VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_aa_ip__programmable_pll
  CLASS BLOCK ;
  FOREIGN sky130_aa_ip__programmable_pll ;
  ORIGIN 172.525 328.515 ;
  SIZE 666.515 BY 935.080 ;
  PIN S6
    ANTENNAGATEAREA 4.600000 ;
    PORT
      LAYER li1 ;
        RECT -110.570 -3.385 -24.980 -3.015 ;
        RECT -25.835 -6.410 -25.575 -3.385 ;
        RECT -21.570 -6.410 -20.730 -6.340 ;
        RECT -25.835 -6.670 -20.730 -6.410 ;
        RECT -21.570 -6.710 -20.730 -6.670 ;
    END
  END S6
  PIN UP_INPUT
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER li1 ;
        RECT 30.055 6.125 30.225 7.440 ;
        RECT 31.035 6.125 31.205 7.440 ;
        RECT 32.015 6.125 32.185 7.440 ;
        RECT 32.995 6.125 33.165 7.440 ;
        RECT 33.975 6.125 34.145 7.440 ;
        RECT 30.055 5.955 34.145 6.125 ;
        RECT 30.055 4.670 30.225 5.955 ;
        RECT 31.035 4.670 31.205 5.955 ;
        RECT 32.015 4.670 32.185 5.955 ;
        RECT 32.995 4.670 33.165 5.955 ;
        RECT 33.975 4.670 34.145 5.955 ;
        RECT 19.925 1.065 20.930 1.325 ;
        RECT -9.030 0.500 20.930 1.065 ;
        RECT -9.030 -9.810 -8.465 0.500 ;
        RECT 19.925 0.380 20.930 0.500 ;
        RECT -131.955 -10.375 -8.465 -9.810 ;
      LAYER met1 ;
        RECT 26.250 7.270 30.260 7.490 ;
        RECT 26.250 6.770 26.470 7.270 ;
        RECT 20.320 6.550 26.470 6.770 ;
        RECT 20.320 1.325 20.540 6.550 ;
        RECT 30.025 6.420 30.255 7.270 ;
        RECT 31.005 6.420 31.235 7.420 ;
        RECT 31.985 6.420 32.215 7.420 ;
        RECT 32.965 6.420 33.195 7.420 ;
        RECT 33.945 6.420 34.175 7.420 ;
        RECT 30.025 4.690 30.255 5.690 ;
        RECT 31.005 4.690 31.235 5.690 ;
        RECT 31.985 4.690 32.215 5.690 ;
        RECT 32.965 4.690 33.195 5.690 ;
        RECT 33.945 4.690 34.175 5.690 ;
        RECT 19.925 0.380 20.930 1.325 ;
    END
  END UP_INPUT
  PIN DN_INPUT
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER li1 ;
        RECT 30.130 -7.325 30.300 -6.010 ;
        RECT 31.110 -7.325 31.280 -6.010 ;
        RECT 32.090 -7.325 32.260 -6.010 ;
        RECT 33.070 -7.325 33.240 -6.010 ;
        RECT 34.050 -7.325 34.220 -6.010 ;
        RECT 30.130 -7.495 34.220 -7.325 ;
        RECT 30.130 -8.780 30.300 -7.495 ;
        RECT 31.110 -8.780 31.280 -7.495 ;
        RECT 32.090 -8.780 32.260 -7.495 ;
        RECT 33.070 -8.780 33.240 -7.495 ;
        RECT 34.050 -8.780 34.220 -7.495 ;
        RECT 21.550 -11.020 22.325 -10.855 ;
        RECT -131.535 -11.500 22.325 -11.020 ;
        RECT 21.550 -11.545 22.325 -11.500 ;
      LAYER met1 ;
        RECT 26.325 -6.180 30.335 -5.960 ;
        RECT 26.325 -6.680 26.545 -6.180 ;
        RECT 21.665 -6.900 26.545 -6.680 ;
        RECT 21.765 -10.855 21.985 -6.900 ;
        RECT 30.100 -7.030 30.330 -6.180 ;
        RECT 31.080 -7.030 31.310 -6.030 ;
        RECT 32.060 -7.030 32.290 -6.030 ;
        RECT 33.040 -7.030 33.270 -6.030 ;
        RECT 34.020 -7.030 34.250 -6.030 ;
        RECT 30.100 -8.760 30.330 -7.760 ;
        RECT 31.080 -8.760 31.310 -7.760 ;
        RECT 32.060 -8.760 32.290 -7.760 ;
        RECT 33.040 -8.760 33.270 -7.760 ;
        RECT 34.020 -8.760 34.250 -7.760 ;
        RECT 21.550 -11.545 22.325 -10.855 ;
    END
  END DN_INPUT
  PIN S2
    ANTENNAGATEAREA 4.600000 ;
    PORT
      LAYER li1 ;
        RECT 21.360 9.355 22.855 9.725 ;
        RECT 22.000 6.330 22.260 9.355 ;
        RECT 26.265 6.330 27.105 6.400 ;
        RECT 22.000 6.215 27.105 6.330 ;
        RECT 21.940 6.070 27.105 6.215 ;
        RECT 21.940 5.330 22.745 6.070 ;
        RECT 26.265 6.030 27.105 6.070 ;
        RECT 21.915 -0.180 22.925 -0.075 ;
        RECT -7.885 -0.425 22.925 -0.180 ;
        RECT -7.905 -0.875 22.925 -0.425 ;
        RECT -7.905 -1.710 -6.615 -0.875 ;
        RECT 21.915 -1.065 22.925 -0.875 ;
        RECT -7.925 -11.965 -6.415 -11.845 ;
        RECT -131.265 -12.665 -6.415 -11.965 ;
        RECT -7.925 -12.920 -6.415 -12.665 ;
      LAYER met1 ;
        RECT 21.940 5.330 22.745 6.215 ;
        RECT 22.040 -0.075 22.535 5.330 ;
        RECT -7.905 -1.710 -6.615 -0.425 ;
        RECT 21.915 -1.065 22.925 -0.075 ;
        RECT -7.585 -11.845 -6.805 -1.710 ;
        RECT -7.925 -12.920 -6.415 -11.845 ;
    END
  END S2
  PIN S3
    ANTENNAGATEAREA 4.600000 ;
    PORT
      LAYER li1 ;
        RECT 16.405 -3.725 17.870 -3.225 ;
        RECT 16.405 -4.095 22.930 -3.725 ;
        RECT 16.405 -4.555 17.870 -4.095 ;
        RECT 22.075 -7.120 22.335 -4.095 ;
        RECT 26.340 -7.120 27.180 -7.050 ;
        RECT 22.075 -7.380 27.180 -7.120 ;
        RECT 26.340 -7.420 27.180 -7.380 ;
        RECT 15.980 -13.140 18.120 -12.695 ;
        RECT -131.055 -14.365 18.120 -13.140 ;
        RECT 15.980 -14.500 18.120 -14.365 ;
      LAYER met1 ;
        RECT 16.405 -4.555 17.870 -3.225 ;
        RECT 16.565 -12.695 17.790 -4.555 ;
        RECT 15.980 -14.500 18.120 -12.695 ;
    END
  END S3
  PIN UP_OUT
    ANTENNADIFFAREA 14.500000 ;
    PORT
      LAYER li1 ;
        RECT 56.560 9.265 56.730 11.305 ;
        RECT 57.740 9.265 57.910 11.305 ;
        RECT 58.920 9.265 59.090 11.305 ;
        RECT 60.100 9.265 60.270 11.305 ;
        RECT 61.280 9.265 61.450 11.305 ;
        RECT 62.460 9.265 62.630 11.305 ;
        RECT 63.640 9.265 63.810 11.305 ;
        RECT 64.820 9.265 64.990 11.305 ;
        RECT 66.000 9.265 66.170 11.305 ;
        RECT 67.180 9.265 67.350 11.305 ;
        RECT 68.360 9.265 68.530 11.305 ;
        RECT 69.540 9.265 69.710 11.305 ;
        RECT 70.720 9.265 70.890 11.305 ;
        RECT 71.900 9.265 72.070 11.305 ;
        RECT 73.080 9.265 73.250 11.305 ;
        RECT 74.260 9.265 74.430 11.305 ;
        RECT 75.440 8.535 75.610 11.305 ;
        RECT 77.610 8.535 78.710 9.165 ;
        RECT 75.440 8.365 78.710 8.535 ;
        RECT 77.610 7.985 78.710 8.365 ;
        RECT 48.400 5.225 48.570 7.265 ;
        RECT 49.580 5.225 49.750 7.265 ;
        RECT 50.760 5.225 50.930 7.265 ;
        RECT 51.940 5.225 52.110 7.265 ;
        RECT 53.120 5.225 53.290 7.265 ;
        RECT 54.300 5.225 54.470 7.265 ;
        RECT 55.480 5.225 55.650 7.265 ;
        RECT 56.660 5.225 56.830 7.265 ;
        RECT 77.200 -14.670 79.265 -14.210 ;
        RECT -130.570 -15.940 79.265 -14.670 ;
        RECT 77.200 -16.055 79.265 -15.940 ;
      LAYER met1 ;
        RECT 56.530 8.930 56.760 11.285 ;
        RECT 57.710 8.930 57.940 11.285 ;
        RECT 58.890 8.930 59.120 11.285 ;
        RECT 60.070 8.930 60.300 11.285 ;
        RECT 61.250 8.930 61.480 11.285 ;
        RECT 62.430 8.930 62.660 11.285 ;
        RECT 63.610 8.930 63.840 11.285 ;
        RECT 64.790 8.930 65.020 11.285 ;
        RECT 65.970 8.930 66.200 11.285 ;
        RECT 67.150 8.930 67.380 11.285 ;
        RECT 68.330 8.930 68.560 11.285 ;
        RECT 69.510 8.930 69.740 11.285 ;
        RECT 70.690 8.930 70.920 11.285 ;
        RECT 71.870 8.930 72.100 11.285 ;
        RECT 73.050 8.930 73.280 11.285 ;
        RECT 74.230 8.930 74.460 11.285 ;
        RECT 75.410 8.930 75.640 11.285 ;
        RECT 56.400 8.560 75.785 8.930 ;
        RECT 56.630 7.980 56.860 8.560 ;
        RECT 77.610 7.985 78.710 9.165 ;
        RECT 48.370 7.750 56.860 7.980 ;
        RECT 48.370 5.245 48.600 7.750 ;
        RECT 49.550 5.245 49.780 7.750 ;
        RECT 50.730 5.245 50.960 7.750 ;
        RECT 51.910 5.245 52.140 7.750 ;
        RECT 53.090 5.245 53.320 7.750 ;
        RECT 54.270 5.245 54.500 7.750 ;
        RECT 55.450 5.245 55.680 7.750 ;
        RECT 56.630 5.245 56.860 7.750 ;
        RECT 77.735 -14.210 78.515 7.985 ;
        RECT 77.200 -16.055 79.265 -14.210 ;
    END
  END UP_OUT
  PIN DN_OUT
    ANTENNADIFFAREA 14.500000 ;
    PORT
      LAYER li1 ;
        RECT 56.355 -4.515 56.525 -2.475 ;
        RECT 57.535 -4.515 57.705 -2.475 ;
        RECT 58.715 -4.515 58.885 -2.475 ;
        RECT 59.895 -4.515 60.065 -2.475 ;
        RECT 61.075 -4.515 61.245 -2.475 ;
        RECT 62.255 -4.515 62.425 -2.475 ;
        RECT 63.435 -4.515 63.605 -2.475 ;
        RECT 64.615 -4.515 64.785 -2.475 ;
        RECT 65.795 -4.515 65.965 -2.475 ;
        RECT 66.975 -4.515 67.145 -2.475 ;
        RECT 68.155 -4.515 68.325 -2.475 ;
        RECT 69.335 -4.515 69.505 -2.475 ;
        RECT 70.515 -4.515 70.685 -2.475 ;
        RECT 71.695 -4.515 71.865 -2.475 ;
        RECT 72.875 -4.515 73.045 -2.475 ;
        RECT 74.055 -4.515 74.225 -2.475 ;
        RECT 75.235 -5.105 75.405 -2.475 ;
        RECT 80.505 -5.105 82.225 -4.355 ;
        RECT 75.235 -5.635 82.225 -5.105 ;
        RECT 80.505 -6.140 82.225 -5.635 ;
        RECT 48.195 -8.555 48.365 -6.515 ;
        RECT 49.375 -8.555 49.545 -6.515 ;
        RECT 50.555 -8.555 50.725 -6.515 ;
        RECT 51.735 -8.555 51.905 -6.515 ;
        RECT 52.915 -8.555 53.085 -6.515 ;
        RECT 54.095 -8.555 54.265 -6.515 ;
        RECT 55.275 -8.555 55.445 -6.515 ;
        RECT 56.455 -8.555 56.625 -6.515 ;
        RECT 80.440 -16.480 82.415 -16.460 ;
        RECT -130.700 -17.930 82.415 -16.480 ;
        RECT 80.440 -18.115 82.415 -17.930 ;
      LAYER met1 ;
        RECT 56.325 -4.850 56.555 -2.495 ;
        RECT 57.505 -4.850 57.735 -2.495 ;
        RECT 58.685 -4.850 58.915 -2.495 ;
        RECT 59.865 -4.850 60.095 -2.495 ;
        RECT 61.045 -4.850 61.275 -2.495 ;
        RECT 62.225 -4.850 62.455 -2.495 ;
        RECT 63.405 -4.850 63.635 -2.495 ;
        RECT 64.585 -4.850 64.815 -2.495 ;
        RECT 65.765 -4.850 65.995 -2.495 ;
        RECT 66.945 -4.850 67.175 -2.495 ;
        RECT 68.125 -4.850 68.355 -2.495 ;
        RECT 69.305 -4.850 69.535 -2.495 ;
        RECT 70.485 -4.850 70.715 -2.495 ;
        RECT 71.665 -4.850 71.895 -2.495 ;
        RECT 72.845 -4.850 73.075 -2.495 ;
        RECT 74.025 -4.850 74.255 -2.495 ;
        RECT 75.205 -4.850 75.435 -2.495 ;
        RECT 56.195 -5.220 75.580 -4.850 ;
        RECT 56.425 -5.800 56.655 -5.220 ;
        RECT 48.165 -6.030 56.655 -5.800 ;
        RECT 48.165 -8.535 48.395 -6.030 ;
        RECT 49.345 -8.535 49.575 -6.030 ;
        RECT 50.525 -8.535 50.755 -6.030 ;
        RECT 51.705 -8.535 51.935 -6.030 ;
        RECT 52.885 -8.535 53.115 -6.030 ;
        RECT 54.065 -8.535 54.295 -6.030 ;
        RECT 55.245 -8.535 55.475 -6.030 ;
        RECT 56.425 -8.535 56.655 -6.030 ;
        RECT 80.505 -6.140 82.225 -4.355 ;
        RECT 80.665 -16.460 81.875 -6.140 ;
        RECT 80.440 -18.115 82.415 -16.460 ;
    END
  END DN_OUT
  PIN ITAIL
    ANTENNAGATEAREA 144.000000 ;
    ANTENNADIFFAREA 2.320000 ;
    PORT
      LAYER li1 ;
        RECT 72.760 39.105 73.975 39.230 ;
        RECT 83.320 39.105 84.805 39.420 ;
        RECT 72.760 38.425 84.805 39.105 ;
        RECT 72.760 38.210 73.975 38.425 ;
        RECT 83.320 38.105 84.805 38.425 ;
        RECT 72.215 30.755 73.455 31.065 ;
        RECT 60.115 30.190 73.455 30.755 ;
        RECT 60.115 28.550 60.680 30.190 ;
        RECT 72.215 30.080 73.455 30.190 ;
        RECT 45.060 27.480 45.490 27.910 ;
        RECT 53.555 27.505 54.185 27.960 ;
        RECT 59.075 27.825 61.475 28.550 ;
        RECT 45.190 23.195 45.360 27.480 ;
        RECT 53.770 23.195 53.940 27.505 ;
        RECT 86.465 -21.680 89.530 -21.175 ;
        RECT 84.875 -21.770 89.530 -21.680 ;
        RECT -131.025 -23.830 89.530 -21.770 ;
        RECT 86.465 -24.240 89.530 -23.830 ;
      LAYER met1 ;
        RECT 72.420 39.280 72.955 39.290 ;
        RECT 72.420 38.745 73.980 39.280 ;
        RECT 72.420 38.210 73.975 38.745 ;
        RECT 72.420 31.065 73.265 38.210 ;
        RECT 72.215 30.080 73.455 31.065 ;
        RECT 45.160 23.215 45.390 27.215 ;
        RECT 53.740 23.215 53.970 27.215 ;
        RECT 82.595 4.545 85.660 40.030 ;
        RECT 82.595 1.480 89.530 4.545 ;
        RECT 86.465 -24.240 89.530 1.480 ;
    END
  END ITAIL
  PIN S4
    ANTENNAGATEAREA 4.600000 ;
    PORT
      LAYER li1 ;
        RECT 90.780 15.550 91.650 15.905 ;
        RECT 90.780 15.180 99.250 15.550 ;
        RECT 90.780 14.925 91.650 15.180 ;
        RECT 98.395 12.155 98.655 15.180 ;
        RECT 102.660 12.155 103.500 12.225 ;
        RECT 98.395 11.895 103.500 12.155 ;
        RECT 102.660 11.855 103.500 11.895 ;
        RECT 89.890 -25.065 92.340 -24.245 ;
        RECT -131.555 -26.995 92.340 -25.065 ;
        RECT 89.890 -27.185 92.340 -26.995 ;
      LAYER met1 ;
        RECT 90.685 15.905 91.620 15.920 ;
        RECT 90.685 14.925 91.650 15.905 ;
        RECT 90.685 -24.245 91.620 14.925 ;
        RECT 89.890 -27.185 92.340 -24.245 ;
    END
  END S4
  PIN VCTRL_IN
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER li1 ;
        RECT 93.145 12.700 93.695 12.745 ;
        RECT 96.705 12.700 97.405 12.895 ;
        RECT 93.145 12.235 97.405 12.700 ;
        RECT 93.145 12.205 93.695 12.235 ;
        RECT 96.705 12.220 97.405 12.235 ;
        RECT 106.450 11.950 106.620 13.265 ;
        RECT 107.430 11.950 107.600 13.265 ;
        RECT 108.410 11.950 108.580 13.265 ;
        RECT 109.390 11.950 109.560 13.265 ;
        RECT 110.370 11.950 110.540 13.265 ;
        RECT 106.450 11.780 110.540 11.950 ;
        RECT 106.450 10.495 106.620 11.780 ;
        RECT 107.430 10.495 107.600 11.780 ;
        RECT 108.410 10.495 108.580 11.780 ;
        RECT 109.390 10.495 109.560 11.780 ;
        RECT 110.370 10.495 110.540 11.780 ;
        RECT 92.670 -28.320 94.950 -27.935 ;
        RECT -131.605 -30.310 94.950 -28.320 ;
        RECT -131.605 -30.490 93.520 -30.310 ;
      LAYER met1 ;
        RECT 102.645 13.095 106.655 13.315 ;
        RECT 93.105 -27.660 93.790 12.785 ;
        RECT 96.705 12.595 97.405 12.895 ;
        RECT 102.645 12.595 102.865 13.095 ;
        RECT 96.705 12.375 102.865 12.595 ;
        RECT 96.705 12.220 97.405 12.375 ;
        RECT 106.420 12.245 106.650 13.095 ;
        RECT 107.400 12.245 107.630 13.245 ;
        RECT 108.380 12.245 108.610 13.245 ;
        RECT 109.360 12.245 109.590 13.245 ;
        RECT 110.340 12.245 110.570 13.245 ;
        RECT 106.420 10.515 106.650 11.515 ;
        RECT 107.400 10.515 107.630 11.515 ;
        RECT 108.380 10.515 108.610 11.515 ;
        RECT 109.360 10.515 109.590 11.515 ;
        RECT 110.340 10.515 110.570 11.515 ;
        RECT 92.120 -30.855 95.405 -27.660 ;
    END
  END VCTRL_IN
  PIN LF_OFFCHIP
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER li1 ;
        RECT 107.310 -4.800 107.480 -3.485 ;
        RECT 108.290 -4.800 108.460 -3.485 ;
        RECT 109.270 -4.800 109.440 -3.485 ;
        RECT 110.250 -4.800 110.420 -3.485 ;
        RECT 111.230 -4.800 111.400 -3.485 ;
        RECT 107.310 -4.970 111.400 -4.800 ;
        RECT 107.310 -6.255 107.480 -4.970 ;
        RECT 108.290 -6.255 108.460 -4.970 ;
        RECT 109.270 -6.255 109.440 -4.970 ;
        RECT 110.250 -6.255 110.420 -4.970 ;
        RECT 111.230 -6.255 111.400 -4.970 ;
        RECT 94.745 -31.730 98.055 -31.465 ;
        RECT -133.265 -33.935 98.055 -31.730 ;
        RECT 94.745 -34.250 98.055 -33.935 ;
      LAYER met1 ;
        RECT 103.505 -3.655 107.515 -3.435 ;
        RECT 96.060 -4.155 96.795 -4.145 ;
        RECT 103.505 -4.155 103.725 -3.655 ;
        RECT 96.060 -4.375 103.725 -4.155 ;
        RECT 96.060 -31.465 97.710 -4.375 ;
        RECT 107.280 -4.505 107.510 -3.655 ;
        RECT 108.260 -4.505 108.490 -3.505 ;
        RECT 109.240 -4.505 109.470 -3.505 ;
        RECT 110.220 -4.505 110.450 -3.505 ;
        RECT 111.200 -4.505 111.430 -3.505 ;
        RECT 107.280 -6.235 107.510 -5.235 ;
        RECT 108.260 -6.235 108.490 -5.235 ;
        RECT 109.240 -6.235 109.470 -5.235 ;
        RECT 110.220 -6.235 110.450 -5.235 ;
        RECT 111.200 -6.235 111.430 -5.235 ;
        RECT 94.745 -34.250 98.055 -31.465 ;
    END
  END LF_OFFCHIP
  PIN S5
    ANTENNAGATEAREA 4.600000 ;
    PORT
      LAYER li1 ;
        RECT 98.615 -1.570 100.110 -1.200 ;
        RECT 99.255 -4.580 99.515 -1.570 ;
        RECT 99.180 -4.595 100.490 -4.580 ;
        RECT 103.520 -4.595 104.360 -4.525 ;
        RECT 99.180 -4.855 104.360 -4.595 ;
        RECT 99.180 -5.645 100.490 -4.855 ;
        RECT 103.520 -4.895 104.360 -4.855 ;
        RECT 99.180 -6.395 100.465 -5.645 ;
        RECT 98.325 -35.500 101.475 -35.125 ;
        RECT -133.730 -37.965 101.475 -35.500 ;
        RECT 98.325 -38.170 101.475 -37.965 ;
      LAYER met1 ;
        RECT 99.180 -6.395 100.465 -4.950 ;
        RECT 99.340 -35.125 100.330 -6.395 ;
        RECT 98.325 -38.170 101.475 -35.125 ;
    END
  END S5
  PIN OUT_CORE
    ANTENNADIFFAREA 14.500000 ;
    PORT
      LAYER li1 ;
        RECT -161.125 -165.950 -130.700 -164.860 ;
        RECT -131.735 -169.465 -130.700 -165.950 ;
        RECT -130.980 -170.095 -130.810 -169.465 ;
        RECT -130.980 -170.265 -128.040 -170.095 ;
        RECT -130.080 -171.445 -128.040 -171.275 ;
        RECT -130.080 -172.625 -128.040 -172.455 ;
        RECT -130.080 -173.805 -128.040 -173.635 ;
        RECT -130.080 -174.985 -128.040 -174.815 ;
        RECT -130.080 -176.165 -128.040 -175.995 ;
        RECT -130.080 -177.345 -128.040 -177.175 ;
        RECT -130.080 -178.525 -128.040 -178.355 ;
        RECT -130.080 -179.705 -128.040 -179.535 ;
        RECT -130.080 -180.885 -128.040 -180.715 ;
        RECT -130.080 -182.065 -128.040 -181.895 ;
        RECT -130.080 -183.245 -128.040 -183.075 ;
        RECT -130.080 -184.425 -128.040 -184.255 ;
        RECT -130.080 -185.605 -128.040 -185.435 ;
        RECT -130.080 -186.785 -128.040 -186.615 ;
        RECT -130.080 -187.965 -128.040 -187.795 ;
        RECT -134.120 -189.045 -132.080 -188.875 ;
        RECT -130.080 -189.145 -128.040 -188.975 ;
        RECT -134.120 -190.225 -132.080 -190.055 ;
        RECT -134.120 -191.405 -132.080 -191.235 ;
        RECT -134.120 -192.585 -132.080 -192.415 ;
        RECT -134.120 -193.765 -132.080 -193.595 ;
        RECT -134.120 -194.945 -132.080 -194.775 ;
        RECT -134.120 -196.125 -132.080 -195.955 ;
        RECT -134.120 -197.305 -132.080 -197.135 ;
      LAYER met1 ;
        RECT -130.785 -170.065 -130.415 -169.920 ;
        RECT -130.785 -170.295 -128.060 -170.065 ;
        RECT -130.785 -171.245 -130.415 -170.295 ;
        RECT -130.785 -171.475 -128.060 -171.245 ;
        RECT -130.785 -172.425 -130.415 -171.475 ;
        RECT -130.785 -172.655 -128.060 -172.425 ;
        RECT -130.785 -173.605 -130.415 -172.655 ;
        RECT -130.785 -173.835 -128.060 -173.605 ;
        RECT -130.785 -174.785 -130.415 -173.835 ;
        RECT -130.785 -175.015 -128.060 -174.785 ;
        RECT -130.785 -175.965 -130.415 -175.015 ;
        RECT -130.785 -176.195 -128.060 -175.965 ;
        RECT -130.785 -177.145 -130.415 -176.195 ;
        RECT -130.785 -177.375 -128.060 -177.145 ;
        RECT -130.785 -178.325 -130.415 -177.375 ;
        RECT -130.785 -178.555 -128.060 -178.325 ;
        RECT -130.785 -179.505 -130.415 -178.555 ;
        RECT -130.785 -179.735 -128.060 -179.505 ;
        RECT -130.785 -180.685 -130.415 -179.735 ;
        RECT -130.785 -180.915 -128.060 -180.685 ;
        RECT -130.785 -181.865 -130.415 -180.915 ;
        RECT -130.785 -182.095 -128.060 -181.865 ;
        RECT -130.785 -183.045 -130.415 -182.095 ;
        RECT -130.785 -183.275 -128.060 -183.045 ;
        RECT -130.785 -184.225 -130.415 -183.275 ;
        RECT -130.785 -184.455 -128.060 -184.225 ;
        RECT -130.785 -185.405 -130.415 -184.455 ;
        RECT -130.785 -185.635 -128.060 -185.405 ;
        RECT -130.785 -186.585 -130.415 -185.635 ;
        RECT -130.785 -186.815 -128.060 -186.585 ;
        RECT -130.785 -187.765 -130.415 -186.815 ;
        RECT -130.785 -187.995 -128.060 -187.765 ;
        RECT -130.785 -188.845 -130.415 -187.995 ;
        RECT -134.100 -188.945 -130.415 -188.845 ;
        RECT -134.100 -189.075 -128.060 -188.945 ;
        RECT -131.595 -190.025 -131.365 -189.075 ;
        RECT -130.785 -189.175 -128.060 -189.075 ;
        RECT -130.785 -189.305 -130.415 -189.175 ;
        RECT -134.100 -190.255 -131.365 -190.025 ;
        RECT -131.595 -191.205 -131.365 -190.255 ;
        RECT -134.100 -191.435 -131.365 -191.205 ;
        RECT -131.595 -192.385 -131.365 -191.435 ;
        RECT -134.100 -192.615 -131.365 -192.385 ;
        RECT -131.595 -193.565 -131.365 -192.615 ;
        RECT -134.100 -193.795 -131.365 -193.565 ;
        RECT -131.595 -194.745 -131.365 -193.795 ;
        RECT -134.100 -194.975 -131.365 -194.745 ;
        RECT -131.595 -195.925 -131.365 -194.975 ;
        RECT -134.100 -196.155 -131.365 -195.925 ;
        RECT -131.595 -197.105 -131.365 -196.155 ;
        RECT -134.100 -197.335 -131.365 -197.105 ;
    END
  END OUT_CORE
  PIN OUT_USB
    ANTENNADIFFAREA 14.500000 ;
    PORT
      LAYER li1 ;
        RECT -163.880 -254.235 -139.430 -253.340 ;
        RECT -140.325 -260.080 -139.430 -254.235 ;
        RECT -140.080 -260.820 -139.910 -260.080 ;
        RECT -140.080 -260.990 -137.140 -260.820 ;
        RECT -139.180 -262.170 -137.140 -262.000 ;
        RECT -139.180 -263.350 -137.140 -263.180 ;
        RECT -139.180 -264.530 -137.140 -264.360 ;
        RECT -139.180 -265.710 -137.140 -265.540 ;
        RECT -139.180 -266.890 -137.140 -266.720 ;
        RECT -139.180 -268.070 -137.140 -267.900 ;
        RECT -139.180 -269.250 -137.140 -269.080 ;
        RECT -139.180 -270.430 -137.140 -270.260 ;
        RECT -139.180 -271.610 -137.140 -271.440 ;
        RECT -139.180 -272.790 -137.140 -272.620 ;
        RECT -139.180 -273.970 -137.140 -273.800 ;
        RECT -139.180 -275.150 -137.140 -274.980 ;
        RECT -139.180 -276.330 -137.140 -276.160 ;
        RECT -139.180 -277.510 -137.140 -277.340 ;
        RECT -139.180 -278.690 -137.140 -278.520 ;
        RECT -143.220 -279.770 -141.180 -279.600 ;
        RECT -139.180 -279.870 -137.140 -279.700 ;
        RECT -143.220 -280.950 -141.180 -280.780 ;
        RECT -143.220 -282.130 -141.180 -281.960 ;
        RECT -143.220 -283.310 -141.180 -283.140 ;
        RECT -143.220 -284.490 -141.180 -284.320 ;
        RECT -143.220 -285.670 -141.180 -285.500 ;
        RECT -143.220 -286.850 -141.180 -286.680 ;
        RECT -143.220 -288.030 -141.180 -287.860 ;
      LAYER met1 ;
        RECT -139.885 -260.790 -139.515 -260.645 ;
        RECT -139.885 -261.020 -137.160 -260.790 ;
        RECT -139.885 -261.970 -139.515 -261.020 ;
        RECT -139.885 -262.200 -137.160 -261.970 ;
        RECT -139.885 -263.150 -139.515 -262.200 ;
        RECT -139.885 -263.380 -137.160 -263.150 ;
        RECT -139.885 -264.330 -139.515 -263.380 ;
        RECT -139.885 -264.560 -137.160 -264.330 ;
        RECT -139.885 -265.510 -139.515 -264.560 ;
        RECT -139.885 -265.740 -137.160 -265.510 ;
        RECT -139.885 -266.690 -139.515 -265.740 ;
        RECT -139.885 -266.920 -137.160 -266.690 ;
        RECT -139.885 -267.870 -139.515 -266.920 ;
        RECT -139.885 -268.100 -137.160 -267.870 ;
        RECT -139.885 -269.050 -139.515 -268.100 ;
        RECT -139.885 -269.280 -137.160 -269.050 ;
        RECT -139.885 -270.230 -139.515 -269.280 ;
        RECT -139.885 -270.460 -137.160 -270.230 ;
        RECT -139.885 -271.410 -139.515 -270.460 ;
        RECT -139.885 -271.640 -137.160 -271.410 ;
        RECT -139.885 -272.590 -139.515 -271.640 ;
        RECT -139.885 -272.820 -137.160 -272.590 ;
        RECT -139.885 -273.770 -139.515 -272.820 ;
        RECT -139.885 -274.000 -137.160 -273.770 ;
        RECT -139.885 -274.950 -139.515 -274.000 ;
        RECT -139.885 -275.180 -137.160 -274.950 ;
        RECT -139.885 -276.130 -139.515 -275.180 ;
        RECT -139.885 -276.360 -137.160 -276.130 ;
        RECT -139.885 -277.310 -139.515 -276.360 ;
        RECT -139.885 -277.540 -137.160 -277.310 ;
        RECT -139.885 -278.490 -139.515 -277.540 ;
        RECT -139.885 -278.720 -137.160 -278.490 ;
        RECT -139.885 -279.570 -139.515 -278.720 ;
        RECT -143.200 -279.670 -139.515 -279.570 ;
        RECT -143.200 -279.800 -137.160 -279.670 ;
        RECT -140.695 -280.750 -140.465 -279.800 ;
        RECT -139.885 -279.900 -137.160 -279.800 ;
        RECT -139.885 -280.030 -139.515 -279.900 ;
        RECT -143.200 -280.980 -140.465 -280.750 ;
        RECT -140.695 -281.930 -140.465 -280.980 ;
        RECT -143.200 -282.160 -140.465 -281.930 ;
        RECT -140.695 -283.110 -140.465 -282.160 ;
        RECT -143.200 -283.340 -140.465 -283.110 ;
        RECT -140.695 -284.290 -140.465 -283.340 ;
        RECT -143.200 -284.520 -140.465 -284.290 ;
        RECT -140.695 -285.470 -140.465 -284.520 ;
        RECT -143.200 -285.700 -140.465 -285.470 ;
        RECT -140.695 -286.650 -140.465 -285.700 ;
        RECT -143.200 -286.880 -140.465 -286.650 ;
        RECT -140.695 -287.830 -140.465 -286.880 ;
        RECT -143.200 -288.060 -140.465 -287.830 ;
    END
  END OUT_USB
  PIN D12
    ANTENNAGATEAREA 10.500000 ;
    PORT
      LAYER li1 ;
        RECT -115.930 -180.955 -115.625 -179.940 ;
        RECT -107.965 -180.955 -107.290 -180.890 ;
        RECT -115.930 -181.125 -107.290 -180.955 ;
        RECT -115.930 -181.130 -115.625 -181.125 ;
        RECT -107.965 -181.160 -107.290 -181.125 ;
        RECT -32.210 -182.275 -31.270 -181.905 ;
        RECT -67.240 -188.225 -66.885 -188.220 ;
        RECT -65.180 -188.225 -64.810 -188.195 ;
        RECT -67.240 -188.230 -64.810 -188.225 ;
        RECT -68.370 -188.420 -64.810 -188.230 ;
        RECT -68.370 -188.430 -67.235 -188.420 ;
        RECT -65.180 -188.550 -64.810 -188.420 ;
        RECT -67.920 -195.575 -67.270 -195.490 ;
        RECT -67.050 -195.575 -66.685 -195.510 ;
        RECT -67.920 -195.780 -66.685 -195.575 ;
        RECT -67.920 -196.240 -67.270 -195.780 ;
        RECT -67.050 -195.810 -66.685 -195.780 ;
        RECT -115.930 -208.555 -115.630 -207.650 ;
        RECT -115.930 -208.760 -106.485 -208.555 ;
        RECT -115.930 -208.835 -115.630 -208.760 ;
        RECT -106.785 -208.785 -106.485 -208.760 ;
        RECT -106.785 -209.065 -106.060 -208.785 ;
        RECT 137.685 -210.385 138.360 -210.355 ;
        RECT 137.585 -210.395 138.360 -210.385 ;
        RECT 134.945 -210.575 138.360 -210.395 ;
        RECT 156.025 -210.540 156.700 -210.510 ;
        RECT 155.925 -210.550 156.700 -210.540 ;
        RECT 42.750 -211.215 43.365 -211.210 ;
        RECT 42.745 -211.430 43.365 -211.215 ;
        RECT 42.745 -215.470 43.035 -211.430 ;
        RECT -31.830 -217.370 -31.135 -217.100 ;
        RECT -26.440 -217.340 -25.745 -217.070 ;
        RECT 42.750 -222.520 43.030 -215.470 ;
        RECT 135.860 -215.710 136.540 -210.575 ;
        RECT 137.585 -210.585 138.360 -210.575 ;
        RECT 137.685 -210.625 138.360 -210.585 ;
        RECT 153.855 -210.730 156.700 -210.550 ;
        RECT 153.855 -215.710 154.535 -210.730 ;
        RECT 155.925 -210.740 156.700 -210.730 ;
        RECT 156.025 -210.780 156.700 -210.740 ;
        RECT 135.860 -216.390 154.535 -215.710 ;
        RECT 135.860 -222.520 136.540 -216.390 ;
        RECT -162.170 -223.200 136.540 -222.520 ;
      LAYER met1 ;
        RECT -115.930 -222.575 -115.625 -179.940 ;
        RECT -32.210 -182.275 -31.530 -181.905 ;
        RECT -32.210 -184.185 -31.955 -182.275 ;
        RECT -32.210 -184.440 47.115 -184.185 ;
        RECT -68.385 -188.470 -67.400 -188.200 ;
        RECT -67.670 -193.625 -67.400 -188.470 ;
        RECT -75.725 -194.505 -67.400 -193.625 ;
        RECT -116.195 -223.190 -115.580 -222.575 ;
        RECT -75.725 -223.200 -74.845 -194.505 ;
        RECT -67.670 -195.490 -67.400 -194.505 ;
        RECT -67.920 -196.240 -67.270 -195.490 ;
        RECT 46.860 -211.190 47.115 -184.440 ;
        RECT -23.925 -211.445 47.115 -211.190 ;
        RECT -31.830 -217.185 -31.135 -217.100 ;
        RECT -26.440 -217.185 -25.745 -217.070 ;
        RECT -31.830 -217.195 -25.745 -217.185 ;
        RECT -23.925 -217.195 -23.785 -211.445 ;
        RECT -31.830 -217.325 -23.785 -217.195 ;
        RECT -31.830 -217.370 -31.135 -217.325 ;
        RECT -26.440 -217.335 -23.785 -217.325 ;
        RECT -26.440 -217.340 -25.745 -217.335 ;
    END
  END D12
  PIN D13
    ANTENNAGATEAREA 7.200000 ;
    PORT
      LAYER li1 ;
        RECT 33.170 -178.530 33.865 -178.260 ;
        RECT 38.560 -178.560 39.255 -178.290 ;
        RECT -114.975 -180.545 -114.670 -179.545 ;
        RECT -108.905 -180.545 -108.230 -180.500 ;
        RECT -114.975 -180.735 -108.230 -180.545 ;
        RECT -108.905 -180.770 -108.230 -180.735 ;
        RECT -114.975 -209.000 -114.675 -208.935 ;
        RECT -108.385 -209.000 -107.660 -208.945 ;
        RECT -114.975 -209.205 -107.660 -209.000 ;
        RECT -114.975 -210.120 -114.675 -209.205 ;
        RECT -108.385 -209.225 -107.660 -209.205 ;
        RECT 179.885 -210.440 180.560 -210.410 ;
        RECT 179.785 -210.450 180.560 -210.440 ;
        RECT 177.145 -210.630 180.560 -210.450 ;
        RECT 198.225 -210.595 198.900 -210.565 ;
        RECT 198.125 -210.605 198.900 -210.595 ;
        RECT 178.060 -215.765 178.740 -210.630 ;
        RECT 179.785 -210.640 180.560 -210.630 ;
        RECT 179.885 -210.680 180.560 -210.640 ;
        RECT 196.055 -210.785 198.900 -210.605 ;
        RECT 196.055 -215.765 196.735 -210.785 ;
        RECT 198.125 -210.795 198.900 -210.785 ;
        RECT 198.225 -210.835 198.900 -210.795 ;
        RECT 178.060 -216.445 196.735 -215.765 ;
        RECT 33.170 -217.370 33.865 -217.100 ;
        RECT 38.560 -217.340 39.255 -217.070 ;
        RECT 43.245 -217.360 43.570 -216.675 ;
        RECT 43.260 -221.160 43.530 -217.360 ;
        RECT 178.060 -223.515 178.740 -216.445 ;
        RECT -162.250 -224.195 178.740 -223.515 ;
      LAYER met1 ;
        RECT 33.170 -178.305 33.865 -178.260 ;
        RECT 38.560 -178.295 39.255 -178.290 ;
        RECT 38.050 -178.305 51.105 -178.295 ;
        RECT 33.170 -178.435 51.105 -178.305 ;
        RECT 33.170 -178.445 39.255 -178.435 ;
        RECT 33.170 -178.530 33.865 -178.445 ;
        RECT 38.560 -178.560 39.255 -178.445 ;
        RECT -114.975 -223.570 -114.670 -179.545 ;
        RECT 33.170 -217.185 33.865 -217.100 ;
        RECT 38.560 -217.185 39.255 -217.070 ;
        RECT 33.170 -217.195 39.255 -217.185 ;
        RECT 43.245 -217.195 43.570 -216.675 ;
        RECT 50.965 -217.195 51.105 -178.435 ;
        RECT 33.170 -217.325 51.105 -217.195 ;
        RECT 33.170 -217.370 33.865 -217.325 ;
        RECT 38.050 -217.335 51.105 -217.325 ;
        RECT 38.560 -217.340 39.255 -217.335 ;
        RECT 43.245 -217.360 43.570 -217.335 ;
        RECT 43.220 -223.545 43.525 -220.525 ;
        RECT -115.240 -224.185 -114.625 -223.570 ;
        RECT 42.955 -224.160 43.570 -223.545 ;
    END
  END D13
  PIN D14
    ANTENNAGATEAREA 7.200000 ;
    PORT
      LAYER li1 ;
        RECT 18.170 -178.530 18.865 -178.260 ;
        RECT 23.560 -178.560 24.255 -178.290 ;
        RECT -114.430 -180.130 -114.125 -179.115 ;
        RECT -110.585 -180.130 -109.910 -180.090 ;
        RECT -114.430 -180.305 -109.910 -180.130 ;
        RECT -110.680 -180.315 -109.910 -180.305 ;
        RECT -110.585 -180.360 -109.910 -180.315 ;
        RECT -114.425 -209.460 -114.125 -209.450 ;
        RECT -110.030 -209.460 -109.305 -209.420 ;
        RECT -114.425 -209.665 -109.305 -209.460 ;
        RECT -114.425 -210.635 -114.125 -209.665 ;
        RECT -110.030 -209.700 -109.305 -209.665 ;
        RECT 224.200 -210.635 224.875 -210.605 ;
        RECT 224.100 -210.645 224.875 -210.635 ;
        RECT 221.460 -210.825 224.875 -210.645 ;
        RECT 242.540 -210.790 243.215 -210.760 ;
        RECT 242.440 -210.800 243.215 -210.790 ;
        RECT 43.465 -214.220 44.080 -214.000 ;
        RECT 18.170 -217.370 18.865 -217.100 ;
        RECT 23.560 -217.340 24.255 -217.070 ;
        RECT 43.785 -221.160 44.055 -214.220 ;
        RECT 222.375 -215.890 223.055 -210.825 ;
        RECT 224.100 -210.835 224.875 -210.825 ;
        RECT 224.200 -210.875 224.875 -210.835 ;
        RECT 240.370 -210.980 243.215 -210.800 ;
        RECT 222.375 -215.960 223.290 -215.890 ;
        RECT 240.370 -215.960 241.050 -210.980 ;
        RECT 242.440 -210.990 243.215 -210.980 ;
        RECT 242.540 -211.030 243.215 -210.990 ;
        RECT 222.375 -216.640 241.050 -215.960 ;
        RECT 222.610 -224.680 223.290 -216.640 ;
        RECT -162.290 -225.360 223.290 -224.680 ;
      LAYER met1 ;
        RECT 18.170 -178.305 18.865 -178.260 ;
        RECT 23.560 -178.295 24.255 -178.290 ;
        RECT 23.560 -178.305 30.355 -178.295 ;
        RECT 18.170 -178.435 30.355 -178.305 ;
        RECT 18.170 -178.445 24.255 -178.435 ;
        RECT 18.170 -178.530 18.865 -178.445 ;
        RECT 23.560 -178.560 24.255 -178.445 ;
        RECT -114.430 -180.305 -114.125 -179.115 ;
        RECT -114.430 -209.450 -114.130 -180.305 ;
        RECT 30.215 -181.425 30.355 -178.435 ;
        RECT 30.215 -181.565 50.350 -181.425 ;
        RECT -114.430 -210.635 -114.125 -209.450 ;
        RECT -114.430 -224.735 -114.130 -210.635 ;
        RECT 43.420 -214.065 44.115 -213.990 ;
        RECT 50.210 -214.065 50.350 -181.565 ;
        RECT 30.215 -214.205 50.350 -214.065 ;
        RECT 18.170 -217.185 18.865 -217.100 ;
        RECT 23.560 -217.185 24.255 -217.070 ;
        RECT 18.170 -217.195 24.255 -217.185 ;
        RECT 30.215 -217.195 30.355 -214.205 ;
        RECT 43.420 -214.225 44.115 -214.205 ;
        RECT 18.170 -217.325 30.355 -217.195 ;
        RECT 18.170 -217.370 18.865 -217.325 ;
        RECT 23.560 -217.335 30.355 -217.325 ;
        RECT 23.560 -217.340 24.255 -217.335 ;
        RECT 43.810 -220.545 44.030 -220.530 ;
        RECT 43.765 -224.710 44.065 -220.545 ;
        RECT -114.710 -225.350 -114.095 -224.735 ;
        RECT 43.485 -225.325 44.100 -224.710 ;
    END
  END D14
  PIN D15
    ANTENNAGATEAREA 7.000000 ;
    PORT
      LAYER li1 ;
        RECT -101.305 -181.730 -100.620 -181.710 ;
        RECT -101.495 -181.740 -100.360 -181.730 ;
        RECT -98.305 -181.740 -97.935 -181.610 ;
        RECT -101.495 -181.930 -97.935 -181.740 ;
        RECT -101.305 -182.000 -100.620 -181.930 ;
        RECT -100.365 -181.935 -97.935 -181.930 ;
        RECT -100.365 -181.940 -100.010 -181.935 ;
        RECT -98.305 -181.965 -97.935 -181.935 ;
        RECT -113.935 -185.325 -113.635 -184.945 ;
        RECT -113.935 -185.525 -113.595 -185.325 ;
        RECT -113.935 -185.910 -113.635 -185.525 ;
        RECT -101.850 -185.910 -101.190 -185.865 ;
        RECT -113.935 -186.110 -101.190 -185.910 ;
        RECT -113.935 -186.130 -113.635 -186.110 ;
        RECT -101.850 -186.130 -101.190 -186.110 ;
        RECT 33.220 -189.785 33.915 -189.515 ;
        RECT 38.610 -189.815 39.305 -189.545 ;
        RECT 33.220 -206.115 33.915 -205.845 ;
        RECT 38.610 -206.085 39.305 -205.815 ;
        RECT 44.165 -206.140 44.890 -205.465 ;
        RECT -104.460 -207.245 -104.170 -206.770 ;
        RECT -102.425 -207.245 -101.710 -207.210 ;
        RECT -104.460 -207.425 -101.710 -207.245 ;
        RECT -104.460 -207.455 -104.170 -207.425 ;
        RECT -102.425 -207.510 -101.710 -207.425 ;
        RECT -113.935 -212.480 -113.645 -212.000 ;
        RECT -104.560 -212.480 -104.270 -212.000 ;
        RECT -113.935 -212.685 -104.270 -212.480 ;
        RECT 44.280 -222.245 44.560 -206.140 ;
        RECT 270.190 -210.465 270.865 -210.435 ;
        RECT 270.090 -210.475 270.865 -210.465 ;
        RECT 267.450 -210.655 270.865 -210.475 ;
        RECT 288.530 -210.620 289.205 -210.590 ;
        RECT 288.430 -210.630 289.205 -210.620 ;
        RECT 268.365 -215.790 269.045 -210.655 ;
        RECT 270.090 -210.665 270.865 -210.655 ;
        RECT 270.190 -210.705 270.865 -210.665 ;
        RECT 286.360 -210.810 289.205 -210.630 ;
        RECT 286.360 -215.790 287.040 -210.810 ;
        RECT 288.430 -210.820 289.205 -210.810 ;
        RECT 288.530 -210.860 289.205 -210.820 ;
        RECT 268.365 -216.470 287.040 -215.790 ;
        RECT 268.365 -225.955 269.045 -216.470 ;
        RECT -162.410 -226.635 269.045 -225.955 ;
      LAYER met1 ;
        RECT -101.305 -182.000 -100.620 -181.710 ;
        RECT -113.935 -226.020 -113.630 -184.940 ;
        RECT -101.270 -185.865 -101.070 -182.000 ;
        RECT -101.850 -185.910 -101.070 -185.865 ;
        RECT -102.085 -186.110 -101.070 -185.910 ;
        RECT -101.850 -186.130 -101.190 -186.110 ;
        RECT 33.220 -189.560 33.915 -189.515 ;
        RECT 38.610 -189.550 39.305 -189.545 ;
        RECT 45.260 -189.550 45.515 -189.510 ;
        RECT 38.610 -189.560 45.515 -189.550 ;
        RECT 33.220 -189.690 45.515 -189.560 ;
        RECT 33.220 -189.700 39.305 -189.690 ;
        RECT 33.220 -189.785 33.915 -189.700 ;
        RECT 38.610 -189.815 39.305 -189.700 ;
        RECT 45.260 -189.765 45.515 -189.690 ;
        RECT 33.220 -205.930 33.915 -205.845 ;
        RECT 38.610 -205.930 39.305 -205.815 ;
        RECT 33.220 -205.940 39.305 -205.930 ;
        RECT 44.165 -205.940 44.890 -205.465 ;
        RECT 45.325 -205.940 45.465 -189.765 ;
        RECT 33.220 -206.070 45.475 -205.940 ;
        RECT 33.220 -206.115 33.915 -206.070 ;
        RECT 38.610 -206.080 45.475 -206.070 ;
        RECT 38.610 -206.085 39.305 -206.080 ;
        RECT 44.165 -206.140 44.890 -206.080 ;
        RECT -104.460 -207.455 -104.170 -206.770 ;
        RECT -104.460 -212.000 -104.285 -207.455 ;
        RECT -104.560 -212.685 -104.270 -212.000 ;
        RECT 44.260 -225.995 44.565 -221.260 ;
        RECT -114.245 -226.635 -113.625 -226.020 ;
        RECT 43.950 -226.610 44.570 -225.995 ;
    END
  END D15
  PIN F_IN
    ANTENNAGATEAREA 34.399998 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT -42.225 569.660 -41.955 570.335 ;
        RECT -42.185 569.560 -41.985 569.660 ;
        RECT -42.175 567.465 -41.995 569.560 ;
        RECT -70.960 562.895 -69.770 563.180 ;
        RECT -42.550 562.895 -41.080 567.465 ;
        RECT -70.960 561.425 -41.080 562.895 ;
        RECT -70.960 561.180 -69.770 561.425 ;
        RECT -42.415 522.840 -42.145 523.515 ;
        RECT -42.375 522.740 -42.175 522.840 ;
        RECT -42.365 520.160 -42.185 522.740 ;
        RECT -70.980 517.765 -69.755 518.325 ;
        RECT -42.715 517.765 -41.790 520.160 ;
        RECT -70.980 516.840 -41.790 517.765 ;
        RECT -70.980 516.415 -69.755 516.840 ;
        RECT -42.500 477.075 -42.230 477.750 ;
        RECT -42.460 476.975 -42.260 477.075 ;
        RECT -42.450 474.830 -42.270 476.975 ;
        RECT -70.930 471.395 -69.770 471.630 ;
        RECT -42.845 471.395 -41.650 474.830 ;
        RECT -70.930 470.200 -41.650 471.395 ;
        RECT -70.930 469.890 -69.770 470.200 ;
        RECT -42.830 433.305 -42.560 433.980 ;
        RECT -42.790 433.205 -42.590 433.305 ;
        RECT -42.780 431.210 -42.600 433.205 ;
        RECT -70.870 428.295 -69.845 428.555 ;
        RECT -43.005 428.295 -42.275 431.210 ;
        RECT -70.870 427.565 -42.275 428.295 ;
        RECT -70.870 427.395 -69.845 427.565 ;
        RECT -43.000 387.315 -42.730 387.990 ;
        RECT -42.960 387.215 -42.760 387.315 ;
        RECT -42.950 384.805 -42.770 387.215 ;
        RECT -70.735 381.700 -70.040 381.960 ;
        RECT -43.465 381.700 -42.735 384.805 ;
        RECT -70.735 380.970 -42.735 381.700 ;
        RECT -70.735 380.700 -70.040 380.970 ;
        RECT -42.805 343.000 -42.535 343.675 ;
        RECT -42.765 342.900 -42.565 343.000 ;
        RECT -42.755 340.800 -42.575 342.900 ;
        RECT -70.965 338.290 -69.950 338.585 ;
        RECT -43.035 338.290 -42.305 340.800 ;
        RECT -70.965 337.560 -42.305 338.290 ;
        RECT -70.965 337.215 -69.950 337.560 ;
        RECT -36.010 305.795 -35.740 306.470 ;
        RECT -35.980 305.695 -35.780 305.795 ;
        RECT -35.970 304.660 -35.790 305.695 ;
        RECT -42.750 300.800 -42.480 301.475 ;
        RECT -42.710 300.700 -42.510 300.800 ;
        RECT -42.700 298.850 -42.520 300.700 ;
        RECT -43.065 297.555 -41.750 298.850 ;
        RECT -70.850 296.085 -69.875 297.190 ;
        RECT -42.990 293.225 -41.965 297.555 ;
        RECT -34.010 294.610 -33.115 298.855 ;
        RECT -34.170 292.960 -32.700 294.610 ;
        RECT -44.115 277.415 -43.745 278.255 ;
        RECT -44.060 277.115 -43.770 277.415 ;
        RECT -41.775 277.360 -41.580 288.255 ;
        RECT -44.065 276.815 -43.405 277.115 ;
        RECT -41.825 276.675 -41.525 277.360 ;
        RECT -41.775 272.630 -41.580 276.675 ;
        RECT -41.830 271.970 -41.530 272.630 ;
        RECT -40.370 272.185 -39.260 272.485 ;
        RECT -44.115 259.800 -43.745 260.345 ;
        RECT -41.775 260.135 -41.580 271.970 ;
        RECT -39.575 271.345 -39.205 272.185 ;
        RECT -39.905 260.135 -39.230 260.265 ;
        RECT -41.775 259.800 -39.230 260.135 ;
        RECT -44.115 259.605 -39.230 259.800 ;
        RECT -44.115 259.505 -43.745 259.605 ;
        RECT -33.815 252.660 -32.585 252.845 ;
        RECT -39.045 251.950 -32.585 252.660 ;
        RECT -39.045 251.765 -38.100 251.950 ;
        RECT -33.815 251.755 -32.585 251.950 ;
        RECT -64.520 236.720 -64.325 247.615 ;
        RECT -34.140 243.455 -32.800 244.075 ;
        RECT -34.150 242.900 -32.800 243.455 ;
        RECT -62.355 236.775 -61.985 237.615 ;
        RECT -64.575 236.035 -64.275 236.720 ;
        RECT -62.330 236.475 -62.040 236.775 ;
        RECT -62.695 236.175 -62.035 236.475 ;
        RECT -64.520 231.990 -64.325 236.035 ;
        RECT -66.840 231.545 -65.730 231.845 ;
        RECT -66.895 230.705 -66.525 231.545 ;
        RECT -64.570 231.330 -64.270 231.990 ;
        RECT -64.520 219.160 -64.325 231.330 ;
        RECT -62.355 219.160 -61.985 219.705 ;
        RECT -64.520 218.965 -61.985 219.160 ;
        RECT -64.520 217.335 -64.325 218.965 ;
        RECT -62.355 218.865 -61.985 218.965 ;
        RECT -82.020 46.625 -81.340 217.335 ;
        RECT -64.850 215.860 -63.835 217.335 ;
        RECT -34.150 215.860 -32.915 242.900 ;
        RECT -70.570 211.525 -69.675 211.630 ;
        RECT -70.570 211.110 -59.935 211.525 ;
        RECT -70.570 210.990 -69.675 211.110 ;
        RECT -60.350 209.665 -59.935 211.110 ;
        RECT -60.440 208.710 -59.905 209.665 ;
        RECT -59.550 159.945 -59.295 160.435 ;
        RECT -56.550 159.945 -56.180 160.045 ;
        RECT -38.230 159.945 -37.860 160.045 ;
        RECT -35.115 159.945 -34.860 160.435 ;
        RECT -59.550 159.750 -54.015 159.945 ;
        RECT -56.550 159.205 -56.180 159.750 ;
        RECT -54.210 147.580 -54.015 159.750 ;
        RECT -39.965 159.750 -34.860 159.945 ;
        RECT -39.965 152.155 -39.770 159.750 ;
        RECT -38.230 159.205 -37.860 159.750 ;
        RECT -38.205 155.635 -37.915 155.810 ;
        RECT -38.230 154.795 -37.860 155.635 ;
        RECT -39.965 152.150 -39.155 152.155 ;
        RECT -39.965 151.780 -38.360 152.150 ;
        RECT -54.265 146.920 -53.965 147.580 ;
        RECT -52.010 147.365 -51.640 148.205 ;
        RECT -52.805 147.065 -51.695 147.365 ;
        RECT -54.210 142.875 -54.015 146.920 ;
        RECT -56.500 142.435 -55.840 142.735 ;
        RECT -56.495 142.135 -56.205 142.435 ;
        RECT -54.260 142.190 -53.960 142.875 ;
        RECT -56.550 141.295 -56.180 142.135 ;
        RECT -54.210 131.295 -54.015 142.190 ;
        RECT -42.770 133.865 -42.400 134.705 ;
        RECT -39.965 133.985 -39.770 151.780 ;
        RECT -42.715 133.805 -42.400 133.865 ;
        RECT -42.715 133.690 -41.680 133.805 ;
        RECT -42.710 133.505 -41.680 133.690 ;
        RECT -40.005 133.325 -39.705 133.985 ;
        RECT -39.965 131.295 -39.770 133.325 ;
        RECT -33.450 70.625 -33.180 71.300 ;
        RECT -33.420 70.525 -33.220 70.625 ;
        RECT -33.410 69.240 -33.230 70.525 ;
        RECT -36.305 68.955 -33.230 69.240 ;
        RECT -36.305 46.910 -35.990 68.955 ;
        RECT -33.410 68.570 -33.230 68.955 ;
        RECT -82.070 45.560 -81.180 46.625 ;
        RECT -36.340 46.405 -35.125 46.910 ;
        RECT -82.020 42.780 -81.340 45.560 ;
        RECT -10.440 5.245 -10.270 6.560 ;
        RECT -9.460 5.245 -9.290 6.560 ;
        RECT -8.480 5.245 -8.310 6.560 ;
        RECT -7.500 5.245 -7.330 6.560 ;
        RECT -6.520 5.245 -6.350 6.560 ;
        RECT -10.440 5.075 -6.350 5.245 ;
        RECT -10.440 3.790 -10.270 5.075 ;
        RECT -9.460 3.790 -9.290 5.075 ;
        RECT -8.480 3.790 -8.310 5.075 ;
        RECT -7.500 3.790 -7.330 5.075 ;
        RECT -6.520 3.790 -6.350 5.075 ;
        RECT -90.195 2.285 -88.020 2.825 ;
        RECT -32.715 2.285 -27.955 2.325 ;
        RECT -112.560 1.600 -27.955 2.285 ;
        RECT -32.715 1.495 -27.955 1.600 ;
        RECT 319.445 -19.130 319.615 -17.815 ;
        RECT 320.425 -19.130 320.595 -17.815 ;
        RECT 321.405 -19.130 321.575 -17.815 ;
        RECT 322.385 -19.130 322.555 -17.815 ;
        RECT 323.365 -19.130 323.535 -17.815 ;
        RECT 319.445 -19.300 323.535 -19.130 ;
        RECT 319.445 -20.585 319.615 -19.300 ;
        RECT 320.425 -20.585 320.595 -19.300 ;
        RECT 321.405 -20.585 321.575 -19.300 ;
        RECT 322.385 -20.585 322.555 -19.300 ;
        RECT 323.365 -20.585 323.535 -19.300 ;
        RECT -33.055 -56.370 -29.685 -55.765 ;
        RECT 306.830 -56.370 311.360 -55.580 ;
        RECT -33.055 -59.195 311.360 -56.370 ;
        RECT -33.055 -59.470 -29.685 -59.195 ;
        RECT 306.830 -59.855 311.360 -59.195 ;
      LAYER met1 ;
        RECT -70.980 294.435 -69.755 573.200 ;
        RECT -36.015 306.110 -35.725 306.505 ;
        RECT -36.015 305.840 -35.180 306.110 ;
        RECT -36.015 305.710 -35.725 305.840 ;
        RECT -35.450 304.740 -35.180 305.840 ;
        RECT -35.450 304.470 -33.460 304.740 ;
        RECT -43.065 297.555 -41.750 298.850 ;
        RECT -33.730 298.615 -33.460 304.470 ;
        RECT -33.930 297.550 -33.265 298.615 ;
        RECT -34.170 294.435 -32.700 294.610 ;
        RECT -70.980 293.710 -32.700 294.435 ;
        RECT -70.980 293.210 -32.500 293.710 ;
        RECT -41.825 277.115 -41.525 277.360 ;
        RECT -44.065 276.815 -41.525 277.115 ;
        RECT -41.825 276.675 -41.525 276.815 ;
        RECT -41.830 272.485 -41.530 272.630 ;
        RECT -41.830 272.185 -39.710 272.485 ;
        RECT -41.830 271.970 -41.530 272.185 ;
        RECT -39.905 260.115 -39.230 260.265 ;
        RECT -39.905 259.740 -38.480 260.115 ;
        RECT -39.905 259.605 -39.230 259.740 ;
        RECT -38.855 252.660 -38.480 259.740 ;
        RECT -39.045 251.765 -38.100 252.660 ;
        RECT -34.260 242.545 -32.500 293.210 ;
        RECT -64.575 236.475 -64.275 236.720 ;
        RECT -64.575 236.175 -62.035 236.475 ;
        RECT -64.575 236.035 -64.275 236.175 ;
        RECT -64.570 231.845 -64.270 231.990 ;
        RECT -66.390 231.545 -64.270 231.845 ;
        RECT -64.570 231.330 -64.270 231.545 ;
        RECT -82.020 215.860 -32.915 217.335 ;
        RECT -70.710 210.600 -69.365 215.860 ;
        RECT -60.440 209.565 -59.905 209.665 ;
        RECT -60.440 209.310 -34.860 209.565 ;
        RECT -60.440 208.710 -59.905 209.310 ;
        RECT -59.550 159.750 -59.295 209.310 ;
        RECT -35.115 159.750 -34.860 209.310 ;
        RECT -54.265 147.365 -53.965 147.580 ;
        RECT -54.265 147.065 -52.145 147.365 ;
        RECT -54.265 146.920 -53.965 147.065 ;
        RECT -54.260 142.735 -53.960 142.875 ;
        RECT -56.500 142.435 -53.960 142.735 ;
        RECT -54.260 142.190 -53.960 142.435 ;
        RECT -40.005 133.805 -39.705 133.985 ;
        RECT -42.340 133.505 -39.705 133.805 ;
        RECT -40.005 133.325 -39.705 133.505 ;
        RECT -36.340 46.845 -35.125 46.910 ;
        RECT -82.070 46.325 -81.180 46.625 ;
        RECT -36.555 46.405 -35.125 46.845 ;
        RECT -36.555 46.325 -35.400 46.405 ;
        RECT -89.180 45.645 -35.400 46.325 ;
        RECT -89.180 2.825 -88.500 45.645 ;
        RECT -82.070 45.560 -81.180 45.645 ;
        RECT -14.245 6.390 -10.235 6.610 ;
        RECT -26.215 5.890 -18.405 6.095 ;
        RECT -14.245 5.890 -14.025 6.390 ;
        RECT -26.215 5.670 -14.025 5.890 ;
        RECT -26.215 5.365 -18.405 5.670 ;
        RECT -10.470 5.540 -10.240 6.390 ;
        RECT -9.490 5.540 -9.260 6.540 ;
        RECT -8.510 5.540 -8.280 6.540 ;
        RECT -7.530 5.540 -7.300 6.540 ;
        RECT -6.550 5.540 -6.320 6.540 ;
        RECT -90.195 1.605 -88.020 2.825 ;
        RECT -26.215 2.365 -25.390 5.365 ;
        RECT -10.470 3.810 -10.240 4.810 ;
        RECT -9.490 3.810 -9.260 4.810 ;
        RECT -8.510 3.810 -8.280 4.810 ;
        RECT -7.530 3.810 -7.300 4.810 ;
        RECT -6.550 3.810 -6.320 4.810 ;
        RECT -32.995 1.945 -25.385 2.365 ;
        RECT -33.000 1.540 -25.385 1.945 ;
        RECT -33.000 1.285 -25.390 1.540 ;
        RECT -33.005 1.120 -25.390 1.285 ;
        RECT -33.005 -55.765 -31.470 1.120 ;
        RECT 315.640 -17.985 319.650 -17.765 ;
        RECT 315.640 -18.485 315.860 -17.985 ;
        RECT 308.275 -18.705 315.860 -18.485 ;
        RECT 308.275 -55.580 310.540 -18.705 ;
        RECT 319.415 -18.835 319.645 -17.985 ;
        RECT 320.395 -18.835 320.625 -17.835 ;
        RECT 321.375 -18.835 321.605 -17.835 ;
        RECT 322.355 -18.835 322.585 -17.835 ;
        RECT 323.335 -18.835 323.565 -17.835 ;
        RECT 319.415 -20.565 319.645 -19.565 ;
        RECT 320.395 -20.565 320.625 -19.565 ;
        RECT 321.375 -20.565 321.605 -19.565 ;
        RECT 322.355 -20.565 322.585 -19.565 ;
        RECT 323.335 -20.565 323.565 -19.565 ;
        RECT -33.055 -59.470 -29.685 -55.765 ;
        RECT 306.830 -59.855 311.360 -55.580 ;
    END
  END F_IN
  PIN D0
    ANTENNAGATEAREA 10.500000 ;
    PORT
      LAYER li1 ;
        RECT -119.420 -98.000 -119.115 -96.985 ;
        RECT -111.455 -98.000 -110.780 -97.935 ;
        RECT -119.420 -98.170 -110.780 -98.000 ;
        RECT -119.420 -98.175 -119.115 -98.170 ;
        RECT -111.455 -98.205 -110.780 -98.170 ;
        RECT -35.700 -99.320 -34.760 -98.950 ;
        RECT -70.730 -105.270 -70.375 -105.265 ;
        RECT -68.670 -105.270 -68.300 -105.240 ;
        RECT -70.730 -105.275 -68.300 -105.270 ;
        RECT -71.860 -105.465 -68.300 -105.275 ;
        RECT -71.860 -105.475 -70.725 -105.465 ;
        RECT -68.670 -105.595 -68.300 -105.465 ;
        RECT -71.410 -112.620 -70.760 -112.535 ;
        RECT -70.540 -112.620 -70.175 -112.555 ;
        RECT -71.410 -112.825 -70.175 -112.620 ;
        RECT -71.410 -113.285 -70.760 -112.825 ;
        RECT -70.540 -112.855 -70.175 -112.825 ;
        RECT -119.420 -125.600 -119.120 -124.695 ;
        RECT -119.420 -125.805 -109.975 -125.600 ;
        RECT -119.420 -125.880 -119.120 -125.805 ;
        RECT -110.275 -125.830 -109.975 -125.805 ;
        RECT -110.275 -126.110 -109.550 -125.830 ;
        RECT 134.195 -127.430 134.870 -127.400 ;
        RECT 134.095 -127.440 134.870 -127.430 ;
        RECT 131.455 -127.620 134.870 -127.440 ;
        RECT 152.535 -127.585 153.210 -127.555 ;
        RECT 152.435 -127.595 153.210 -127.585 ;
        RECT 39.260 -128.260 39.875 -128.255 ;
        RECT 39.255 -128.475 39.875 -128.260 ;
        RECT 39.255 -132.515 39.545 -128.475 ;
        RECT -35.320 -134.415 -34.625 -134.145 ;
        RECT -29.930 -134.385 -29.235 -134.115 ;
        RECT 39.260 -139.565 39.540 -132.515 ;
        RECT 132.370 -132.755 133.050 -127.620 ;
        RECT 134.095 -127.630 134.870 -127.620 ;
        RECT 134.195 -127.670 134.870 -127.630 ;
        RECT 150.365 -127.775 153.210 -127.595 ;
        RECT 150.365 -132.755 151.045 -127.775 ;
        RECT 152.435 -127.785 153.210 -127.775 ;
        RECT 152.535 -127.825 153.210 -127.785 ;
        RECT 132.370 -133.435 151.045 -132.755 ;
        RECT 132.370 -139.565 133.050 -133.435 ;
        RECT -162.825 -140.245 133.050 -139.565 ;
      LAYER met1 ;
        RECT -119.420 -139.620 -119.115 -96.985 ;
        RECT -35.700 -99.320 -35.020 -98.950 ;
        RECT -35.700 -101.230 -35.445 -99.320 ;
        RECT -35.700 -101.485 43.625 -101.230 ;
        RECT -71.875 -105.515 -70.890 -105.245 ;
        RECT -71.160 -110.670 -70.890 -105.515 ;
        RECT -79.215 -111.550 -70.890 -110.670 ;
        RECT -119.685 -140.235 -119.070 -139.620 ;
        RECT -79.215 -140.245 -78.335 -111.550 ;
        RECT -71.160 -112.535 -70.890 -111.550 ;
        RECT -71.410 -113.285 -70.760 -112.535 ;
        RECT 43.370 -128.235 43.625 -101.485 ;
        RECT -27.415 -128.490 43.625 -128.235 ;
        RECT -35.320 -134.230 -34.625 -134.145 ;
        RECT -29.930 -134.230 -29.235 -134.115 ;
        RECT -35.320 -134.240 -29.235 -134.230 ;
        RECT -27.415 -134.240 -27.275 -128.490 ;
        RECT -35.320 -134.370 -27.275 -134.240 ;
        RECT -35.320 -134.415 -34.625 -134.370 ;
        RECT -29.930 -134.380 -27.275 -134.370 ;
        RECT -29.930 -134.385 -29.235 -134.380 ;
    END
  END D0
  PIN D1
    ANTENNAGATEAREA 7.200000 ;
    PORT
      LAYER li1 ;
        RECT 29.680 -95.575 30.375 -95.305 ;
        RECT 35.070 -95.605 35.765 -95.335 ;
        RECT -118.465 -97.590 -118.160 -96.590 ;
        RECT -112.395 -97.590 -111.720 -97.545 ;
        RECT -118.465 -97.780 -111.720 -97.590 ;
        RECT -112.395 -97.815 -111.720 -97.780 ;
        RECT -118.465 -126.045 -118.165 -125.980 ;
        RECT -111.875 -126.045 -111.150 -125.990 ;
        RECT -118.465 -126.250 -111.150 -126.045 ;
        RECT -118.465 -127.165 -118.165 -126.250 ;
        RECT -111.875 -126.270 -111.150 -126.250 ;
        RECT 176.395 -127.485 177.070 -127.455 ;
        RECT 176.295 -127.495 177.070 -127.485 ;
        RECT 173.655 -127.675 177.070 -127.495 ;
        RECT 194.735 -127.640 195.410 -127.610 ;
        RECT 194.635 -127.650 195.410 -127.640 ;
        RECT 174.570 -132.810 175.250 -127.675 ;
        RECT 176.295 -127.685 177.070 -127.675 ;
        RECT 176.395 -127.725 177.070 -127.685 ;
        RECT 192.565 -127.830 195.410 -127.650 ;
        RECT 192.565 -132.810 193.245 -127.830 ;
        RECT 194.635 -127.840 195.410 -127.830 ;
        RECT 194.735 -127.880 195.410 -127.840 ;
        RECT 174.570 -133.490 193.245 -132.810 ;
        RECT 29.680 -134.415 30.375 -134.145 ;
        RECT 35.070 -134.385 35.765 -134.115 ;
        RECT 39.755 -134.405 40.080 -133.720 ;
        RECT 39.770 -138.205 40.040 -134.405 ;
        RECT 174.570 -140.560 175.250 -133.490 ;
        RECT -162.690 -141.240 175.250 -140.560 ;
      LAYER met1 ;
        RECT 29.680 -95.350 30.375 -95.305 ;
        RECT 35.070 -95.340 35.765 -95.335 ;
        RECT 34.560 -95.350 47.615 -95.340 ;
        RECT 29.680 -95.480 47.615 -95.350 ;
        RECT 29.680 -95.490 35.765 -95.480 ;
        RECT 29.680 -95.575 30.375 -95.490 ;
        RECT 35.070 -95.605 35.765 -95.490 ;
        RECT -118.465 -140.615 -118.160 -96.590 ;
        RECT 29.680 -134.230 30.375 -134.145 ;
        RECT 35.070 -134.230 35.765 -134.115 ;
        RECT 29.680 -134.240 35.765 -134.230 ;
        RECT 39.755 -134.240 40.080 -133.720 ;
        RECT 47.475 -134.240 47.615 -95.480 ;
        RECT 29.680 -134.370 47.615 -134.240 ;
        RECT 29.680 -134.415 30.375 -134.370 ;
        RECT 34.560 -134.380 47.615 -134.370 ;
        RECT 35.070 -134.385 35.765 -134.380 ;
        RECT 39.755 -134.405 40.080 -134.380 ;
        RECT 39.730 -140.590 40.035 -137.570 ;
        RECT -118.730 -141.230 -118.115 -140.615 ;
        RECT 39.465 -141.205 40.080 -140.590 ;
    END
  END D1
  PIN D2
    ANTENNAGATEAREA 7.200000 ;
    PORT
      LAYER li1 ;
        RECT 14.680 -95.575 15.375 -95.305 ;
        RECT 20.070 -95.605 20.765 -95.335 ;
        RECT -117.920 -97.175 -117.615 -96.160 ;
        RECT -114.075 -97.175 -113.400 -97.135 ;
        RECT -117.920 -97.350 -113.400 -97.175 ;
        RECT -114.170 -97.360 -113.400 -97.350 ;
        RECT -114.075 -97.405 -113.400 -97.360 ;
        RECT -117.915 -126.505 -117.615 -126.495 ;
        RECT -113.520 -126.505 -112.795 -126.465 ;
        RECT -117.915 -126.710 -112.795 -126.505 ;
        RECT -117.915 -127.680 -117.615 -126.710 ;
        RECT -113.520 -126.745 -112.795 -126.710 ;
        RECT 220.710 -127.680 221.385 -127.650 ;
        RECT 220.610 -127.690 221.385 -127.680 ;
        RECT 217.970 -127.870 221.385 -127.690 ;
        RECT 239.050 -127.835 239.725 -127.805 ;
        RECT 238.950 -127.845 239.725 -127.835 ;
        RECT 39.975 -131.265 40.590 -131.045 ;
        RECT 14.680 -134.415 15.375 -134.145 ;
        RECT 20.070 -134.385 20.765 -134.115 ;
        RECT 40.295 -138.205 40.565 -131.265 ;
        RECT 218.885 -132.935 219.565 -127.870 ;
        RECT 220.610 -127.880 221.385 -127.870 ;
        RECT 220.710 -127.920 221.385 -127.880 ;
        RECT 236.880 -128.025 239.725 -127.845 ;
        RECT 218.885 -133.005 219.800 -132.935 ;
        RECT 236.880 -133.005 237.560 -128.025 ;
        RECT 238.950 -128.035 239.725 -128.025 ;
        RECT 239.050 -128.075 239.725 -128.035 ;
        RECT 218.885 -133.685 237.560 -133.005 ;
        RECT 219.120 -141.725 219.800 -133.685 ;
        RECT -162.690 -142.405 219.800 -141.725 ;
      LAYER met1 ;
        RECT 14.680 -95.350 15.375 -95.305 ;
        RECT 20.070 -95.340 20.765 -95.335 ;
        RECT 20.070 -95.350 26.865 -95.340 ;
        RECT 14.680 -95.480 26.865 -95.350 ;
        RECT 14.680 -95.490 20.765 -95.480 ;
        RECT 14.680 -95.575 15.375 -95.490 ;
        RECT 20.070 -95.605 20.765 -95.490 ;
        RECT -117.920 -97.350 -117.615 -96.160 ;
        RECT -117.920 -126.495 -117.620 -97.350 ;
        RECT 26.725 -98.470 26.865 -95.480 ;
        RECT 26.725 -98.610 46.860 -98.470 ;
        RECT -117.920 -127.680 -117.615 -126.495 ;
        RECT -117.920 -141.780 -117.620 -127.680 ;
        RECT 39.930 -131.110 40.625 -131.035 ;
        RECT 46.720 -131.110 46.860 -98.610 ;
        RECT 26.725 -131.250 46.860 -131.110 ;
        RECT 14.680 -134.230 15.375 -134.145 ;
        RECT 20.070 -134.230 20.765 -134.115 ;
        RECT 14.680 -134.240 20.765 -134.230 ;
        RECT 26.725 -134.240 26.865 -131.250 ;
        RECT 39.930 -131.270 40.625 -131.250 ;
        RECT 14.680 -134.370 26.865 -134.240 ;
        RECT 14.680 -134.415 15.375 -134.370 ;
        RECT 20.070 -134.380 26.865 -134.370 ;
        RECT 20.070 -134.385 20.765 -134.380 ;
        RECT 40.320 -137.590 40.540 -137.575 ;
        RECT 40.275 -141.755 40.575 -137.590 ;
        RECT -118.200 -142.395 -117.585 -141.780 ;
        RECT 39.995 -142.370 40.610 -141.755 ;
    END
  END D2
  PIN D3
    ANTENNAGATEAREA 7.000000 ;
    PORT
      LAYER li1 ;
        RECT -104.795 -98.775 -104.110 -98.755 ;
        RECT -104.985 -98.785 -103.850 -98.775 ;
        RECT -101.795 -98.785 -101.425 -98.655 ;
        RECT -104.985 -98.975 -101.425 -98.785 ;
        RECT -104.795 -99.045 -104.110 -98.975 ;
        RECT -103.855 -98.980 -101.425 -98.975 ;
        RECT -103.855 -98.985 -103.500 -98.980 ;
        RECT -101.795 -99.010 -101.425 -98.980 ;
        RECT -117.425 -102.370 -117.125 -101.990 ;
        RECT -117.425 -102.570 -117.085 -102.370 ;
        RECT -117.425 -102.955 -117.125 -102.570 ;
        RECT -105.340 -102.955 -104.680 -102.910 ;
        RECT -117.425 -103.155 -104.680 -102.955 ;
        RECT -117.425 -103.175 -117.125 -103.155 ;
        RECT -105.340 -103.175 -104.680 -103.155 ;
        RECT 29.730 -106.830 30.425 -106.560 ;
        RECT 35.120 -106.860 35.815 -106.590 ;
        RECT 29.730 -123.160 30.425 -122.890 ;
        RECT 35.120 -123.130 35.815 -122.860 ;
        RECT 40.675 -123.185 41.400 -122.510 ;
        RECT -107.950 -124.290 -107.660 -123.815 ;
        RECT -105.915 -124.290 -105.200 -124.255 ;
        RECT -107.950 -124.470 -105.200 -124.290 ;
        RECT -107.950 -124.500 -107.660 -124.470 ;
        RECT -105.915 -124.555 -105.200 -124.470 ;
        RECT -117.425 -129.525 -117.135 -129.045 ;
        RECT -108.050 -129.525 -107.760 -129.045 ;
        RECT -117.425 -129.730 -107.760 -129.525 ;
        RECT 40.790 -139.290 41.070 -123.185 ;
        RECT 266.700 -127.510 267.375 -127.480 ;
        RECT 266.600 -127.520 267.375 -127.510 ;
        RECT 263.960 -127.700 267.375 -127.520 ;
        RECT 285.040 -127.665 285.715 -127.635 ;
        RECT 284.940 -127.675 285.715 -127.665 ;
        RECT 264.875 -132.835 265.555 -127.700 ;
        RECT 266.600 -127.710 267.375 -127.700 ;
        RECT 266.700 -127.750 267.375 -127.710 ;
        RECT 282.870 -127.855 285.715 -127.675 ;
        RECT 282.870 -132.835 283.550 -127.855 ;
        RECT 284.940 -127.865 285.715 -127.855 ;
        RECT 285.040 -127.905 285.715 -127.865 ;
        RECT 264.875 -133.515 283.550 -132.835 ;
        RECT 264.875 -143.000 265.555 -133.515 ;
        RECT -162.960 -143.680 265.555 -143.000 ;
      LAYER met1 ;
        RECT -104.795 -99.045 -104.110 -98.755 ;
        RECT -117.425 -143.065 -117.120 -101.985 ;
        RECT -104.760 -102.910 -104.560 -99.045 ;
        RECT -105.340 -102.955 -104.560 -102.910 ;
        RECT -105.575 -103.155 -104.560 -102.955 ;
        RECT -105.340 -103.175 -104.680 -103.155 ;
        RECT 29.730 -106.605 30.425 -106.560 ;
        RECT 35.120 -106.595 35.815 -106.590 ;
        RECT 41.770 -106.595 42.025 -106.555 ;
        RECT 35.120 -106.605 42.025 -106.595 ;
        RECT 29.730 -106.735 42.025 -106.605 ;
        RECT 29.730 -106.745 35.815 -106.735 ;
        RECT 29.730 -106.830 30.425 -106.745 ;
        RECT 35.120 -106.860 35.815 -106.745 ;
        RECT 41.770 -106.810 42.025 -106.735 ;
        RECT 29.730 -122.975 30.425 -122.890 ;
        RECT 35.120 -122.975 35.815 -122.860 ;
        RECT 29.730 -122.985 35.815 -122.975 ;
        RECT 40.675 -122.985 41.400 -122.510 ;
        RECT 41.835 -122.985 41.975 -106.810 ;
        RECT 29.730 -123.115 41.985 -122.985 ;
        RECT 29.730 -123.160 30.425 -123.115 ;
        RECT 35.120 -123.125 41.985 -123.115 ;
        RECT 35.120 -123.130 35.815 -123.125 ;
        RECT 40.675 -123.185 41.400 -123.125 ;
        RECT -107.950 -124.500 -107.660 -123.815 ;
        RECT -107.950 -129.045 -107.775 -124.500 ;
        RECT -108.050 -129.730 -107.760 -129.045 ;
        RECT 40.770 -143.040 41.075 -138.305 ;
        RECT -117.735 -143.680 -117.115 -143.065 ;
        RECT 40.460 -143.655 41.080 -143.040 ;
    END
  END D3
  PIN D4
    ANTENNAGATEAREA 7.000000 ;
    PORT
      LAYER li1 ;
        RECT 2.180 -95.575 2.875 -95.305 ;
        RECT 7.570 -95.605 8.265 -95.335 ;
        RECT -105.270 -98.305 -104.585 -98.220 ;
        RECT -104.120 -98.295 -103.445 -98.265 ;
        RECT -104.220 -98.305 -103.445 -98.295 ;
        RECT -105.270 -98.485 -103.445 -98.305 ;
        RECT -105.270 -98.510 -104.585 -98.485 ;
        RECT -104.220 -98.495 -103.445 -98.485 ;
        RECT -104.120 -98.535 -103.445 -98.495 ;
        RECT -116.860 -102.540 -116.555 -101.650 ;
        RECT -105.420 -102.540 -105.155 -102.060 ;
        RECT -116.860 -102.720 -105.155 -102.540 ;
        RECT -116.860 -102.730 -116.555 -102.720 ;
        RECT -107.575 -124.735 -107.285 -124.670 ;
        RECT -107.030 -124.735 -106.300 -124.655 ;
        RECT -107.575 -124.915 -106.300 -124.735 ;
        RECT -107.575 -125.355 -107.285 -124.915 ;
        RECT -107.030 -124.955 -106.300 -124.915 ;
        RECT 310.470 -127.180 311.145 -127.150 ;
        RECT 310.370 -127.190 311.145 -127.180 ;
        RECT 307.730 -127.370 311.145 -127.190 ;
        RECT 328.810 -127.335 329.485 -127.305 ;
        RECT 328.710 -127.345 329.485 -127.335 ;
        RECT -116.860 -129.920 -116.570 -129.905 ;
        RECT -107.585 -129.920 -107.295 -129.440 ;
        RECT -116.860 -130.125 -107.295 -129.920 ;
        RECT -116.860 -130.590 -116.570 -130.125 ;
        RECT 41.350 -130.550 42.135 -130.350 ;
        RECT 2.180 -134.415 2.875 -134.145 ;
        RECT 7.570 -134.385 8.265 -134.115 ;
        RECT 41.350 -138.205 41.620 -130.550 ;
        RECT 308.645 -132.505 309.325 -127.370 ;
        RECT 310.370 -127.380 311.145 -127.370 ;
        RECT 310.470 -127.420 311.145 -127.380 ;
        RECT 326.640 -127.525 329.485 -127.345 ;
        RECT 326.640 -132.505 327.320 -127.525 ;
        RECT 328.710 -127.535 329.485 -127.525 ;
        RECT 328.810 -127.575 329.485 -127.535 ;
        RECT 308.645 -133.185 327.320 -132.505 ;
        RECT 41.445 -144.430 42.125 -144.420 ;
        RECT 308.645 -144.430 309.325 -133.185 ;
        RECT -165.005 -145.110 309.325 -144.430 ;
        RECT -165.005 -145.135 -114.705 -145.110 ;
      LAYER met1 ;
        RECT 2.180 -95.350 2.875 -95.305 ;
        RECT 7.570 -95.340 8.265 -95.335 ;
        RECT 7.570 -95.350 10.260 -95.340 ;
        RECT 2.180 -95.480 10.260 -95.350 ;
        RECT 2.180 -95.490 8.265 -95.480 ;
        RECT 2.180 -95.575 2.875 -95.490 ;
        RECT 7.570 -95.605 8.265 -95.490 ;
        RECT -105.270 -98.305 -104.585 -98.220 ;
        RECT -105.410 -98.510 -104.585 -98.305 ;
        RECT -116.860 -144.485 -116.555 -101.650 ;
        RECT -105.410 -102.060 -105.230 -98.510 ;
        RECT 10.120 -99.205 10.260 -95.480 ;
        RECT 10.120 -99.345 46.065 -99.205 ;
        RECT -105.420 -102.720 -105.155 -102.060 ;
        RECT -107.575 -124.690 -107.285 -124.670 ;
        RECT -107.580 -125.355 -107.285 -124.690 ;
        RECT -107.580 -129.440 -107.365 -125.355 ;
        RECT -107.585 -130.125 -107.295 -129.440 ;
        RECT 41.495 -130.375 42.215 -130.340 ;
        RECT 45.925 -130.375 46.065 -99.345 ;
        RECT 10.120 -130.515 46.065 -130.375 ;
        RECT 2.180 -134.230 2.875 -134.145 ;
        RECT 7.570 -134.230 8.265 -134.115 ;
        RECT 2.180 -134.240 8.265 -134.230 ;
        RECT 10.120 -134.240 10.260 -130.515 ;
        RECT 41.495 -130.575 42.215 -130.515 ;
        RECT 2.180 -134.370 10.260 -134.240 ;
        RECT 2.180 -134.415 2.875 -134.370 ;
        RECT 7.570 -134.380 10.260 -134.370 ;
        RECT 7.570 -134.385 8.265 -134.380 ;
        RECT 41.335 -144.460 41.640 -137.575 ;
        RECT -117.205 -144.490 -116.555 -144.485 ;
        RECT 40.990 -144.465 41.640 -144.460 ;
        RECT -117.205 -144.655 -116.550 -144.490 ;
        RECT 40.990 -144.630 41.645 -144.465 ;
        RECT -117.200 -145.080 -116.550 -144.655 ;
        RECT 40.995 -145.055 41.645 -144.630 ;
    END
  END D4
  PIN D5
    ANTENNAGATEAREA 7.000000 ;
    PORT
      LAYER li1 ;
        RECT -10.320 -95.575 -9.625 -95.305 ;
        RECT -4.930 -95.605 -4.235 -95.335 ;
        RECT -116.195 -108.330 -113.560 -108.320 ;
        RECT -111.505 -108.330 -111.135 -108.200 ;
        RECT -116.195 -108.520 -111.135 -108.330 ;
        RECT -116.195 -109.045 -115.995 -108.520 ;
        RECT -113.565 -108.525 -111.135 -108.520 ;
        RECT -113.565 -108.530 -113.210 -108.525 ;
        RECT -111.505 -108.555 -111.135 -108.525 ;
        RECT -116.280 -110.230 -115.980 -109.045 ;
        RECT -103.370 -124.295 -103.080 -123.820 ;
        RECT -101.390 -124.295 -100.675 -124.260 ;
        RECT -103.370 -124.475 -100.675 -124.295 ;
        RECT -103.370 -124.505 -103.080 -124.475 ;
        RECT -101.390 -124.560 -100.675 -124.475 ;
        RECT 356.235 -127.095 356.910 -127.065 ;
        RECT 356.135 -127.105 356.910 -127.095 ;
        RECT 353.495 -127.285 356.910 -127.105 ;
        RECT 374.575 -127.250 375.250 -127.220 ;
        RECT 374.475 -127.260 375.250 -127.250 ;
        RECT -116.290 -130.315 -116.000 -130.310 ;
        RECT -103.480 -130.315 -103.190 -129.835 ;
        RECT 42.145 -129.915 42.760 -129.695 ;
        RECT -116.290 -130.520 -103.190 -130.315 ;
        RECT -116.290 -130.995 -116.000 -130.520 ;
        RECT 42.420 -132.070 42.690 -129.915 ;
        RECT 41.925 -132.340 42.690 -132.070 ;
        RECT -10.320 -134.415 -9.625 -134.145 ;
        RECT -4.930 -134.385 -4.235 -134.115 ;
        RECT 41.925 -138.205 42.195 -132.340 ;
        RECT 354.410 -132.420 355.090 -127.285 ;
        RECT 356.135 -127.295 356.910 -127.285 ;
        RECT 356.235 -127.335 356.910 -127.295 ;
        RECT 372.405 -127.440 375.250 -127.260 ;
        RECT 372.405 -132.420 373.085 -127.440 ;
        RECT 374.475 -127.450 375.250 -127.440 ;
        RECT 374.575 -127.490 375.250 -127.450 ;
        RECT 354.410 -133.100 373.085 -132.420 ;
        RECT 354.410 -145.925 355.090 -133.100 ;
        RECT -163.775 -146.605 355.090 -145.925 ;
      LAYER met1 ;
        RECT -10.320 -95.350 -9.625 -95.305 ;
        RECT -4.930 -95.340 -4.235 -95.335 ;
        RECT -4.930 -95.350 -2.070 -95.340 ;
        RECT -10.320 -95.480 -2.070 -95.350 ;
        RECT -10.320 -95.490 -4.235 -95.480 ;
        RECT -10.320 -95.575 -9.625 -95.490 ;
        RECT -4.930 -95.605 -4.235 -95.490 ;
        RECT -2.210 -99.805 -2.070 -95.480 ;
        RECT -2.210 -99.945 45.255 -99.805 ;
        RECT -116.290 -145.125 -115.970 -109.010 ;
        RECT -103.370 -124.505 -103.080 -123.820 ;
        RECT -103.370 -129.835 -103.195 -124.505 ;
        RECT 42.125 -129.775 42.840 -129.685 ;
        RECT 45.115 -129.775 45.255 -99.945 ;
        RECT -103.480 -130.520 -103.190 -129.835 ;
        RECT -2.210 -129.915 45.255 -129.775 ;
        RECT -10.320 -134.230 -9.625 -134.145 ;
        RECT -4.930 -134.230 -4.235 -134.115 ;
        RECT -10.320 -134.240 -4.235 -134.230 ;
        RECT -2.210 -134.240 -2.070 -129.915 ;
        RECT 42.125 -129.920 42.840 -129.915 ;
        RECT -10.320 -134.370 -2.070 -134.240 ;
        RECT -10.320 -134.415 -9.625 -134.370 ;
        RECT -4.930 -134.380 -2.070 -134.370 ;
        RECT -4.930 -134.385 -4.235 -134.380 ;
        RECT 41.905 -145.100 42.225 -137.555 ;
        RECT -116.300 -145.985 -115.970 -145.125 ;
        RECT 41.895 -145.960 42.225 -145.100 ;
        RECT -116.405 -145.990 -115.970 -145.985 ;
        RECT 41.790 -145.965 42.225 -145.960 ;
        RECT -116.405 -146.605 -115.790 -145.990 ;
        RECT 41.790 -146.580 42.405 -145.965 ;
    END
  END D5
  PIN D6
    ANTENNAGATEAREA 7.000000 ;
    PORT
      LAYER li1 ;
        RECT -22.820 -95.575 -22.125 -95.305 ;
        RECT -17.430 -95.605 -16.735 -95.335 ;
        RECT -115.565 -107.850 -115.265 -106.855 ;
        RECT -113.830 -107.840 -113.155 -107.810 ;
        RECT -113.930 -107.850 -113.155 -107.840 ;
        RECT -115.565 -108.030 -113.155 -107.850 ;
        RECT -115.565 -108.040 -115.265 -108.030 ;
        RECT -113.930 -108.040 -113.155 -108.030 ;
        RECT -113.830 -108.080 -113.155 -108.040 ;
        RECT -102.985 -124.740 -102.695 -124.680 ;
        RECT -102.505 -124.740 -101.775 -124.660 ;
        RECT -102.985 -124.920 -101.775 -124.740 ;
        RECT -102.985 -125.365 -102.695 -124.920 ;
        RECT -102.505 -124.960 -101.775 -124.920 ;
        RECT 403.055 -126.905 403.730 -126.875 ;
        RECT 402.955 -126.915 403.730 -126.905 ;
        RECT 400.315 -127.095 403.730 -126.915 ;
        RECT 421.395 -127.060 422.070 -127.030 ;
        RECT 421.295 -127.070 422.070 -127.060 ;
        RECT 42.925 -129.240 43.665 -129.000 ;
        RECT -103.015 -130.700 -102.725 -130.220 ;
        RECT -115.565 -130.905 -102.725 -130.700 ;
        RECT -115.565 -131.385 -115.275 -130.905 ;
        RECT -22.820 -134.415 -22.125 -134.145 ;
        RECT -17.430 -134.385 -16.735 -134.115 ;
        RECT 42.645 -137.730 42.915 -137.580 ;
        RECT 43.135 -137.730 43.405 -129.240 ;
        RECT 401.230 -132.230 401.910 -127.095 ;
        RECT 402.955 -127.105 403.730 -127.095 ;
        RECT 403.055 -127.145 403.730 -127.105 ;
        RECT 419.225 -127.250 422.070 -127.070 ;
        RECT 419.225 -132.230 419.905 -127.250 ;
        RECT 421.295 -127.260 422.070 -127.250 ;
        RECT 421.395 -127.300 422.070 -127.260 ;
        RECT 401.230 -132.910 419.905 -132.230 ;
        RECT 42.645 -138.000 43.405 -137.730 ;
        RECT 42.645 -138.205 42.915 -138.000 ;
        RECT 401.350 -147.775 402.030 -132.910 ;
        RECT -164.585 -148.455 402.030 -147.775 ;
      LAYER met1 ;
        RECT -22.820 -95.350 -22.125 -95.305 ;
        RECT -17.430 -95.340 -16.735 -95.335 ;
        RECT -17.430 -95.350 -14.490 -95.340 ;
        RECT -22.820 -95.480 -14.490 -95.350 ;
        RECT -22.820 -95.490 -16.735 -95.480 ;
        RECT -22.820 -95.575 -22.125 -95.490 ;
        RECT -17.430 -95.605 -16.735 -95.490 ;
        RECT -14.630 -100.500 -14.490 -95.480 ;
        RECT -14.630 -100.680 44.460 -100.500 ;
        RECT -115.565 -147.825 -115.265 -106.855 ;
        RECT -102.985 -125.365 -102.695 -124.680 ;
        RECT -102.985 -130.220 -102.810 -125.365 ;
        RECT 42.925 -129.040 43.665 -129.000 ;
        RECT 44.280 -129.040 44.460 -100.680 ;
        RECT -14.630 -129.220 44.460 -129.040 ;
        RECT -103.015 -130.905 -102.725 -130.220 ;
        RECT -22.820 -134.230 -22.125 -134.145 ;
        RECT -17.430 -134.230 -16.735 -134.115 ;
        RECT -22.820 -134.240 -16.735 -134.230 ;
        RECT -14.630 -134.240 -14.490 -129.220 ;
        RECT 42.925 -129.240 43.665 -129.220 ;
        RECT -22.820 -134.370 -14.490 -134.240 ;
        RECT -22.820 -134.415 -22.125 -134.370 ;
        RECT -17.430 -134.380 -14.490 -134.370 ;
        RECT -17.430 -134.385 -16.735 -134.380 ;
        RECT 42.630 -147.800 42.930 -137.375 ;
        RECT -115.650 -148.440 -115.035 -147.825 ;
        RECT 42.545 -148.415 43.160 -147.800 ;
    END
  END D6
  PIN D7
    ANTENNAGATEAREA 10.500000 ;
    PORT
      LAYER li1 ;
        RECT -60.170 319.100 -59.900 319.775 ;
        RECT -60.130 319.000 -59.930 319.100 ;
        RECT -60.120 317.610 -59.940 319.000 ;
        RECT -65.780 316.930 -59.940 317.610 ;
        RECT -65.780 299.615 -65.100 316.930 ;
        RECT -60.015 300.760 -59.745 301.435 ;
        RECT -59.975 300.660 -59.775 300.760 ;
        RECT -59.965 299.615 -59.785 300.660 ;
        RECT -72.590 298.935 -59.785 299.615 ;
        RECT -72.590 206.105 -71.910 298.935 ;
        RECT -59.965 298.020 -59.785 298.935 ;
        RECT -60.820 206.110 -60.600 206.440 ;
        RECT -64.860 206.105 -60.600 206.110 ;
        RECT -72.590 205.825 -60.600 206.105 ;
        RECT -72.590 22.360 -71.910 205.825 ;
        RECT -64.860 205.820 -60.605 205.825 ;
        RECT -66.730 136.635 -66.460 137.330 ;
        RECT -66.760 131.245 -66.490 131.940 ;
        RECT -31.665 130.865 -31.295 131.805 ;
        RECT -37.940 97.895 -37.585 98.265 ;
        RECT -45.200 96.025 -44.900 96.390 ;
        RECT -37.810 96.190 -37.615 97.895 ;
        RECT -45.170 95.805 -44.965 96.025 ;
        RECT -37.810 95.840 -37.610 96.190 ;
        RECT -37.820 95.835 -37.610 95.840 ;
        RECT -45.630 95.155 -44.880 95.805 ;
        RECT -37.820 94.705 -37.620 95.835 ;
        RECT -58.455 56.590 -58.175 57.015 ;
        RECT -58.455 56.290 -57.945 56.590 ;
        RECT -58.150 47.445 -57.945 56.290 ;
        RECT -30.550 55.110 -30.280 55.785 ;
        RECT -30.515 47.450 -30.345 55.110 ;
        RECT -58.225 47.145 -57.040 47.445 ;
        RECT -30.520 47.145 -29.330 47.450 ;
        RECT -102.580 21.680 -71.910 22.360 ;
      LAYER met1 ;
        RECT -60.835 209.935 -33.575 210.190 ;
        RECT -60.835 139.290 -60.580 209.935 ;
        RECT -66.725 139.150 -60.580 139.290 ;
        RECT -66.725 137.330 -66.585 139.150 ;
        RECT -66.730 136.635 -66.460 137.330 ;
        RECT -66.715 131.940 -66.575 136.635 ;
        RECT -66.760 131.245 -66.490 131.940 ;
        RECT -33.830 131.120 -33.575 209.935 ;
        RECT -31.665 131.120 -31.295 131.545 ;
        RECT -33.830 130.865 -31.295 131.120 ;
        RECT -45.630 95.675 -44.880 95.805 ;
        RECT -45.630 95.405 -37.590 95.675 ;
        RECT -45.630 95.155 -44.880 95.405 ;
        RECT -43.895 88.230 -43.015 95.405 ;
        RECT -37.860 94.690 -37.590 95.405 ;
        RECT -72.590 87.350 -43.015 88.230 ;
        RECT -72.580 47.450 -71.965 47.495 ;
        RECT -72.580 47.145 -29.330 47.450 ;
        RECT -72.580 46.880 -71.965 47.145 ;
    END
  END D7
  PIN D8
    ANTENNAGATEAREA 7.200000 ;
    PORT
      LAYER li1 ;
        RECT -60.225 361.300 -59.955 361.975 ;
        RECT -60.185 361.200 -59.985 361.300 ;
        RECT -60.175 359.810 -59.995 361.200 ;
        RECT -65.835 359.130 -59.995 359.810 ;
        RECT -65.835 341.815 -65.155 359.130 ;
        RECT -60.070 342.960 -59.800 343.635 ;
        RECT -60.030 342.860 -59.830 342.960 ;
        RECT -60.020 341.815 -59.840 342.860 ;
        RECT -73.585 341.135 -59.840 341.815 ;
        RECT -73.585 27.445 -72.905 341.135 ;
        RECT -60.020 340.220 -59.840 341.135 ;
        RECT -66.750 206.605 -66.065 206.645 ;
        RECT -70.550 206.335 -66.065 206.605 ;
        RECT -66.750 206.320 -66.065 206.335 ;
        RECT -66.730 201.635 -66.460 202.330 ;
        RECT -27.950 201.635 -27.680 202.330 ;
        RECT -66.760 196.245 -66.490 196.940 ;
        RECT -27.920 196.245 -27.650 196.940 ;
        RECT -58.615 54.690 -58.335 55.415 ;
        RECT -58.595 48.400 -58.390 54.690 ;
        RECT -30.160 54.170 -29.890 54.845 ;
        RECT -30.125 48.405 -29.935 54.170 ;
        RECT -59.510 48.100 -58.325 48.400 ;
        RECT -30.125 48.100 -28.935 48.405 ;
        RECT -99.900 26.765 -72.905 27.445 ;
        RECT -73.585 26.550 -72.905 26.765 ;
      LAYER met1 ;
        RECT -66.725 214.040 -27.685 214.180 ;
        RECT -66.725 206.645 -66.585 214.040 ;
        RECT -73.550 206.600 -72.935 206.645 ;
        RECT -73.550 206.295 -69.915 206.600 ;
        RECT -66.750 206.320 -66.065 206.645 ;
        RECT -73.550 206.030 -72.935 206.295 ;
        RECT -66.725 202.330 -66.585 206.320 ;
        RECT -27.825 202.330 -27.685 214.040 ;
        RECT -66.730 201.635 -66.460 202.330 ;
        RECT -27.950 201.635 -27.680 202.330 ;
        RECT -66.725 201.125 -66.575 201.635 ;
        RECT -66.715 196.940 -66.575 201.125 ;
        RECT -27.835 201.125 -27.685 201.635 ;
        RECT -27.835 196.940 -27.695 201.125 ;
        RECT -66.760 196.245 -66.490 196.940 ;
        RECT -27.920 196.245 -27.650 196.940 ;
        RECT -73.575 48.405 -72.960 48.450 ;
        RECT -73.575 48.100 -28.935 48.405 ;
        RECT -73.575 47.835 -72.960 48.100 ;
    END
  END D8
  PIN D9
    ANTENNAGATEAREA 7.200000 ;
    PORT
      LAYER li1 ;
        RECT -60.420 405.615 -60.150 406.290 ;
        RECT -60.380 405.515 -60.180 405.615 ;
        RECT -60.370 404.125 -60.190 405.515 ;
        RECT -66.030 403.445 -60.190 404.125 ;
        RECT -66.030 386.365 -65.350 403.445 ;
        RECT -60.265 387.275 -59.995 387.950 ;
        RECT -60.225 387.175 -60.025 387.275 ;
        RECT -74.750 386.130 -65.280 386.365 ;
        RECT -60.215 386.130 -60.035 387.175 ;
        RECT -74.750 385.685 -60.035 386.130 ;
        RECT -74.750 35.765 -74.070 385.685 ;
        RECT -66.030 385.450 -60.035 385.685 ;
        RECT -60.215 384.535 -60.035 385.450 ;
        RECT -63.610 207.130 -63.390 207.155 ;
        RECT -70.550 206.860 -63.390 207.130 ;
        RECT -63.610 206.540 -63.390 206.860 ;
        RECT -66.730 186.635 -66.460 187.330 ;
        RECT -27.950 186.635 -27.680 187.330 ;
        RECT -66.760 181.245 -66.490 181.940 ;
        RECT -27.920 181.245 -27.650 181.940 ;
        RECT -59.090 53.045 -58.810 53.770 ;
        RECT -59.055 48.950 -58.850 53.045 ;
        RECT -29.750 52.490 -29.480 53.165 ;
        RECT -29.705 52.395 -29.520 52.490 ;
        RECT -29.695 48.950 -29.520 52.395 ;
        RECT -60.025 48.650 -58.840 48.950 ;
        RECT -29.695 48.645 -28.505 48.950 ;
        RECT -99.255 35.085 -74.070 35.765 ;
      LAYER met1 ;
        RECT -63.595 213.285 -30.815 213.425 ;
        RECT -63.595 207.190 -63.455 213.285 ;
        RECT -74.715 207.140 -74.100 207.175 ;
        RECT -74.715 207.105 -69.935 207.140 ;
        RECT -74.715 206.885 -69.920 207.105 ;
        RECT -74.715 206.840 -69.935 206.885 ;
        RECT -74.715 206.560 -74.100 206.840 ;
        RECT -63.615 206.495 -63.380 207.190 ;
        RECT -63.595 193.430 -63.455 206.495 ;
        RECT -66.725 193.290 -63.455 193.430 ;
        RECT -30.955 193.430 -30.815 213.285 ;
        RECT -30.955 193.290 -27.685 193.430 ;
        RECT -66.725 187.330 -66.585 193.290 ;
        RECT -27.825 187.330 -27.685 193.290 ;
        RECT -66.730 186.635 -66.460 187.330 ;
        RECT -27.950 186.635 -27.680 187.330 ;
        RECT -66.715 181.940 -66.575 186.635 ;
        RECT -27.835 181.940 -27.695 186.635 ;
        RECT -66.760 181.245 -66.490 181.940 ;
        RECT -27.920 181.245 -27.650 181.940 ;
        RECT -74.740 48.945 -74.125 48.980 ;
        RECT -60.025 48.945 -58.840 48.950 ;
        RECT -29.695 48.945 -28.505 48.950 ;
        RECT -74.740 48.645 -28.505 48.945 ;
        RECT -74.740 48.365 -74.125 48.645 ;
    END
  END D9
  PIN D10
    ANTENNAGATEAREA 7.000000 ;
    PORT
      LAYER li1 ;
        RECT -60.250 451.605 -59.980 452.280 ;
        RECT -60.210 451.505 -60.010 451.605 ;
        RECT -60.200 450.115 -60.020 451.505 ;
        RECT -65.860 449.435 -60.020 450.115 ;
        RECT -65.860 432.120 -65.180 449.435 ;
        RECT -60.095 433.265 -59.825 433.940 ;
        RECT -60.055 433.165 -59.855 433.265 ;
        RECT -60.045 432.120 -59.865 433.165 ;
        RECT -76.025 431.440 -59.865 432.120 ;
        RECT -76.025 39.280 -75.345 431.440 ;
        RECT -60.045 430.525 -59.865 431.440 ;
        RECT -55.530 207.635 -54.855 207.965 ;
        RECT -71.635 207.355 -54.855 207.635 ;
        RECT -55.530 207.240 -54.855 207.355 ;
        RECT -55.475 201.685 -55.205 202.380 ;
        RECT -39.205 201.685 -38.935 202.380 ;
        RECT -55.505 196.295 -55.235 196.990 ;
        RECT -39.175 196.295 -38.905 196.990 ;
        RECT -31.355 64.770 -31.000 65.140 ;
        RECT -31.325 63.065 -31.130 64.770 ;
        RECT -31.330 62.715 -31.130 63.065 ;
        RECT -31.330 62.710 -31.120 62.715 ;
        RECT -31.320 62.455 -31.120 62.710 ;
        RECT -56.900 60.650 -56.600 61.365 ;
        RECT -35.520 61.225 -35.255 61.885 ;
        RECT -31.390 61.770 -31.100 62.455 ;
        RECT -31.320 61.580 -31.120 61.770 ;
        RECT -56.815 58.905 -56.635 60.650 ;
        RECT -62.075 58.515 -61.390 58.805 ;
        RECT -56.845 58.615 -56.160 58.905 ;
        RECT -62.075 49.430 -61.870 58.515 ;
        RECT -35.500 49.440 -35.300 61.225 ;
        RECT -34.915 49.440 -34.715 49.480 ;
        RECT -62.075 49.140 -61.390 49.430 ;
        RECT -35.520 49.140 -34.335 49.440 ;
        RECT -95.000 38.600 -75.345 39.280 ;
      LAYER met1 ;
        RECT -55.470 208.540 -55.330 208.550 ;
        RECT -39.155 208.540 -38.900 208.590 ;
        RECT -55.470 208.400 -38.900 208.540 ;
        RECT -55.470 207.965 -55.330 208.400 ;
        RECT -39.155 208.335 -38.900 208.400 ;
        RECT -76.000 207.640 -75.385 207.645 ;
        RECT -76.000 207.335 -70.650 207.640 ;
        RECT -76.000 207.025 -75.385 207.335 ;
        RECT -55.530 207.240 -54.855 207.965 ;
        RECT -55.470 202.380 -55.330 207.240 ;
        RECT -39.080 202.380 -38.940 208.335 ;
        RECT -55.475 201.685 -55.205 202.380 ;
        RECT -39.205 201.685 -38.935 202.380 ;
        RECT -55.460 196.990 -55.320 201.685 ;
        RECT -39.090 196.990 -38.950 201.685 ;
        RECT -55.505 196.295 -55.235 196.990 ;
        RECT -39.175 196.295 -38.905 196.990 ;
        RECT -31.390 62.005 -31.100 62.455 ;
        RECT -35.500 61.885 -31.100 62.005 ;
        RECT -35.520 61.805 -31.100 61.885 ;
        RECT -35.520 61.225 -35.255 61.805 ;
        RECT -31.390 61.770 -31.100 61.805 ;
        RECT -35.500 60.990 -35.300 61.225 ;
        RECT -62.075 58.790 -61.390 58.805 ;
        RECT -56.845 58.790 -56.160 58.905 ;
        RECT -62.075 58.615 -56.160 58.790 ;
        RECT -62.075 58.515 -61.390 58.615 ;
        RECT -76.025 49.445 -75.410 49.450 ;
        RECT -76.025 49.140 -34.330 49.445 ;
        RECT -76.025 48.830 -75.410 49.140 ;
    END
  END D10
  PIN D16
    ANTENNAGATEAREA 10.500000 ;
    PORT
      LAYER li1 ;
        RECT -112.415 -271.510 -112.110 -270.495 ;
        RECT -104.450 -271.510 -103.775 -271.445 ;
        RECT -112.415 -271.680 -103.775 -271.510 ;
        RECT -112.415 -271.685 -112.110 -271.680 ;
        RECT -104.450 -271.715 -103.775 -271.680 ;
        RECT -28.695 -272.830 -27.755 -272.460 ;
        RECT -63.725 -278.780 -63.370 -278.775 ;
        RECT -61.665 -278.780 -61.295 -278.750 ;
        RECT -63.725 -278.785 -61.295 -278.780 ;
        RECT -64.855 -278.975 -61.295 -278.785 ;
        RECT -64.855 -278.985 -63.720 -278.975 ;
        RECT -61.665 -279.105 -61.295 -278.975 ;
        RECT -64.405 -286.130 -63.755 -286.045 ;
        RECT -63.535 -286.130 -63.170 -286.065 ;
        RECT -64.405 -286.335 -63.170 -286.130 ;
        RECT -64.405 -286.795 -63.755 -286.335 ;
        RECT -63.535 -286.365 -63.170 -286.335 ;
        RECT -112.415 -299.110 -112.115 -298.205 ;
        RECT -112.415 -299.315 -102.970 -299.110 ;
        RECT -112.415 -299.390 -112.115 -299.315 ;
        RECT -103.270 -299.340 -102.970 -299.315 ;
        RECT -103.270 -299.620 -102.545 -299.340 ;
        RECT 141.200 -300.940 141.875 -300.910 ;
        RECT 141.100 -300.950 141.875 -300.940 ;
        RECT 138.460 -301.130 141.875 -300.950 ;
        RECT 159.540 -301.095 160.215 -301.065 ;
        RECT 159.440 -301.105 160.215 -301.095 ;
        RECT 46.265 -301.770 46.880 -301.765 ;
        RECT 46.260 -301.985 46.880 -301.770 ;
        RECT 46.260 -306.025 46.550 -301.985 ;
        RECT -28.315 -307.925 -27.620 -307.655 ;
        RECT -22.925 -307.895 -22.230 -307.625 ;
        RECT 46.265 -313.075 46.545 -306.025 ;
        RECT 139.375 -306.265 140.055 -301.130 ;
        RECT 141.100 -301.140 141.875 -301.130 ;
        RECT 141.200 -301.180 141.875 -301.140 ;
        RECT 157.370 -301.285 160.215 -301.105 ;
        RECT 157.370 -306.265 158.050 -301.285 ;
        RECT 159.440 -301.295 160.215 -301.285 ;
        RECT 159.540 -301.335 160.215 -301.295 ;
        RECT 139.375 -306.945 158.050 -306.265 ;
        RECT 139.375 -313.075 140.055 -306.945 ;
        RECT -165.310 -313.755 140.055 -313.075 ;
      LAYER met1 ;
        RECT -112.415 -313.130 -112.110 -270.495 ;
        RECT -28.695 -272.830 -28.015 -272.460 ;
        RECT -28.695 -274.740 -28.440 -272.830 ;
        RECT -28.695 -274.995 50.630 -274.740 ;
        RECT -64.870 -279.025 -63.885 -278.755 ;
        RECT -64.155 -284.180 -63.885 -279.025 ;
        RECT -72.210 -285.060 -63.885 -284.180 ;
        RECT -112.680 -313.745 -112.065 -313.130 ;
        RECT -72.210 -313.755 -71.330 -285.060 ;
        RECT -64.155 -286.045 -63.885 -285.060 ;
        RECT -64.405 -286.795 -63.755 -286.045 ;
        RECT 50.375 -301.745 50.630 -274.995 ;
        RECT -20.410 -302.000 50.630 -301.745 ;
        RECT -28.315 -307.740 -27.620 -307.655 ;
        RECT -22.925 -307.740 -22.230 -307.625 ;
        RECT -28.315 -307.750 -22.230 -307.740 ;
        RECT -20.410 -307.750 -20.270 -302.000 ;
        RECT -28.315 -307.880 -20.270 -307.750 ;
        RECT -28.315 -307.925 -27.620 -307.880 ;
        RECT -22.925 -307.890 -20.270 -307.880 ;
        RECT -22.925 -307.895 -22.230 -307.890 ;
    END
  END D16
  PIN D17
    ANTENNAGATEAREA 7.200000 ;
    PORT
      LAYER li1 ;
        RECT 36.685 -269.085 37.380 -268.815 ;
        RECT 42.075 -269.115 42.770 -268.845 ;
        RECT -111.460 -271.100 -111.155 -270.100 ;
        RECT -105.390 -271.100 -104.715 -271.055 ;
        RECT -111.460 -271.290 -104.715 -271.100 ;
        RECT -105.390 -271.325 -104.715 -271.290 ;
        RECT -111.460 -299.555 -111.160 -299.490 ;
        RECT -104.870 -299.555 -104.145 -299.500 ;
        RECT -111.460 -299.760 -104.145 -299.555 ;
        RECT -111.460 -300.675 -111.160 -299.760 ;
        RECT -104.870 -299.780 -104.145 -299.760 ;
        RECT 183.400 -300.995 184.075 -300.965 ;
        RECT 183.300 -301.005 184.075 -300.995 ;
        RECT 180.660 -301.185 184.075 -301.005 ;
        RECT 201.740 -301.150 202.415 -301.120 ;
        RECT 201.640 -301.160 202.415 -301.150 ;
        RECT 181.575 -306.320 182.255 -301.185 ;
        RECT 183.300 -301.195 184.075 -301.185 ;
        RECT 183.400 -301.235 184.075 -301.195 ;
        RECT 199.570 -301.340 202.415 -301.160 ;
        RECT 199.570 -306.320 200.250 -301.340 ;
        RECT 201.640 -301.350 202.415 -301.340 ;
        RECT 201.740 -301.390 202.415 -301.350 ;
        RECT 181.575 -307.000 200.250 -306.320 ;
        RECT 36.685 -307.925 37.380 -307.655 ;
        RECT 42.075 -307.895 42.770 -307.625 ;
        RECT 46.760 -307.915 47.085 -307.230 ;
        RECT 46.775 -311.715 47.045 -307.915 ;
        RECT 181.575 -314.070 182.255 -307.000 ;
        RECT -167.315 -314.750 182.255 -314.070 ;
      LAYER met1 ;
        RECT 36.685 -268.860 37.380 -268.815 ;
        RECT 42.075 -268.850 42.770 -268.845 ;
        RECT 41.565 -268.860 54.620 -268.850 ;
        RECT 36.685 -268.990 54.620 -268.860 ;
        RECT 36.685 -269.000 42.770 -268.990 ;
        RECT 36.685 -269.085 37.380 -269.000 ;
        RECT 42.075 -269.115 42.770 -269.000 ;
        RECT -111.460 -314.125 -111.155 -270.100 ;
        RECT 36.685 -307.740 37.380 -307.655 ;
        RECT 42.075 -307.740 42.770 -307.625 ;
        RECT 36.685 -307.750 42.770 -307.740 ;
        RECT 46.760 -307.750 47.085 -307.230 ;
        RECT 54.480 -307.750 54.620 -268.990 ;
        RECT 36.685 -307.880 54.620 -307.750 ;
        RECT 36.685 -307.925 37.380 -307.880 ;
        RECT 41.565 -307.890 54.620 -307.880 ;
        RECT 42.075 -307.895 42.770 -307.890 ;
        RECT 46.760 -307.915 47.085 -307.890 ;
        RECT 46.735 -314.100 47.040 -311.080 ;
        RECT -111.725 -314.740 -111.110 -314.125 ;
        RECT 46.470 -314.715 47.085 -314.100 ;
    END
  END D17
  PIN D18
    ANTENNAGATEAREA 7.200000 ;
    PORT
      LAYER li1 ;
        RECT 21.685 -269.085 22.380 -268.815 ;
        RECT 27.075 -269.115 27.770 -268.845 ;
        RECT -110.915 -270.685 -110.610 -269.670 ;
        RECT -107.070 -270.685 -106.395 -270.645 ;
        RECT -110.915 -270.860 -106.395 -270.685 ;
        RECT -107.165 -270.870 -106.395 -270.860 ;
        RECT -107.070 -270.915 -106.395 -270.870 ;
        RECT -110.910 -300.015 -110.610 -300.005 ;
        RECT -106.515 -300.015 -105.790 -299.975 ;
        RECT -110.910 -300.220 -105.790 -300.015 ;
        RECT -110.910 -301.190 -110.610 -300.220 ;
        RECT -106.515 -300.255 -105.790 -300.220 ;
        RECT 227.715 -301.190 228.390 -301.160 ;
        RECT 227.615 -301.200 228.390 -301.190 ;
        RECT 224.975 -301.380 228.390 -301.200 ;
        RECT 246.055 -301.345 246.730 -301.315 ;
        RECT 245.955 -301.355 246.730 -301.345 ;
        RECT 46.980 -304.775 47.595 -304.555 ;
        RECT 21.685 -307.925 22.380 -307.655 ;
        RECT 27.075 -307.895 27.770 -307.625 ;
        RECT 47.300 -311.715 47.570 -304.775 ;
        RECT 225.890 -306.445 226.570 -301.380 ;
        RECT 227.615 -301.390 228.390 -301.380 ;
        RECT 227.715 -301.430 228.390 -301.390 ;
        RECT 243.885 -301.535 246.730 -301.355 ;
        RECT 225.890 -306.515 226.805 -306.445 ;
        RECT 243.885 -306.515 244.565 -301.535 ;
        RECT 245.955 -301.545 246.730 -301.535 ;
        RECT 246.055 -301.585 246.730 -301.545 ;
        RECT 225.890 -307.195 244.565 -306.515 ;
        RECT 226.125 -315.235 226.805 -307.195 ;
        RECT -164.955 -315.915 226.805 -315.235 ;
      LAYER met1 ;
        RECT 21.685 -268.860 22.380 -268.815 ;
        RECT 27.075 -268.850 27.770 -268.845 ;
        RECT 27.075 -268.860 33.870 -268.850 ;
        RECT 21.685 -268.990 33.870 -268.860 ;
        RECT 21.685 -269.000 27.770 -268.990 ;
        RECT 21.685 -269.085 22.380 -269.000 ;
        RECT 27.075 -269.115 27.770 -269.000 ;
        RECT -110.915 -270.860 -110.610 -269.670 ;
        RECT -110.915 -300.005 -110.615 -270.860 ;
        RECT 33.730 -271.980 33.870 -268.990 ;
        RECT 33.730 -272.120 53.865 -271.980 ;
        RECT -110.915 -301.190 -110.610 -300.005 ;
        RECT -110.915 -315.290 -110.615 -301.190 ;
        RECT 46.935 -304.620 47.630 -304.545 ;
        RECT 53.725 -304.620 53.865 -272.120 ;
        RECT 33.730 -304.760 53.865 -304.620 ;
        RECT 21.685 -307.740 22.380 -307.655 ;
        RECT 27.075 -307.740 27.770 -307.625 ;
        RECT 21.685 -307.750 27.770 -307.740 ;
        RECT 33.730 -307.750 33.870 -304.760 ;
        RECT 46.935 -304.780 47.630 -304.760 ;
        RECT 21.685 -307.880 33.870 -307.750 ;
        RECT 21.685 -307.925 22.380 -307.880 ;
        RECT 27.075 -307.890 33.870 -307.880 ;
        RECT 27.075 -307.895 27.770 -307.890 ;
        RECT 47.325 -311.100 47.545 -311.085 ;
        RECT 47.280 -315.265 47.580 -311.100 ;
        RECT -111.195 -315.905 -110.580 -315.290 ;
        RECT 47.000 -315.880 47.615 -315.265 ;
    END
  END D18
  PIN D19
    ANTENNAGATEAREA 7.000000 ;
    PORT
      LAYER li1 ;
        RECT -97.790 -272.285 -97.105 -272.265 ;
        RECT -97.980 -272.295 -96.845 -272.285 ;
        RECT -94.790 -272.295 -94.420 -272.165 ;
        RECT -97.980 -272.485 -94.420 -272.295 ;
        RECT -97.790 -272.555 -97.105 -272.485 ;
        RECT -96.850 -272.490 -94.420 -272.485 ;
        RECT -96.850 -272.495 -96.495 -272.490 ;
        RECT -94.790 -272.520 -94.420 -272.490 ;
        RECT -110.420 -275.880 -110.120 -275.500 ;
        RECT -110.420 -276.080 -110.080 -275.880 ;
        RECT -110.420 -276.465 -110.120 -276.080 ;
        RECT -98.335 -276.465 -97.675 -276.420 ;
        RECT -110.420 -276.665 -97.675 -276.465 ;
        RECT -110.420 -276.685 -110.120 -276.665 ;
        RECT -98.335 -276.685 -97.675 -276.665 ;
        RECT 36.735 -280.340 37.430 -280.070 ;
        RECT 42.125 -280.370 42.820 -280.100 ;
        RECT 36.735 -296.670 37.430 -296.400 ;
        RECT 42.125 -296.640 42.820 -296.370 ;
        RECT 47.680 -296.695 48.405 -296.020 ;
        RECT -100.945 -297.800 -100.655 -297.325 ;
        RECT -98.910 -297.800 -98.195 -297.765 ;
        RECT -100.945 -297.980 -98.195 -297.800 ;
        RECT -100.945 -298.010 -100.655 -297.980 ;
        RECT -98.910 -298.065 -98.195 -297.980 ;
        RECT -110.420 -303.035 -110.130 -302.555 ;
        RECT -101.045 -303.035 -100.755 -302.555 ;
        RECT -110.420 -303.240 -100.755 -303.035 ;
        RECT 47.795 -312.800 48.075 -296.695 ;
        RECT 273.705 -301.020 274.380 -300.990 ;
        RECT 273.605 -301.030 274.380 -301.020 ;
        RECT 270.965 -301.210 274.380 -301.030 ;
        RECT 292.045 -301.175 292.720 -301.145 ;
        RECT 291.945 -301.185 292.720 -301.175 ;
        RECT 271.880 -306.345 272.560 -301.210 ;
        RECT 273.605 -301.220 274.380 -301.210 ;
        RECT 273.705 -301.260 274.380 -301.220 ;
        RECT 289.875 -301.365 292.720 -301.185 ;
        RECT 289.875 -306.345 290.555 -301.365 ;
        RECT 291.945 -301.375 292.720 -301.365 ;
        RECT 292.045 -301.415 292.720 -301.375 ;
        RECT 271.880 -307.025 290.555 -306.345 ;
        RECT 271.880 -316.510 272.560 -307.025 ;
        RECT -164.880 -317.190 272.560 -316.510 ;
      LAYER met1 ;
        RECT -97.790 -272.555 -97.105 -272.265 ;
        RECT -110.420 -316.575 -110.115 -275.495 ;
        RECT -97.755 -276.420 -97.555 -272.555 ;
        RECT -98.335 -276.465 -97.555 -276.420 ;
        RECT -98.570 -276.665 -97.555 -276.465 ;
        RECT -98.335 -276.685 -97.675 -276.665 ;
        RECT 36.735 -280.115 37.430 -280.070 ;
        RECT 42.125 -280.105 42.820 -280.100 ;
        RECT 48.775 -280.105 49.030 -280.065 ;
        RECT 42.125 -280.115 49.030 -280.105 ;
        RECT 36.735 -280.245 49.030 -280.115 ;
        RECT 36.735 -280.255 42.820 -280.245 ;
        RECT 36.735 -280.340 37.430 -280.255 ;
        RECT 42.125 -280.370 42.820 -280.255 ;
        RECT 48.775 -280.320 49.030 -280.245 ;
        RECT 36.735 -296.485 37.430 -296.400 ;
        RECT 42.125 -296.485 42.820 -296.370 ;
        RECT 36.735 -296.495 42.820 -296.485 ;
        RECT 47.680 -296.495 48.405 -296.020 ;
        RECT 48.840 -296.495 48.980 -280.320 ;
        RECT 36.735 -296.625 48.990 -296.495 ;
        RECT 36.735 -296.670 37.430 -296.625 ;
        RECT 42.125 -296.635 48.990 -296.625 ;
        RECT 42.125 -296.640 42.820 -296.635 ;
        RECT 47.680 -296.695 48.405 -296.635 ;
        RECT -100.945 -298.010 -100.655 -297.325 ;
        RECT -100.945 -302.555 -100.770 -298.010 ;
        RECT -101.045 -303.240 -100.755 -302.555 ;
        RECT 47.775 -316.550 48.080 -311.815 ;
        RECT -110.730 -317.190 -110.110 -316.575 ;
        RECT 47.465 -317.165 48.085 -316.550 ;
    END
  END D19
  PIN OUTB
    ANTENNAGATEAREA 34.399998 ;
    ANTENNADIFFAREA 14.500000 ;
    PORT
      LAYER li1 ;
        RECT 272.950 13.150 273.120 15.190 ;
        RECT 274.130 13.150 274.300 15.190 ;
        RECT 275.310 13.150 275.480 15.190 ;
        RECT 276.490 13.150 276.660 15.190 ;
        RECT 277.670 13.150 277.840 15.190 ;
        RECT 278.850 13.150 279.020 15.190 ;
        RECT 280.030 13.150 280.200 15.190 ;
        RECT 281.210 13.150 281.380 15.190 ;
        RECT 282.390 13.150 282.560 15.190 ;
        RECT 283.570 13.150 283.740 15.190 ;
        RECT 284.750 13.150 284.920 15.190 ;
        RECT 285.930 13.150 286.100 15.190 ;
        RECT 287.110 13.150 287.280 15.190 ;
        RECT 288.290 13.150 288.460 15.190 ;
        RECT 289.470 13.150 289.640 15.190 ;
        RECT 290.650 13.150 290.820 15.190 ;
        RECT 291.830 12.420 292.000 15.190 ;
        RECT 293.555 12.420 294.650 12.985 ;
        RECT 291.830 12.250 294.650 12.420 ;
        RECT 293.555 11.670 294.650 12.250 ;
        RECT 264.790 9.110 264.960 11.150 ;
        RECT 265.970 9.110 266.140 11.150 ;
        RECT 267.150 9.110 267.320 11.150 ;
        RECT 268.330 9.110 268.500 11.150 ;
        RECT 269.510 9.110 269.680 11.150 ;
        RECT 270.690 9.110 270.860 11.150 ;
        RECT 271.870 9.110 272.040 11.150 ;
        RECT 273.050 9.110 273.220 11.150 ;
        RECT -157.335 -45.300 -152.850 -43.985 ;
        RECT 294.565 -45.300 299.300 -44.155 ;
        RECT -171.415 -48.565 299.300 -45.300 ;
        RECT -157.335 -50.070 -152.850 -48.565 ;
        RECT 294.565 -49.545 299.300 -48.565 ;
        RECT 83.340 -274.080 84.515 -273.965 ;
        RECT -88.935 -274.385 -88.260 -274.345 ;
        RECT -89.035 -274.395 -88.260 -274.385 ;
        RECT -90.990 -274.575 -88.260 -274.395 ;
        RECT -113.155 -277.155 -112.650 -276.290 ;
        RECT -90.605 -277.155 -90.320 -274.575 ;
        RECT -89.035 -274.585 -88.260 -274.575 ;
        RECT -88.935 -274.615 -88.260 -274.585 ;
        RECT 56.300 -275.305 84.515 -274.080 ;
        RECT 92.195 -274.980 93.285 -273.750 ;
        RECT 133.400 -274.280 135.050 -273.865 ;
        RECT 56.300 -275.315 83.895 -275.305 ;
        RECT -113.155 -277.470 -90.320 -277.155 ;
        RECT 0.190 -276.280 0.875 -276.025 ;
        RECT -113.155 -277.505 -112.650 -277.470 ;
        RECT 0.190 -279.025 0.385 -276.280 ;
        RECT -4.765 -279.080 -3.925 -279.025 ;
        RECT -4.765 -279.370 -3.750 -279.080 ;
        RECT -4.765 -279.395 -3.925 -279.370 ;
        RECT -0.355 -279.395 0.485 -279.025 ;
        RECT 92.390 -279.265 93.100 -274.980 ;
        RECT 133.400 -275.175 139.295 -274.280 ;
        RECT 133.400 -275.335 135.050 -275.175 ;
        RECT 146.235 -276.945 146.910 -276.905 ;
        RECT 146.135 -276.955 146.910 -276.945 ;
        RECT 145.100 -277.135 146.910 -276.955 ;
        RECT 146.135 -277.145 146.910 -277.135 ;
        RECT 146.235 -277.175 146.910 -277.145 ;
        RECT -7.780 -280.320 -7.410 -279.525 ;
        RECT -26.235 -280.935 -25.575 -280.870 ;
        RECT -7.780 -280.935 -7.405 -280.320 ;
        RECT 0.190 -280.935 0.385 -279.395 ;
        RECT 92.205 -280.210 93.100 -279.265 ;
        RECT -28.265 -281.130 0.385 -280.935 ;
        RECT 100.045 -281.070 100.705 -280.395 ;
        RECT 111.785 -280.425 112.625 -280.370 ;
        RECT 111.785 -280.740 112.925 -280.425 ;
        RECT -26.235 -281.170 -25.575 -281.130 ;
        RECT 100.045 -282.745 100.575 -281.070 ;
        RECT 112.625 -281.535 112.925 -280.740 ;
        RECT 112.410 -282.745 113.070 -282.695 ;
        RECT 117.115 -282.745 117.800 -282.690 ;
        RECT -26.055 -283.565 -25.755 -282.845 ;
        RECT 100.045 -282.940 128.695 -282.745 ;
        RECT -26.055 -283.875 -24.855 -283.565 ;
        RECT -25.870 -283.880 -24.855 -283.875 ;
        RECT -25.695 -283.935 -24.855 -283.880 ;
        RECT 100.045 -284.910 100.240 -282.940 ;
        RECT 112.410 -282.995 113.070 -282.940 ;
        RECT 117.115 -282.990 117.800 -282.940 ;
        RECT 137.995 -283.130 139.290 -282.915 ;
        RECT 133.665 -283.685 139.290 -283.130 ;
        RECT 310.640 -283.435 315.270 -282.815 ;
        RECT 357.280 -283.350 360.600 -282.955 ;
        RECT 401.865 -283.160 407.905 -282.245 ;
        RECT 410.100 -283.150 410.775 -283.120 ;
        RECT 410.000 -283.160 410.775 -283.150 ;
        RECT 363.280 -283.340 363.955 -283.310 ;
        RECT 363.180 -283.350 363.955 -283.340 ;
        RECT 317.515 -283.425 318.190 -283.395 ;
        RECT 317.415 -283.435 318.190 -283.425 ;
        RECT 141.240 -283.675 141.915 -283.645 ;
        RECT 141.140 -283.685 141.915 -283.675 ;
        RECT 133.665 -283.865 141.915 -283.685 ;
        RECT 133.665 -284.155 139.290 -283.865 ;
        RECT 141.140 -283.875 141.915 -283.865 ;
        RECT 141.240 -283.915 141.915 -283.875 ;
        RECT 178.000 -283.740 181.240 -283.470 ;
        RECT 183.440 -283.730 184.115 -283.700 ;
        RECT 183.340 -283.740 184.115 -283.730 ;
        RECT 137.995 -284.230 139.290 -284.155 ;
        RECT 178.000 -283.920 184.115 -283.740 ;
        RECT 268.005 -283.765 271.650 -283.440 ;
        RECT 310.640 -283.615 318.190 -283.435 ;
        RECT 273.745 -283.755 274.420 -283.725 ;
        RECT 273.645 -283.765 274.420 -283.755 ;
        RECT 178.000 -284.200 181.240 -283.920 ;
        RECT 183.340 -283.930 184.115 -283.920 ;
        RECT 183.440 -283.970 184.115 -283.930 ;
        RECT 221.410 -283.935 225.245 -283.900 ;
        RECT 227.755 -283.925 228.430 -283.895 ;
        RECT 227.655 -283.935 228.430 -283.925 ;
        RECT 221.410 -284.115 228.430 -283.935 ;
        RECT 99.945 -285.280 100.785 -284.910 ;
        RECT 117.255 -284.935 117.555 -284.570 ;
        RECT 117.855 -284.935 118.695 -284.910 ;
        RECT 117.255 -285.225 118.695 -284.935 ;
        RECT 117.255 -285.230 117.555 -285.225 ;
        RECT 117.855 -285.280 118.695 -285.225 ;
        RECT -12.195 -292.860 -11.355 -292.805 ;
        RECT -12.495 -293.175 -11.355 -292.860 ;
        RECT -12.495 -293.970 -12.195 -293.175 ;
        RECT -17.370 -295.180 -16.685 -295.125 ;
        RECT -12.640 -295.180 -11.980 -295.130 ;
        RECT -28.265 -295.375 0.385 -295.180 ;
        RECT -17.370 -295.425 -16.685 -295.375 ;
        RECT -12.640 -295.430 -11.980 -295.375 ;
        RECT -18.265 -297.370 -17.425 -297.345 ;
        RECT -17.125 -297.370 -16.825 -297.005 ;
        RECT 0.190 -297.345 0.385 -295.375 ;
        RECT -18.265 -297.660 -16.825 -297.370 ;
        RECT -18.265 -297.715 -17.425 -297.660 ;
        RECT -17.125 -297.665 -16.825 -297.660 ;
        RECT -0.355 -297.715 0.485 -297.345 ;
        RECT 0.190 -300.460 0.385 -297.715 ;
        RECT 0.190 -300.715 0.875 -300.460 ;
        RECT 49.150 -301.100 50.105 -301.070 ;
        RECT 49.150 -301.515 51.965 -301.100 ;
        RECT 49.150 -301.605 50.105 -301.515 ;
        RECT 51.550 -310.840 51.965 -301.515 ;
        RECT 59.305 -303.520 60.145 -303.150 ;
        RECT 76.615 -303.205 76.915 -303.200 ;
        RECT 77.215 -303.205 78.055 -303.150 ;
        RECT 76.615 -303.495 78.055 -303.205 ;
        RECT 56.300 -305.490 57.775 -305.000 ;
        RECT 59.405 -305.490 59.600 -303.520 ;
        RECT 76.615 -303.860 76.915 -303.495 ;
        RECT 77.215 -303.520 78.055 -303.495 ;
        RECT 71.770 -305.490 72.430 -305.435 ;
        RECT 76.475 -305.490 77.160 -305.440 ;
        RECT 56.300 -305.685 88.055 -305.490 ;
        RECT 56.300 -306.015 57.775 -305.685 ;
        RECT 71.770 -305.735 72.430 -305.685 ;
        RECT 76.475 -305.740 77.160 -305.685 ;
        RECT 71.985 -307.690 72.285 -306.895 ;
        RECT 71.145 -308.005 72.285 -307.690 ;
        RECT 71.145 -308.060 71.985 -308.005 ;
        RECT 51.430 -311.735 52.070 -310.840 ;
        RECT 136.525 -312.015 137.630 -311.040 ;
        RECT 178.000 -311.115 178.730 -284.200 ;
        RECT 221.410 -284.630 225.245 -284.115 ;
        RECT 227.655 -284.125 228.430 -284.115 ;
        RECT 227.755 -284.165 228.430 -284.125 ;
        RECT 268.005 -283.945 274.420 -283.765 ;
        RECT 268.005 -284.170 271.650 -283.945 ;
        RECT 273.645 -283.955 274.420 -283.945 ;
        RECT 273.745 -283.995 274.420 -283.955 ;
        RECT 310.640 -284.010 315.270 -283.615 ;
        RECT 317.415 -283.625 318.190 -283.615 ;
        RECT 317.515 -283.665 318.190 -283.625 ;
        RECT 357.280 -283.530 363.955 -283.350 ;
        RECT 357.280 -283.880 360.600 -283.530 ;
        RECT 363.180 -283.540 363.955 -283.530 ;
        RECT 363.280 -283.580 363.955 -283.540 ;
        RECT 401.865 -283.340 410.775 -283.160 ;
        RECT 401.865 -283.715 407.905 -283.340 ;
        RECT 410.000 -283.350 410.775 -283.340 ;
        RECT 410.100 -283.390 410.775 -283.350 ;
        RECT 177.655 -312.130 179.025 -311.115 ;
        RECT 221.410 -311.205 222.140 -284.630 ;
        RECT 268.005 -311.010 268.735 -284.170 ;
        RECT 310.640 -310.935 311.835 -284.010 ;
        RECT 357.280 -310.920 358.205 -283.880 ;
        RECT 221.140 -311.900 222.400 -311.205 ;
        RECT 267.835 -312.035 268.995 -311.010 ;
        RECT 310.330 -312.095 312.070 -310.935 ;
        RECT 356.855 -312.145 358.765 -310.920 ;
        RECT 401.865 -310.935 403.335 -283.715 ;
        RECT 401.620 -312.125 403.620 -310.935 ;
        RECT -158.395 -319.180 -152.600 -318.125 ;
        RECT -158.395 -322.505 -152.610 -319.180 ;
        RECT -114.000 -322.505 -112.935 -322.345 ;
        RECT -158.395 -323.185 57.775 -322.505 ;
        RECT -158.395 -324.325 -152.610 -323.185 ;
        RECT -114.000 -323.235 -112.935 -323.185 ;
      LAYER met1 ;
        RECT 272.920 12.815 273.150 15.170 ;
        RECT 274.100 12.815 274.330 15.170 ;
        RECT 275.280 12.815 275.510 15.170 ;
        RECT 276.460 12.815 276.690 15.170 ;
        RECT 277.640 12.815 277.870 15.170 ;
        RECT 278.820 12.815 279.050 15.170 ;
        RECT 280.000 12.815 280.230 15.170 ;
        RECT 281.180 12.815 281.410 15.170 ;
        RECT 282.360 12.815 282.590 15.170 ;
        RECT 283.540 12.815 283.770 15.170 ;
        RECT 284.720 12.815 284.950 15.170 ;
        RECT 285.900 12.815 286.130 15.170 ;
        RECT 287.080 12.815 287.310 15.170 ;
        RECT 288.260 12.815 288.490 15.170 ;
        RECT 289.440 12.815 289.670 15.170 ;
        RECT 290.620 12.815 290.850 15.170 ;
        RECT 291.800 12.815 292.030 15.170 ;
        RECT 272.790 12.445 292.175 12.815 ;
        RECT 273.020 11.865 273.250 12.445 ;
        RECT 264.760 11.635 273.250 11.865 ;
        RECT 264.760 9.130 264.990 11.635 ;
        RECT 265.940 9.130 266.170 11.635 ;
        RECT 267.120 9.130 267.350 11.635 ;
        RECT 268.300 9.130 268.530 11.635 ;
        RECT 269.480 9.130 269.710 11.635 ;
        RECT 270.660 9.130 270.890 11.635 ;
        RECT 271.840 9.130 272.070 11.635 ;
        RECT 273.020 9.130 273.250 11.635 ;
        RECT 293.530 11.300 298.080 13.520 ;
        RECT -158.395 -312.985 -152.610 -43.395 ;
        RECT 295.860 -44.155 298.080 11.300 ;
        RECT 294.565 -49.545 299.300 -44.155 ;
        RECT 82.985 -273.865 134.150 -273.665 ;
        RECT 0.190 -276.280 50.005 -276.025 ;
        RECT -113.155 -276.565 -112.650 -276.290 ;
        RECT -113.915 -277.505 -112.650 -276.565 ;
        RECT -113.915 -277.720 -112.715 -277.505 ;
        RECT -158.395 -319.180 -152.600 -312.985 ;
        RECT -158.395 -324.325 -152.610 -319.180 ;
        RECT -113.915 -322.345 -113.235 -277.720 ;
        RECT -26.235 -281.170 -25.575 -280.870 ;
        RECT -26.055 -283.505 -25.755 -281.170 ;
        RECT -17.370 -295.425 -16.685 -295.125 ;
        RECT -12.495 -295.130 -12.195 -293.310 ;
        RECT -17.125 -297.665 -16.825 -295.425 ;
        RECT -12.640 -295.430 -11.980 -295.130 ;
        RECT 49.750 -300.460 50.005 -276.280 ;
        RECT 0.190 -300.715 50.005 -300.460 ;
        RECT 49.750 -301.070 50.005 -300.715 ;
        RECT 49.150 -301.605 50.105 -301.070 ;
        RECT 56.300 -310.530 57.775 -274.080 ;
        RECT 82.985 -275.335 135.050 -273.865 ;
        RECT 137.990 -274.625 139.055 -274.430 ;
        RECT 137.990 -274.895 145.180 -274.625 ;
        RECT 137.990 -275.095 139.055 -274.895 ;
        RECT 82.985 -275.425 134.875 -275.335 ;
        RECT 92.205 -279.645 93.100 -279.265 ;
        RECT 92.205 -280.020 100.555 -279.645 ;
        RECT 92.205 -280.210 93.100 -280.020 ;
        RECT 100.180 -280.395 100.555 -280.020 ;
        RECT 100.045 -281.070 100.705 -280.395 ;
        RECT 112.625 -282.695 112.925 -280.875 ;
        RECT 112.410 -282.995 113.070 -282.695 ;
        RECT 117.115 -282.990 117.800 -282.690 ;
        RECT 117.255 -285.230 117.555 -282.990 ;
        RECT 71.770 -305.735 72.430 -305.435 ;
        RECT 76.615 -305.440 76.915 -303.200 ;
        RECT 71.985 -307.555 72.285 -305.735 ;
        RECT 76.475 -305.740 77.160 -305.440 ;
        RECT 51.040 -311.875 57.775 -310.530 ;
        RECT -114.000 -323.235 -112.935 -322.345 ;
        RECT 56.300 -323.185 57.775 -311.875 ;
        RECT 133.650 -310.920 134.875 -275.425 ;
        RECT 144.910 -276.345 145.180 -274.895 ;
        RECT 144.910 -276.615 146.550 -276.345 ;
        RECT 146.280 -276.890 146.550 -276.615 ;
        RECT 146.150 -277.180 146.945 -276.890 ;
        RECT 137.995 -284.230 139.290 -282.915 ;
        RECT 133.650 -312.145 413.640 -310.920 ;
    END
  END OUTB
  PIN OUT
    ANTENNAGATEAREA 34.399998 ;
    ANTENNADIFFAREA 14.500000 ;
    PORT
      LAYER li1 ;
        RECT 271.935 -1.405 272.105 0.635 ;
        RECT 273.115 -1.405 273.285 0.635 ;
        RECT 274.295 -1.405 274.465 0.635 ;
        RECT 275.475 -1.405 275.645 0.635 ;
        RECT 276.655 -1.405 276.825 0.635 ;
        RECT 277.835 -1.405 278.005 0.635 ;
        RECT 279.015 -1.405 279.185 0.635 ;
        RECT 280.195 -1.405 280.365 0.635 ;
        RECT 281.375 -1.405 281.545 0.635 ;
        RECT 282.555 -1.405 282.725 0.635 ;
        RECT 283.735 -1.405 283.905 0.635 ;
        RECT 284.915 -1.405 285.085 0.635 ;
        RECT 286.095 -1.405 286.265 0.635 ;
        RECT 287.275 -1.405 287.445 0.635 ;
        RECT 288.455 -1.405 288.625 0.635 ;
        RECT 289.635 -1.405 289.805 0.635 ;
        RECT 290.815 -2.135 290.985 0.635 ;
        RECT 303.065 -2.135 305.390 -1.690 ;
        RECT 290.815 -2.305 305.390 -2.135 ;
        RECT 291.620 -3.090 305.390 -2.305 ;
        RECT 303.065 -3.345 305.390 -3.090 ;
        RECT 263.775 -5.445 263.945 -3.405 ;
        RECT 264.955 -5.445 265.125 -3.405 ;
        RECT 266.135 -5.445 266.305 -3.405 ;
        RECT 267.315 -5.445 267.485 -3.405 ;
        RECT 268.495 -5.445 268.665 -3.405 ;
        RECT 269.675 -5.445 269.845 -3.405 ;
        RECT 270.855 -5.445 271.025 -3.405 ;
        RECT 272.035 -5.445 272.205 -3.405 ;
        RECT -145.865 -49.915 -142.360 -49.910 ;
        RECT 302.115 -49.915 307.270 -48.085 ;
        RECT -146.735 -52.610 307.270 -49.915 ;
        RECT -147.820 -53.405 307.270 -52.610 ;
        RECT -147.820 -58.755 -141.430 -53.405 ;
        RECT 302.115 -53.655 307.270 -53.405 ;
        RECT -145.865 -62.975 -142.360 -58.755 ;
        RECT -171.845 -66.480 -142.360 -62.975 ;
        RECT 79.825 -183.525 81.000 -183.410 ;
        RECT -92.450 -183.830 -91.775 -183.790 ;
        RECT -92.550 -183.840 -91.775 -183.830 ;
        RECT -94.505 -184.020 -91.775 -183.840 ;
        RECT -116.670 -186.600 -116.165 -185.735 ;
        RECT -94.120 -186.600 -93.835 -184.020 ;
        RECT -92.550 -184.030 -91.775 -184.020 ;
        RECT -92.450 -184.060 -91.775 -184.030 ;
        RECT 52.785 -184.750 81.000 -183.525 ;
        RECT 88.680 -184.425 89.770 -183.195 ;
        RECT 129.885 -183.725 131.535 -183.310 ;
        RECT 52.785 -184.760 80.380 -184.750 ;
        RECT -116.670 -186.915 -93.835 -186.600 ;
        RECT -3.325 -185.725 -2.640 -185.470 ;
        RECT -116.670 -186.950 -116.165 -186.915 ;
        RECT -3.325 -188.470 -3.130 -185.725 ;
        RECT -8.280 -188.525 -7.440 -188.470 ;
        RECT -8.280 -188.815 -7.265 -188.525 ;
        RECT -8.280 -188.840 -7.440 -188.815 ;
        RECT -3.870 -188.840 -3.030 -188.470 ;
        RECT 88.875 -188.710 89.585 -184.425 ;
        RECT 129.885 -184.620 135.780 -183.725 ;
        RECT 129.885 -184.780 131.535 -184.620 ;
        RECT 142.720 -186.390 143.395 -186.350 ;
        RECT 142.620 -186.400 143.395 -186.390 ;
        RECT 141.585 -186.580 143.395 -186.400 ;
        RECT 142.620 -186.590 143.395 -186.580 ;
        RECT 142.720 -186.620 143.395 -186.590 ;
        RECT -11.295 -189.765 -10.925 -188.970 ;
        RECT -29.750 -190.380 -29.090 -190.315 ;
        RECT -11.295 -190.380 -10.920 -189.765 ;
        RECT -3.325 -190.380 -3.130 -188.840 ;
        RECT 88.690 -189.655 89.585 -188.710 ;
        RECT -31.780 -190.575 -3.130 -190.380 ;
        RECT 96.530 -190.515 97.190 -189.840 ;
        RECT 108.270 -189.870 109.110 -189.815 ;
        RECT 108.270 -190.185 109.410 -189.870 ;
        RECT -29.750 -190.615 -29.090 -190.575 ;
        RECT 96.530 -192.190 97.060 -190.515 ;
        RECT 109.110 -190.980 109.410 -190.185 ;
        RECT 108.895 -192.190 109.555 -192.140 ;
        RECT 113.600 -192.190 114.285 -192.135 ;
        RECT -29.570 -193.010 -29.270 -192.290 ;
        RECT 96.530 -192.385 125.180 -192.190 ;
        RECT -29.570 -193.320 -28.370 -193.010 ;
        RECT -29.385 -193.325 -28.370 -193.320 ;
        RECT -29.210 -193.380 -28.370 -193.325 ;
        RECT 96.530 -194.355 96.725 -192.385 ;
        RECT 108.895 -192.440 109.555 -192.385 ;
        RECT 113.600 -192.435 114.285 -192.385 ;
        RECT 134.480 -192.575 135.775 -192.360 ;
        RECT 130.150 -193.130 135.775 -192.575 ;
        RECT 307.125 -192.880 311.755 -192.260 ;
        RECT 353.765 -192.795 357.085 -192.400 ;
        RECT 398.350 -192.605 404.390 -191.690 ;
        RECT 406.585 -192.595 407.260 -192.565 ;
        RECT 406.485 -192.605 407.260 -192.595 ;
        RECT 359.765 -192.785 360.440 -192.755 ;
        RECT 359.665 -192.795 360.440 -192.785 ;
        RECT 314.000 -192.870 314.675 -192.840 ;
        RECT 313.900 -192.880 314.675 -192.870 ;
        RECT 137.725 -193.120 138.400 -193.090 ;
        RECT 137.625 -193.130 138.400 -193.120 ;
        RECT 130.150 -193.310 138.400 -193.130 ;
        RECT 130.150 -193.600 135.775 -193.310 ;
        RECT 137.625 -193.320 138.400 -193.310 ;
        RECT 137.725 -193.360 138.400 -193.320 ;
        RECT 174.485 -193.185 177.725 -192.915 ;
        RECT 179.925 -193.175 180.600 -193.145 ;
        RECT 179.825 -193.185 180.600 -193.175 ;
        RECT 134.480 -193.675 135.775 -193.600 ;
        RECT 174.485 -193.365 180.600 -193.185 ;
        RECT 264.490 -193.210 268.135 -192.885 ;
        RECT 307.125 -193.060 314.675 -192.880 ;
        RECT 270.230 -193.200 270.905 -193.170 ;
        RECT 270.130 -193.210 270.905 -193.200 ;
        RECT 174.485 -193.645 177.725 -193.365 ;
        RECT 179.825 -193.375 180.600 -193.365 ;
        RECT 179.925 -193.415 180.600 -193.375 ;
        RECT 217.895 -193.380 221.730 -193.345 ;
        RECT 224.240 -193.370 224.915 -193.340 ;
        RECT 224.140 -193.380 224.915 -193.370 ;
        RECT 217.895 -193.560 224.915 -193.380 ;
        RECT 96.430 -194.725 97.270 -194.355 ;
        RECT 113.740 -194.380 114.040 -194.015 ;
        RECT 114.340 -194.380 115.180 -194.355 ;
        RECT 113.740 -194.670 115.180 -194.380 ;
        RECT 113.740 -194.675 114.040 -194.670 ;
        RECT 114.340 -194.725 115.180 -194.670 ;
        RECT -15.710 -202.305 -14.870 -202.250 ;
        RECT -16.010 -202.620 -14.870 -202.305 ;
        RECT -16.010 -203.415 -15.710 -202.620 ;
        RECT -20.885 -204.625 -20.200 -204.570 ;
        RECT -16.155 -204.625 -15.495 -204.575 ;
        RECT -31.780 -204.820 -3.130 -204.625 ;
        RECT -20.885 -204.870 -20.200 -204.820 ;
        RECT -16.155 -204.875 -15.495 -204.820 ;
        RECT -21.780 -206.815 -20.940 -206.790 ;
        RECT -20.640 -206.815 -20.340 -206.450 ;
        RECT -3.325 -206.790 -3.130 -204.820 ;
        RECT -21.780 -207.105 -20.340 -206.815 ;
        RECT -21.780 -207.160 -20.940 -207.105 ;
        RECT -20.640 -207.110 -20.340 -207.105 ;
        RECT -3.870 -207.160 -3.030 -206.790 ;
        RECT -3.325 -209.905 -3.130 -207.160 ;
        RECT -3.325 -210.160 -2.640 -209.905 ;
        RECT 45.635 -210.545 46.590 -210.515 ;
        RECT 45.635 -210.960 48.450 -210.545 ;
        RECT 45.635 -211.050 46.590 -210.960 ;
        RECT 48.035 -220.285 48.450 -210.960 ;
        RECT 55.790 -212.965 56.630 -212.595 ;
        RECT 73.100 -212.650 73.400 -212.645 ;
        RECT 73.700 -212.650 74.540 -212.595 ;
        RECT 73.100 -212.940 74.540 -212.650 ;
        RECT 52.785 -214.935 54.260 -214.445 ;
        RECT 55.890 -214.935 56.085 -212.965 ;
        RECT 73.100 -213.305 73.400 -212.940 ;
        RECT 73.700 -212.965 74.540 -212.940 ;
        RECT 68.255 -214.935 68.915 -214.880 ;
        RECT 72.960 -214.935 73.645 -214.885 ;
        RECT 52.785 -215.130 84.540 -214.935 ;
        RECT 52.785 -215.460 54.260 -215.130 ;
        RECT 68.255 -215.180 68.915 -215.130 ;
        RECT 72.960 -215.185 73.645 -215.130 ;
        RECT 68.470 -217.135 68.770 -216.340 ;
        RECT 67.630 -217.450 68.770 -217.135 ;
        RECT 67.630 -217.505 68.470 -217.450 ;
        RECT 47.915 -221.180 48.555 -220.285 ;
        RECT 133.010 -221.460 134.115 -220.485 ;
        RECT 174.485 -220.560 175.215 -193.645 ;
        RECT 217.895 -194.075 221.730 -193.560 ;
        RECT 224.140 -193.570 224.915 -193.560 ;
        RECT 224.240 -193.610 224.915 -193.570 ;
        RECT 264.490 -193.390 270.905 -193.210 ;
        RECT 264.490 -193.615 268.135 -193.390 ;
        RECT 270.130 -193.400 270.905 -193.390 ;
        RECT 270.230 -193.440 270.905 -193.400 ;
        RECT 307.125 -193.455 311.755 -193.060 ;
        RECT 313.900 -193.070 314.675 -193.060 ;
        RECT 314.000 -193.110 314.675 -193.070 ;
        RECT 353.765 -192.975 360.440 -192.795 ;
        RECT 353.765 -193.325 357.085 -192.975 ;
        RECT 359.665 -192.985 360.440 -192.975 ;
        RECT 359.765 -193.025 360.440 -192.985 ;
        RECT 398.350 -192.785 407.260 -192.605 ;
        RECT 398.350 -193.160 404.390 -192.785 ;
        RECT 406.485 -192.795 407.260 -192.785 ;
        RECT 406.585 -192.835 407.260 -192.795 ;
        RECT 174.140 -221.575 175.510 -220.560 ;
        RECT 217.895 -220.650 218.625 -194.075 ;
        RECT 264.490 -220.455 265.220 -193.615 ;
        RECT 307.125 -220.380 308.320 -193.455 ;
        RECT 353.765 -220.365 354.690 -193.325 ;
        RECT 217.625 -221.345 218.885 -220.650 ;
        RECT 264.320 -221.480 265.480 -220.455 ;
        RECT 306.815 -221.540 308.555 -220.380 ;
        RECT 353.340 -221.590 355.250 -220.365 ;
        RECT 398.350 -220.380 399.820 -193.160 ;
        RECT 398.105 -221.570 400.105 -220.380 ;
        RECT -147.900 -231.950 -140.785 -227.055 ;
        RECT -117.515 -231.950 -116.450 -231.790 ;
        RECT -147.900 -232.630 54.260 -231.950 ;
        RECT -117.515 -232.680 -116.450 -232.630 ;
      LAYER met1 ;
        RECT 271.905 -1.740 272.135 0.615 ;
        RECT 273.085 -1.740 273.315 0.615 ;
        RECT 274.265 -1.740 274.495 0.615 ;
        RECT 275.445 -1.740 275.675 0.615 ;
        RECT 276.625 -1.740 276.855 0.615 ;
        RECT 277.805 -1.740 278.035 0.615 ;
        RECT 278.985 -1.740 279.215 0.615 ;
        RECT 280.165 -1.740 280.395 0.615 ;
        RECT 281.345 -1.740 281.575 0.615 ;
        RECT 282.525 -1.740 282.755 0.615 ;
        RECT 283.705 -1.740 283.935 0.615 ;
        RECT 284.885 -1.740 285.115 0.615 ;
        RECT 286.065 -1.740 286.295 0.615 ;
        RECT 287.245 -1.740 287.475 0.615 ;
        RECT 288.425 -1.740 288.655 0.615 ;
        RECT 289.605 -1.740 289.835 0.615 ;
        RECT 290.785 -1.740 291.015 0.615 ;
        RECT 271.775 -2.110 291.160 -1.740 ;
        RECT 272.005 -2.690 272.235 -2.110 ;
        RECT 263.745 -2.920 272.235 -2.690 ;
        RECT 263.745 -5.425 263.975 -2.920 ;
        RECT 264.925 -5.425 265.155 -2.920 ;
        RECT 266.105 -5.425 266.335 -2.920 ;
        RECT 267.285 -5.425 267.515 -2.920 ;
        RECT 268.465 -5.425 268.695 -2.920 ;
        RECT 269.645 -5.425 269.875 -2.920 ;
        RECT 270.825 -5.425 271.055 -2.920 ;
        RECT 272.005 -5.425 272.235 -2.920 ;
        RECT 302.745 -48.085 305.795 -1.140 ;
        RECT -147.900 -232.360 -140.785 -52.530 ;
        RECT 302.115 -53.655 307.270 -48.085 ;
        RECT 79.470 -183.310 130.635 -183.110 ;
        RECT -3.325 -185.725 46.490 -185.470 ;
        RECT -116.670 -186.010 -116.165 -185.735 ;
        RECT -117.430 -186.950 -116.165 -186.010 ;
        RECT -117.430 -187.165 -116.230 -186.950 ;
        RECT -117.430 -231.790 -116.750 -187.165 ;
        RECT -29.750 -190.615 -29.090 -190.315 ;
        RECT -29.570 -192.950 -29.270 -190.615 ;
        RECT -20.885 -204.870 -20.200 -204.570 ;
        RECT -16.010 -204.575 -15.710 -202.755 ;
        RECT -20.640 -207.110 -20.340 -204.870 ;
        RECT -16.155 -204.875 -15.495 -204.575 ;
        RECT 46.235 -209.905 46.490 -185.725 ;
        RECT -3.325 -210.160 46.490 -209.905 ;
        RECT 46.235 -210.515 46.490 -210.160 ;
        RECT 45.635 -211.050 46.590 -210.515 ;
        RECT 52.785 -219.975 54.260 -183.525 ;
        RECT 79.470 -184.780 131.535 -183.310 ;
        RECT 134.475 -184.070 135.540 -183.875 ;
        RECT 134.475 -184.340 141.665 -184.070 ;
        RECT 134.475 -184.540 135.540 -184.340 ;
        RECT 79.470 -184.870 131.360 -184.780 ;
        RECT 88.690 -189.090 89.585 -188.710 ;
        RECT 88.690 -189.465 97.040 -189.090 ;
        RECT 88.690 -189.655 89.585 -189.465 ;
        RECT 96.665 -189.840 97.040 -189.465 ;
        RECT 96.530 -190.515 97.190 -189.840 ;
        RECT 109.110 -192.140 109.410 -190.320 ;
        RECT 108.895 -192.440 109.555 -192.140 ;
        RECT 113.600 -192.435 114.285 -192.135 ;
        RECT 113.740 -194.675 114.040 -192.435 ;
        RECT 68.255 -215.180 68.915 -214.880 ;
        RECT 73.100 -214.885 73.400 -212.645 ;
        RECT 68.470 -217.000 68.770 -215.180 ;
        RECT 72.960 -215.185 73.645 -214.885 ;
        RECT 47.525 -221.320 54.260 -219.975 ;
        RECT -117.515 -232.680 -116.450 -231.790 ;
        RECT 52.785 -232.630 54.260 -221.320 ;
        RECT 130.135 -220.365 131.360 -184.870 ;
        RECT 141.395 -185.790 141.665 -184.340 ;
        RECT 141.395 -186.060 143.035 -185.790 ;
        RECT 142.765 -186.335 143.035 -186.060 ;
        RECT 142.635 -186.625 143.430 -186.335 ;
        RECT 134.480 -193.675 135.775 -192.360 ;
        RECT 130.135 -221.590 410.125 -220.365 ;
    END
  END OUT
  PIN PRE_SCALAR
    ANTENNADIFFAREA 14.500000 ;
    PORT
      LAYER li1 ;
        RECT -67.045 7.125 -66.875 9.895 ;
        RECT -65.865 7.855 -65.695 9.895 ;
        RECT -64.685 7.855 -64.515 9.895 ;
        RECT -63.505 7.855 -63.335 9.895 ;
        RECT -62.325 7.855 -62.155 9.895 ;
        RECT -61.145 7.855 -60.975 9.895 ;
        RECT -59.965 7.855 -59.795 9.895 ;
        RECT -58.785 7.855 -58.615 9.895 ;
        RECT -57.605 7.855 -57.435 9.895 ;
        RECT -56.425 7.855 -56.255 9.895 ;
        RECT -55.245 7.855 -55.075 9.895 ;
        RECT -54.065 7.855 -53.895 9.895 ;
        RECT -52.885 7.855 -52.715 9.895 ;
        RECT -51.705 7.855 -51.535 9.895 ;
        RECT -50.525 7.855 -50.355 9.895 ;
        RECT -49.345 7.855 -49.175 9.895 ;
        RECT -48.165 7.855 -47.995 9.895 ;
        RECT -113.320 6.955 -66.875 7.125 ;
        RECT -48.265 3.815 -48.095 5.855 ;
        RECT -47.085 3.815 -46.915 5.855 ;
        RECT -45.905 3.815 -45.735 5.855 ;
        RECT -44.725 3.815 -44.555 5.855 ;
        RECT -43.545 3.815 -43.375 5.855 ;
        RECT -42.365 3.815 -42.195 5.855 ;
        RECT -41.185 3.815 -41.015 5.855 ;
        RECT -40.005 3.815 -39.835 5.855 ;
      LAYER met1 ;
        RECT -67.075 7.520 -66.845 9.875 ;
        RECT -65.895 7.520 -65.665 9.875 ;
        RECT -64.715 7.520 -64.485 9.875 ;
        RECT -63.535 7.520 -63.305 9.875 ;
        RECT -62.355 7.520 -62.125 9.875 ;
        RECT -61.175 7.520 -60.945 9.875 ;
        RECT -59.995 7.520 -59.765 9.875 ;
        RECT -58.815 7.520 -58.585 9.875 ;
        RECT -57.635 7.520 -57.405 9.875 ;
        RECT -56.455 7.520 -56.225 9.875 ;
        RECT -55.275 7.520 -55.045 9.875 ;
        RECT -54.095 7.520 -53.865 9.875 ;
        RECT -52.915 7.520 -52.685 9.875 ;
        RECT -51.735 7.520 -51.505 9.875 ;
        RECT -50.555 7.520 -50.325 9.875 ;
        RECT -49.375 7.520 -49.145 9.875 ;
        RECT -48.195 7.520 -47.965 9.875 ;
        RECT -67.220 7.150 -47.835 7.520 ;
        RECT -48.295 6.570 -48.065 7.150 ;
        RECT -48.295 6.340 -39.805 6.570 ;
        RECT -48.295 3.835 -48.065 6.340 ;
        RECT -47.115 3.835 -46.885 6.340 ;
        RECT -45.935 3.835 -45.705 6.340 ;
        RECT -44.755 3.835 -44.525 6.340 ;
        RECT -43.575 3.835 -43.345 6.340 ;
        RECT -42.395 3.835 -42.165 6.340 ;
        RECT -41.215 3.835 -40.985 6.340 ;
        RECT -40.035 3.835 -39.805 6.340 ;
    END
  END PRE_SCALAR
  PIN S1
    ANTENNAGATEAREA 4.600000 ;
    PORT
      LAYER li1 ;
        RECT -19.135 8.475 -17.640 8.845 ;
        RECT -18.495 5.450 -18.235 8.475 ;
        RECT -14.230 5.450 -13.390 5.520 ;
        RECT -18.495 5.190 -13.390 5.450 ;
        RECT -18.475 1.060 -18.215 5.190 ;
        RECT -14.230 5.150 -13.390 5.190 ;
        RECT -114.810 0.800 -18.215 1.060 ;
    END
  END S1
  PIN S7
    ANTENNAGATEAREA 4.600000 ;
    PORT
      LAYER li1 ;
        RECT 310.750 -15.900 312.245 -15.530 ;
        RECT 311.390 -18.925 311.650 -15.900 ;
        RECT 315.655 -18.925 316.495 -18.855 ;
        RECT 311.390 -19.185 316.495 -18.925 ;
        RECT 312.160 -20.695 313.895 -19.185 ;
        RECT 315.655 -19.225 316.495 -19.185 ;
        RECT 311.230 -62.730 315.360 -62.205 ;
        RECT -134.980 -65.605 315.360 -62.730 ;
        RECT -134.980 -69.955 -132.105 -65.605 ;
        RECT 311.230 -65.900 315.360 -65.605 ;
        RECT -172.525 -72.830 -132.105 -69.955 ;
      LAYER met1 ;
        RECT 312.160 -20.695 313.895 -18.930 ;
        RECT 312.325 -62.205 313.660 -20.695 ;
        RECT 311.230 -65.900 315.360 -62.205 ;
    END
  END S7
  PIN DIV_OUT
    ANTENNADIFFAREA 14.500000 ;
    PORT
      LAYER li1 ;
        RECT -56.465 -78.660 -56.295 -76.620 ;
        RECT -55.285 -78.660 -55.115 -76.620 ;
        RECT -54.105 -78.660 -53.935 -76.620 ;
        RECT -52.925 -78.660 -52.755 -76.620 ;
        RECT -51.745 -78.660 -51.575 -76.620 ;
        RECT -50.565 -78.660 -50.395 -76.620 ;
        RECT -49.385 -78.660 -49.215 -76.620 ;
        RECT -48.205 -78.660 -48.035 -76.620 ;
        RECT -171.465 -79.760 -75.570 -79.460 ;
        RECT -171.465 -79.930 -75.075 -79.760 ;
        RECT -171.465 -80.110 -75.570 -79.930 ;
        RECT -75.245 -82.700 -75.075 -79.930 ;
        RECT -74.065 -82.700 -73.895 -80.660 ;
        RECT -72.885 -82.700 -72.715 -80.660 ;
        RECT -71.705 -82.700 -71.535 -80.660 ;
        RECT -70.525 -82.700 -70.355 -80.660 ;
        RECT -69.345 -82.700 -69.175 -80.660 ;
        RECT -68.165 -82.700 -67.995 -80.660 ;
        RECT -66.985 -82.700 -66.815 -80.660 ;
        RECT -65.805 -82.700 -65.635 -80.660 ;
        RECT -64.625 -82.700 -64.455 -80.660 ;
        RECT -63.445 -82.700 -63.275 -80.660 ;
        RECT -62.265 -82.700 -62.095 -80.660 ;
        RECT -61.085 -82.700 -60.915 -80.660 ;
        RECT -59.905 -82.700 -59.735 -80.660 ;
        RECT -58.725 -82.700 -58.555 -80.660 ;
        RECT -57.545 -82.700 -57.375 -80.660 ;
        RECT -56.365 -82.700 -56.195 -80.660 ;
      LAYER met1 ;
        RECT -56.495 -79.145 -56.265 -76.640 ;
        RECT -55.315 -79.145 -55.085 -76.640 ;
        RECT -54.135 -79.145 -53.905 -76.640 ;
        RECT -52.955 -79.145 -52.725 -76.640 ;
        RECT -51.775 -79.145 -51.545 -76.640 ;
        RECT -50.595 -79.145 -50.365 -76.640 ;
        RECT -49.415 -79.145 -49.185 -76.640 ;
        RECT -48.235 -79.145 -48.005 -76.640 ;
        RECT -56.495 -79.375 -48.005 -79.145 ;
        RECT -56.495 -79.955 -56.265 -79.375 ;
        RECT -75.420 -80.325 -56.035 -79.955 ;
        RECT -75.275 -82.680 -75.045 -80.325 ;
        RECT -74.095 -82.680 -73.865 -80.325 ;
        RECT -72.915 -82.680 -72.685 -80.325 ;
        RECT -71.735 -82.680 -71.505 -80.325 ;
        RECT -70.555 -82.680 -70.325 -80.325 ;
        RECT -69.375 -82.680 -69.145 -80.325 ;
        RECT -68.195 -82.680 -67.965 -80.325 ;
        RECT -67.015 -82.680 -66.785 -80.325 ;
        RECT -65.835 -82.680 -65.605 -80.325 ;
        RECT -64.655 -82.680 -64.425 -80.325 ;
        RECT -63.475 -82.680 -63.245 -80.325 ;
        RECT -62.295 -82.680 -62.065 -80.325 ;
        RECT -61.115 -82.680 -60.885 -80.325 ;
        RECT -59.935 -82.680 -59.705 -80.325 ;
        RECT -58.755 -82.680 -58.525 -80.325 ;
        RECT -57.575 -82.680 -57.345 -80.325 ;
        RECT -56.395 -82.680 -56.165 -80.325 ;
    END
  END DIV_OUT
  PIN VDD
    ANTENNAGATEAREA 14.000000 ;
    ANTENNADIFFAREA 3074.406982 ;
    PORT
      LAYER nwell ;
        RECT -55.705 599.615 -53.835 599.775 ;
        RECT -60.505 596.185 -53.835 599.615 ;
        RECT -60.505 595.750 -53.800 596.185 ;
        RECT -60.505 595.380 -52.830 595.750 ;
        RECT -58.480 594.290 -52.830 595.380 ;
        RECT -58.445 593.140 -52.830 594.290 ;
        RECT -58.445 591.865 -52.905 593.140 ;
        RECT -58.445 591.190 -52.685 591.865 ;
        RECT -58.480 590.755 -52.685 591.190 ;
        RECT -59.450 588.275 -52.685 590.755 ;
        RECT -59.450 588.145 -54.735 588.275 ;
        RECT -41.875 587.040 -37.510 594.425 ;
        RECT -55.550 581.275 -53.680 581.435 ;
        RECT -38.285 581.315 -36.415 581.475 ;
        RECT -60.350 577.845 -53.680 581.275 ;
        RECT -43.085 577.885 -36.415 581.315 ;
        RECT -60.350 577.410 -53.645 577.845 ;
        RECT -43.085 577.450 -36.380 577.885 ;
        RECT -60.350 577.040 -52.675 577.410 ;
        RECT -43.085 577.080 -35.410 577.450 ;
        RECT -58.325 575.950 -52.675 577.040 ;
        RECT -41.060 575.990 -35.410 577.080 ;
        RECT -58.290 574.800 -52.675 575.950 ;
        RECT -41.025 574.840 -35.410 575.990 ;
        RECT -58.290 573.525 -52.750 574.800 ;
        RECT -41.025 573.565 -35.485 574.840 ;
        RECT -58.290 572.850 -52.530 573.525 ;
        RECT -41.025 572.890 -35.265 573.565 ;
        RECT -58.325 572.415 -52.530 572.850 ;
        RECT -41.060 572.455 -35.265 572.890 ;
        RECT -59.295 569.935 -52.530 572.415 ;
        RECT -42.030 569.975 -35.265 572.455 ;
        RECT -59.295 569.805 -54.580 569.935 ;
        RECT -42.030 569.845 -37.315 569.975 ;
        RECT -55.895 552.795 -54.025 552.955 ;
        RECT -60.695 549.365 -54.025 552.795 ;
        RECT -60.695 548.930 -53.990 549.365 ;
        RECT -60.695 548.560 -53.020 548.930 ;
        RECT -58.670 547.470 -53.020 548.560 ;
        RECT -58.635 546.320 -53.020 547.470 ;
        RECT -58.635 545.045 -53.095 546.320 ;
        RECT -58.635 544.370 -52.875 545.045 ;
        RECT -58.670 543.935 -52.875 544.370 ;
        RECT -59.640 541.455 -52.875 543.935 ;
        RECT -59.640 541.325 -54.925 541.455 ;
        RECT -42.065 540.220 -37.700 547.605 ;
        RECT -55.740 534.455 -53.870 534.615 ;
        RECT -38.475 534.495 -36.605 534.655 ;
        RECT -60.540 531.025 -53.870 534.455 ;
        RECT -43.275 531.065 -36.605 534.495 ;
        RECT -60.540 530.590 -53.835 531.025 ;
        RECT -43.275 530.630 -36.570 531.065 ;
        RECT -60.540 530.220 -52.865 530.590 ;
        RECT -43.275 530.260 -35.600 530.630 ;
        RECT -58.515 529.130 -52.865 530.220 ;
        RECT -41.250 529.170 -35.600 530.260 ;
        RECT -58.480 527.980 -52.865 529.130 ;
        RECT -41.215 528.020 -35.600 529.170 ;
        RECT -58.480 526.705 -52.940 527.980 ;
        RECT -41.215 526.745 -35.675 528.020 ;
        RECT -58.480 526.030 -52.720 526.705 ;
        RECT -41.215 526.070 -35.455 526.745 ;
        RECT -58.515 525.595 -52.720 526.030 ;
        RECT -41.250 525.635 -35.455 526.070 ;
        RECT -59.485 523.115 -52.720 525.595 ;
        RECT -42.220 523.155 -35.455 525.635 ;
        RECT -59.485 522.985 -54.770 523.115 ;
        RECT -42.220 523.025 -37.505 523.155 ;
        RECT -55.980 507.030 -54.110 507.190 ;
        RECT -60.780 503.600 -54.110 507.030 ;
        RECT -60.780 503.165 -54.075 503.600 ;
        RECT -60.780 502.795 -53.105 503.165 ;
        RECT -58.755 501.705 -53.105 502.795 ;
        RECT -58.720 500.555 -53.105 501.705 ;
        RECT -58.720 499.280 -53.180 500.555 ;
        RECT -58.720 498.605 -52.960 499.280 ;
        RECT -58.755 498.170 -52.960 498.605 ;
        RECT -59.725 495.690 -52.960 498.170 ;
        RECT -59.725 495.560 -55.010 495.690 ;
        RECT -42.150 494.455 -37.785 501.840 ;
        RECT -55.825 488.690 -53.955 488.850 ;
        RECT -38.560 488.730 -36.690 488.890 ;
        RECT -60.625 485.260 -53.955 488.690 ;
        RECT -43.360 485.300 -36.690 488.730 ;
        RECT -60.625 484.825 -53.920 485.260 ;
        RECT -43.360 484.865 -36.655 485.300 ;
        RECT -60.625 484.455 -52.950 484.825 ;
        RECT -43.360 484.495 -35.685 484.865 ;
        RECT -58.600 483.365 -52.950 484.455 ;
        RECT -41.335 483.405 -35.685 484.495 ;
        RECT -58.565 482.215 -52.950 483.365 ;
        RECT -41.300 482.255 -35.685 483.405 ;
        RECT -58.565 480.940 -53.025 482.215 ;
        RECT -41.300 480.980 -35.760 482.255 ;
        RECT -58.565 480.265 -52.805 480.940 ;
        RECT -41.300 480.305 -35.540 480.980 ;
        RECT -58.600 479.830 -52.805 480.265 ;
        RECT -41.335 479.870 -35.540 480.305 ;
        RECT -59.570 477.350 -52.805 479.830 ;
        RECT -42.305 477.390 -35.540 479.870 ;
        RECT -59.570 477.220 -54.855 477.350 ;
        RECT -42.305 477.260 -37.590 477.390 ;
        RECT -56.310 463.260 -54.440 463.420 ;
        RECT -61.110 459.830 -54.440 463.260 ;
        RECT -61.110 459.395 -54.405 459.830 ;
        RECT -61.110 459.025 -53.435 459.395 ;
        RECT -59.085 457.935 -53.435 459.025 ;
        RECT -59.050 456.785 -53.435 457.935 ;
        RECT -59.050 455.510 -53.510 456.785 ;
        RECT -59.050 454.835 -53.290 455.510 ;
        RECT -59.085 454.400 -53.290 454.835 ;
        RECT -60.055 451.920 -53.290 454.400 ;
        RECT -60.055 451.790 -55.340 451.920 ;
        RECT -42.480 450.685 -38.115 458.070 ;
        RECT -56.155 444.920 -54.285 445.080 ;
        RECT -38.890 444.960 -37.020 445.120 ;
        RECT -60.955 441.490 -54.285 444.920 ;
        RECT -43.690 441.530 -37.020 444.960 ;
        RECT -60.955 441.055 -54.250 441.490 ;
        RECT -43.690 441.095 -36.985 441.530 ;
        RECT -60.955 440.685 -53.280 441.055 ;
        RECT -43.690 440.725 -36.015 441.095 ;
        RECT -58.930 439.595 -53.280 440.685 ;
        RECT -41.665 439.635 -36.015 440.725 ;
        RECT -58.895 438.445 -53.280 439.595 ;
        RECT -41.630 438.485 -36.015 439.635 ;
        RECT -58.895 437.170 -53.355 438.445 ;
        RECT -41.630 437.210 -36.090 438.485 ;
        RECT -58.895 436.495 -53.135 437.170 ;
        RECT -41.630 436.535 -35.870 437.210 ;
        RECT -58.930 436.060 -53.135 436.495 ;
        RECT -41.665 436.100 -35.870 436.535 ;
        RECT -59.900 433.580 -53.135 436.060 ;
        RECT -42.635 433.620 -35.870 436.100 ;
        RECT -59.900 433.450 -55.185 433.580 ;
        RECT -42.635 433.490 -37.920 433.620 ;
        RECT -56.480 417.270 -54.610 417.430 ;
        RECT -61.280 413.840 -54.610 417.270 ;
        RECT -61.280 413.405 -54.575 413.840 ;
        RECT -61.280 413.035 -53.605 413.405 ;
        RECT -59.255 411.945 -53.605 413.035 ;
        RECT -59.220 410.795 -53.605 411.945 ;
        RECT -59.220 409.520 -53.680 410.795 ;
        RECT -59.220 408.845 -53.460 409.520 ;
        RECT -59.255 408.410 -53.460 408.845 ;
        RECT -60.225 405.930 -53.460 408.410 ;
        RECT -60.225 405.800 -55.510 405.930 ;
        RECT -42.650 404.695 -38.285 412.080 ;
        RECT -56.325 398.930 -54.455 399.090 ;
        RECT -39.060 398.970 -37.190 399.130 ;
        RECT -61.125 395.500 -54.455 398.930 ;
        RECT -43.860 395.540 -37.190 398.970 ;
        RECT -61.125 395.065 -54.420 395.500 ;
        RECT -43.860 395.105 -37.155 395.540 ;
        RECT -61.125 394.695 -53.450 395.065 ;
        RECT -43.860 394.735 -36.185 395.105 ;
        RECT -59.100 393.605 -53.450 394.695 ;
        RECT -41.835 393.645 -36.185 394.735 ;
        RECT -59.065 392.455 -53.450 393.605 ;
        RECT -41.800 392.495 -36.185 393.645 ;
        RECT -59.065 391.180 -53.525 392.455 ;
        RECT -41.800 391.220 -36.260 392.495 ;
        RECT -59.065 390.505 -53.305 391.180 ;
        RECT -41.800 390.545 -36.040 391.220 ;
        RECT -59.100 390.070 -53.305 390.505 ;
        RECT -41.835 390.110 -36.040 390.545 ;
        RECT -60.070 387.590 -53.305 390.070 ;
        RECT -42.805 387.630 -36.040 390.110 ;
        RECT -60.070 387.460 -55.355 387.590 ;
        RECT -42.805 387.500 -38.090 387.630 ;
        RECT -56.285 372.955 -54.415 373.115 ;
        RECT -61.085 369.525 -54.415 372.955 ;
        RECT -61.085 369.090 -54.380 369.525 ;
        RECT -61.085 368.720 -53.410 369.090 ;
        RECT -59.060 367.630 -53.410 368.720 ;
        RECT -59.025 366.480 -53.410 367.630 ;
        RECT -59.025 365.205 -53.485 366.480 ;
        RECT -59.025 364.530 -53.265 365.205 ;
        RECT -59.060 364.095 -53.265 364.530 ;
        RECT -60.030 361.615 -53.265 364.095 ;
        RECT -60.030 361.485 -55.315 361.615 ;
        RECT -42.455 360.380 -38.090 367.765 ;
        RECT -56.130 354.615 -54.260 354.775 ;
        RECT -38.865 354.655 -36.995 354.815 ;
        RECT -60.930 351.185 -54.260 354.615 ;
        RECT -43.665 351.225 -36.995 354.655 ;
        RECT -60.930 350.750 -54.225 351.185 ;
        RECT -43.665 350.790 -36.960 351.225 ;
        RECT -60.930 350.380 -53.255 350.750 ;
        RECT -43.665 350.420 -35.990 350.790 ;
        RECT -58.905 349.290 -53.255 350.380 ;
        RECT -41.640 349.330 -35.990 350.420 ;
        RECT -58.870 348.140 -53.255 349.290 ;
        RECT -41.605 348.180 -35.990 349.330 ;
        RECT -58.870 346.865 -53.330 348.140 ;
        RECT -41.605 346.905 -36.065 348.180 ;
        RECT -58.870 346.190 -53.110 346.865 ;
        RECT -41.605 346.230 -35.845 346.905 ;
        RECT -58.905 345.755 -53.110 346.190 ;
        RECT -41.640 345.795 -35.845 346.230 ;
        RECT -59.875 343.275 -53.110 345.755 ;
        RECT -42.610 343.315 -35.845 345.795 ;
        RECT -59.875 343.145 -55.160 343.275 ;
        RECT -42.610 343.185 -37.895 343.315 ;
        RECT -56.230 330.755 -54.360 330.915 ;
        RECT -61.030 327.325 -54.360 330.755 ;
        RECT -61.030 326.890 -54.325 327.325 ;
        RECT -61.030 326.520 -53.355 326.890 ;
        RECT -59.005 325.430 -53.355 326.520 ;
        RECT -58.970 324.280 -53.355 325.430 ;
        RECT -58.970 323.005 -53.430 324.280 ;
        RECT -58.970 322.330 -53.210 323.005 ;
        RECT -59.005 321.895 -53.210 322.330 ;
        RECT -59.975 319.415 -53.210 321.895 ;
        RECT -59.975 319.285 -55.260 319.415 ;
        RECT -42.400 318.180 -38.035 325.565 ;
        RECT -56.075 312.415 -54.205 312.575 ;
        RECT -38.810 312.455 -36.940 312.615 ;
        RECT -60.875 308.985 -54.205 312.415 ;
        RECT -43.610 309.025 -36.940 312.455 ;
        RECT -60.875 308.550 -54.170 308.985 ;
        RECT -43.610 308.590 -36.905 309.025 ;
        RECT -60.875 308.180 -53.200 308.550 ;
        RECT -43.610 308.220 -35.935 308.590 ;
        RECT -58.850 307.090 -53.200 308.180 ;
        RECT -41.585 307.130 -35.935 308.220 ;
        RECT -58.815 305.940 -53.200 307.090 ;
        RECT -41.550 305.980 -35.935 307.130 ;
        RECT -58.815 304.665 -53.275 305.940 ;
        RECT -41.550 304.705 -36.010 305.980 ;
        RECT -58.815 303.990 -53.055 304.665 ;
        RECT -41.550 304.030 -35.790 304.705 ;
        RECT -58.850 303.555 -53.055 303.990 ;
        RECT -41.585 303.595 -35.790 304.030 ;
        RECT -59.820 301.075 -53.055 303.555 ;
        RECT -42.555 301.115 -35.790 303.595 ;
        RECT -59.820 300.945 -55.105 301.075 ;
        RECT -42.555 300.985 -37.840 301.115 ;
        RECT -57.715 276.200 -52.555 289.830 ;
        RECT -46.415 275.935 -44.145 289.615 ;
        RECT -39.175 276.045 -36.905 289.550 ;
        RECT -57.675 271.800 -55.410 274.900 ;
        RECT -46.410 274.660 -44.145 275.935 ;
        RECT -50.525 272.050 -44.145 274.660 ;
        RECT -47.755 271.995 -44.145 272.050 ;
        RECT -57.735 269.630 -55.445 269.785 ;
        RECT -57.740 262.505 -55.445 269.630 ;
        RECT -46.410 264.550 -44.145 271.995 ;
        RECT -39.205 275.870 -36.905 276.045 ;
        RECT -39.205 271.840 -36.910 275.870 ;
        RECT -46.410 262.845 -44.090 264.550 ;
        RECT -39.175 264.240 -36.910 271.840 ;
        RECT -57.680 257.925 -54.275 261.100 ;
        RECT -46.410 257.945 -44.145 262.845 ;
        RECT -57.680 253.195 -54.275 256.370 ;
        RECT -46.410 253.220 -41.545 257.945 ;
        RECT -46.410 253.215 -44.145 253.220 ;
        RECT -69.195 235.405 -66.925 248.910 ;
        RECT -69.195 235.230 -66.895 235.405 ;
        RECT -69.190 231.200 -66.895 235.230 ;
        RECT -61.955 235.295 -59.685 248.975 ;
        RECT -69.190 223.600 -66.925 231.200 ;
        RECT -61.955 223.910 -59.690 235.295 ;
        RECT -62.010 222.205 -59.690 223.910 ;
        RECT -61.955 219.185 -59.690 222.205 ;
        RECT -70.115 194.100 -67.740 203.685 ;
        RECT -70.115 194.095 -68.105 194.100 ;
        RECT -70.115 179.100 -67.740 188.685 ;
        RECT -58.860 184.110 -56.485 203.735 ;
        RECT -37.925 184.110 -35.550 203.735 ;
        RECT -26.670 194.100 -24.295 203.685 ;
        RECT -26.305 194.095 -24.295 194.100 ;
        RECT -58.860 181.500 -55.915 184.110 ;
        RECT -38.495 181.500 -35.550 184.110 ;
        RECT -58.860 181.065 -56.885 181.500 ;
        RECT -37.525 181.065 -35.550 181.500 ;
        RECT -70.115 179.095 -68.105 179.100 ;
        RECT -70.115 166.600 -67.740 176.185 ;
        RECT -58.860 176.085 -56.920 181.065 ;
        RECT -37.490 176.085 -35.550 181.065 ;
        RECT -26.670 179.100 -24.295 188.685 ;
        RECT -26.305 179.095 -24.295 179.100 ;
        RECT -58.860 173.475 -55.925 176.085 ;
        RECT -38.485 173.475 -35.550 176.085 ;
        RECT -58.860 173.040 -56.895 173.475 ;
        RECT -37.515 173.040 -35.550 173.475 ;
        RECT -58.860 168.065 -56.930 173.040 ;
        RECT -37.480 168.065 -35.550 173.040 ;
        RECT -70.115 166.595 -68.105 166.600 ;
        RECT -70.115 154.100 -67.740 163.685 ;
        RECT -58.860 158.135 -56.495 168.065 ;
        RECT -37.915 158.135 -35.550 168.065 ;
        RECT -26.670 166.600 -24.295 176.185 ;
        RECT -26.305 166.595 -24.295 166.600 ;
        RECT -58.860 156.705 -56.580 158.135 ;
        RECT -37.830 156.705 -35.550 158.135 ;
        RECT -58.860 155.000 -56.525 156.705 ;
        RECT -70.115 154.095 -68.105 154.100 ;
        RECT -70.115 141.600 -67.740 151.185 ;
        RECT -70.115 141.595 -68.105 141.600 ;
        RECT -70.115 129.100 -67.740 138.685 ;
        RECT -58.860 129.935 -56.580 155.000 ;
        RECT -51.610 147.710 -49.345 155.310 ;
        RECT -51.640 143.680 -49.345 147.710 ;
        RECT -45.065 147.710 -42.800 155.310 ;
        RECT -37.885 155.000 -35.550 156.705 ;
        RECT -45.065 143.680 -42.770 147.710 ;
        RECT -51.640 143.505 -49.340 143.680 ;
        RECT -51.610 130.000 -49.340 143.505 ;
        RECT -45.070 143.505 -42.770 143.680 ;
        RECT -45.070 130.000 -42.800 143.505 ;
        RECT -37.830 129.935 -35.550 155.000 ;
        RECT -26.670 154.100 -24.295 163.685 ;
        RECT -26.305 154.095 -24.295 154.100 ;
        RECT -26.670 141.600 -24.295 151.185 ;
        RECT -26.305 141.595 -24.295 141.600 ;
        RECT -33.960 131.285 -31.695 134.385 ;
        RECT -26.670 129.100 -24.295 138.685 ;
        RECT -70.115 129.095 -68.105 129.100 ;
        RECT -26.305 129.095 -24.295 129.100 ;
        RECT -52.360 122.085 -47.975 126.320 ;
        RECT -27.690 121.950 -23.305 126.185 ;
        RECT -57.510 117.335 -55.245 120.355 ;
        RECT -32.875 117.335 -30.610 120.355 ;
        RECT -57.510 115.630 -55.190 117.335 ;
        RECT -57.510 104.245 -55.245 115.630 ;
        RECT -50.275 108.340 -48.010 115.940 ;
        RECT -57.515 90.565 -55.245 104.245 ;
        RECT -50.305 104.310 -48.010 108.340 ;
        RECT -32.875 115.630 -30.555 117.335 ;
        RECT -43.870 107.225 -42.000 107.385 ;
        RECT -50.305 104.135 -48.005 104.310 ;
        RECT -50.275 90.630 -48.005 104.135 ;
        RECT -43.870 103.795 -37.200 107.225 ;
        RECT -32.875 104.245 -30.610 115.630 ;
        RECT -25.640 108.340 -23.375 115.940 ;
        RECT -43.905 103.360 -37.200 103.795 ;
        RECT -44.875 102.990 -37.200 103.360 ;
        RECT -44.875 101.900 -39.225 102.990 ;
        RECT -44.875 100.750 -39.260 101.900 ;
        RECT -44.800 99.475 -39.260 100.750 ;
        RECT -45.020 98.800 -39.260 99.475 ;
        RECT -45.020 98.365 -39.225 98.800 ;
        RECT -45.020 95.885 -38.255 98.365 ;
        RECT -42.970 95.755 -38.255 95.885 ;
        RECT -32.880 90.565 -30.610 104.245 ;
        RECT -25.670 104.310 -23.375 108.340 ;
        RECT -25.670 104.135 -23.370 104.310 ;
        RECT -25.640 90.630 -23.370 104.135 ;
        RECT -63.990 82.280 -62.120 82.440 ;
        RECT -38.990 82.280 -37.120 82.440 ;
        RECT -63.990 78.850 -57.320 82.280 ;
        RECT -38.990 78.850 -32.320 82.280 ;
        RECT -64.025 78.415 -57.320 78.850 ;
        RECT -39.025 78.415 -32.320 78.850 ;
        RECT -64.995 78.045 -57.320 78.415 ;
        RECT -39.995 78.045 -32.320 78.415 ;
        RECT -64.995 76.955 -59.345 78.045 ;
        RECT -39.995 76.955 -34.345 78.045 ;
        RECT -64.995 75.805 -59.380 76.955 ;
        RECT -39.995 75.805 -34.380 76.955 ;
        RECT -64.920 74.530 -59.380 75.805 ;
        RECT -39.920 74.530 -34.380 75.805 ;
        RECT -65.140 73.855 -59.380 74.530 ;
        RECT -40.140 73.855 -34.380 74.530 ;
        RECT -65.140 73.420 -59.345 73.855 ;
        RECT -40.140 73.420 -34.345 73.855 ;
        RECT -65.140 70.940 -58.375 73.420 ;
        RECT -40.140 70.940 -33.375 73.420 ;
        RECT -63.090 70.810 -58.375 70.940 ;
        RECT -38.090 70.810 -33.375 70.940 ;
        RECT -39.255 68.910 -36.965 69.065 ;
        RECT -56.350 63.800 -52.945 66.975 ;
        RECT -56.345 59.275 -52.940 62.450 ;
        RECT -39.255 61.785 -36.960 68.910 ;
        RECT -29.680 65.675 -27.810 69.265 ;
        RECT -29.715 65.240 -27.810 65.675 ;
        RECT -30.685 62.630 -27.810 65.240 ;
        RECT -29.575 59.760 -27.285 59.915 ;
        RECT -70.465 51.715 -68.170 58.840 ;
        RECT -57.700 53.245 -52.975 57.970 ;
        RECT -39.225 55.965 -37.355 59.555 ;
        RECT -39.260 55.530 -37.355 55.965 ;
        RECT -40.230 52.920 -37.355 55.530 ;
        RECT -29.575 52.635 -27.280 59.760 ;
        RECT -70.460 51.560 -68.170 51.715 ;
        RECT 72.345 45.265 79.750 51.075 ;
        RECT 78.320 44.030 79.740 45.265 ;
        RECT 40.480 33.170 63.825 39.595 ;
        RECT 40.950 32.945 63.570 33.170 ;
        RECT 98.730 15.580 110.780 18.060 ;
        RECT 211.800 15.630 225.480 15.635 ;
        RECT 195.690 13.365 225.480 15.630 ;
        RECT 198.710 13.310 200.415 13.365 ;
        RECT 254.240 12.860 292.240 16.705 ;
        RECT -67.285 7.565 -29.285 11.410 ;
        RECT -18.160 8.875 -6.110 11.355 ;
        RECT 22.335 9.755 34.385 12.235 ;
        RECT 8.585 9.415 9.605 9.635 ;
        RECT 2.885 9.405 4.565 9.415 ;
        RECT 8.585 9.405 14.895 9.415 ;
        RECT -13.910 2.640 -6.110 5.120 ;
        RECT 2.885 4.905 14.895 9.405 ;
        RECT 37.850 8.975 75.850 12.820 ;
        RECT 102.980 9.345 110.780 11.825 ;
        RECT 140.305 10.620 146.350 11.910 ;
        RECT 140.305 10.265 147.785 10.620 ;
        RECT 138.365 7.030 147.785 10.265 ;
        RECT 164.580 10.585 170.625 11.875 ;
        RECT 164.580 10.230 172.060 10.585 ;
        RECT 146.345 7.025 147.785 7.030 ;
        RECT 2.885 4.895 4.565 4.905 ;
        RECT 8.585 4.895 14.895 4.905 ;
        RECT 8.585 4.675 9.605 4.895 ;
        RECT 26.585 3.520 34.385 6.000 ;
        RECT 151.410 1.890 158.380 9.510 ;
        RECT 162.640 6.995 172.060 10.230 ;
        RECT 170.620 6.990 172.060 6.995 ;
        RECT 175.085 2.005 182.055 9.620 ;
        RECT 183.690 2.220 190.660 9.405 ;
        RECT 207.705 8.395 211.910 8.425 ;
        RECT 200.105 6.130 225.415 8.395 ;
        RECT 227.655 6.580 230.755 8.845 ;
        RECT 211.735 6.125 225.415 6.130 ;
        RECT -25.500 -2.985 -13.450 -0.505 ;
        RECT 22.410 -3.695 34.460 -1.215 ;
        RECT 37.645 -4.805 75.645 -0.960 ;
        RECT 99.590 -1.170 111.640 1.310 ;
        RECT 253.225 -1.695 291.225 2.150 ;
        RECT -21.250 -9.220 -13.450 -6.740 ;
        RECT 103.840 -7.405 111.640 -4.925 ;
        RECT 26.660 -9.930 34.460 -7.450 ;
        RECT 253.225 -16.930 291.225 -13.085 ;
        RECT 311.725 -15.500 323.775 -13.020 ;
        RECT 315.975 -21.735 323.775 -19.255 ;
        RECT -75.485 -84.215 -37.485 -80.370 ;
        RECT -75.935 -91.030 -62.255 -91.025 ;
        RECT -75.935 -93.295 -50.625 -91.030 ;
        RECT -62.430 -93.325 -58.225 -93.295 ;
        RECT -113.930 -94.940 -106.805 -94.935 ;
        RECT -113.930 -97.230 -106.650 -94.940 ;
        RECT -44.615 -95.345 -40.380 -90.960 ;
        RECT -37.470 -93.960 -27.880 -91.950 ;
        RECT -24.970 -93.960 -15.380 -91.950 ;
        RECT -12.470 -93.960 -2.880 -91.950 ;
        RECT 0.030 -93.960 9.620 -91.950 ;
        RECT 12.530 -93.960 22.120 -91.950 ;
        RECT 27.530 -93.960 37.120 -91.950 ;
        RECT -37.465 -94.325 -27.880 -93.960 ;
        RECT -24.965 -94.325 -15.380 -93.960 ;
        RECT -12.465 -94.325 -2.880 -93.960 ;
        RECT 0.035 -94.325 9.620 -93.960 ;
        RECT 12.535 -94.325 22.120 -93.960 ;
        RECT 27.535 -94.325 37.120 -93.960 ;
        RECT -103.935 -97.335 -97.300 -95.465 ;
        RECT -103.935 -97.370 -100.890 -97.335 ;
        RECT -103.935 -98.340 -101.325 -97.370 ;
        RECT -50.935 -98.265 -49.230 -98.210 ;
        RECT -95.755 -102.000 -93.145 -101.030 ;
        RECT -88.520 -102.000 -84.285 -99.975 ;
        RECT -76.000 -100.530 -46.210 -98.265 ;
        RECT -76.000 -100.535 -62.320 -100.530 ;
        RECT -35.280 -101.615 -32.180 -99.350 ;
        RECT -95.755 -102.035 -92.710 -102.000 ;
        RECT -89.610 -102.035 -84.285 -102.000 ;
        RECT -104.780 -104.620 -97.655 -104.615 ;
        RECT -113.645 -106.880 -107.010 -105.010 ;
        RECT -113.645 -106.915 -110.600 -106.880 ;
        RECT -104.780 -106.910 -97.500 -104.620 ;
        RECT -95.755 -104.775 -84.285 -102.035 ;
        RECT -95.755 -105.745 -84.125 -104.775 ;
        RECT -95.625 -106.645 -84.125 -105.745 ;
        RECT -95.625 -106.680 -87.715 -106.645 ;
        RECT -113.645 -107.885 -111.035 -106.915 ;
        RECT -95.625 -107.575 -88.150 -106.680 ;
        RECT -95.625 -107.795 -92.035 -107.575 ;
        RECT -90.760 -107.650 -88.150 -107.575 ;
        RECT -70.810 -106.880 -68.200 -105.910 ;
        RECT -63.575 -106.880 -59.340 -104.855 ;
        RECT -36.630 -105.135 37.170 -103.205 ;
        RECT 310.825 -103.415 314.415 -103.195 ;
        RECT 356.590 -103.330 360.180 -103.110 ;
        RECT 403.410 -103.140 407.000 -102.920 ;
        RECT 408.275 -103.140 410.885 -103.065 ;
        RECT 361.455 -103.330 364.065 -103.255 ;
        RECT 315.690 -103.415 318.300 -103.340 ;
        RECT 134.550 -103.665 138.140 -103.445 ;
        RECT 139.415 -103.665 142.025 -103.590 ;
        RECT 134.550 -104.560 142.025 -103.665 ;
        RECT 176.750 -103.720 180.340 -103.500 ;
        RECT 181.615 -103.720 184.225 -103.645 ;
        RECT 109.305 -104.565 122.985 -104.560 ;
        RECT -36.630 -105.485 1.500 -105.135 ;
        RECT 6.475 -105.145 37.170 -105.135 ;
        RECT 6.475 -105.170 9.520 -105.145 ;
        RECT -11.565 -105.540 -9.860 -105.485 ;
        RECT -8.430 -105.570 1.500 -105.485 ;
        RECT 6.910 -106.140 9.520 -105.170 ;
        RECT 14.500 -105.180 37.170 -105.145 ;
        RECT 14.935 -105.580 37.170 -105.180 ;
        RECT 14.935 -106.150 17.545 -105.580 ;
        RECT 97.675 -106.830 122.985 -104.565 ;
        RECT 134.550 -104.595 142.460 -104.560 ;
        RECT 134.550 -105.495 146.050 -104.595 ;
        RECT 134.420 -106.465 146.050 -105.495 ;
        RECT 176.750 -104.615 184.225 -103.720 ;
        RECT 221.065 -103.915 224.655 -103.695 ;
        RECT 267.055 -103.745 270.645 -103.525 ;
        RECT 271.920 -103.745 274.530 -103.670 ;
        RECT 225.930 -103.915 228.540 -103.840 ;
        RECT 176.750 -104.650 184.660 -104.615 ;
        RECT 176.750 -105.550 188.250 -104.650 ;
        RECT 105.275 -106.860 109.480 -106.830 ;
        RECT -70.810 -106.915 -67.765 -106.880 ;
        RECT -64.665 -106.915 -59.340 -106.880 ;
        RECT -70.810 -109.655 -59.340 -106.915 ;
        RECT -70.810 -110.625 -59.180 -109.655 ;
        RECT -23.060 -110.455 -18.855 -110.425 ;
        RECT -70.680 -111.525 -59.180 -110.625 ;
        RECT -70.680 -111.560 -62.770 -111.525 ;
        RECT -70.680 -112.455 -63.205 -111.560 ;
        RECT -70.680 -112.675 -67.090 -112.455 ;
        RECT -65.815 -112.530 -63.205 -112.455 ;
        RECT -36.565 -112.720 -11.255 -110.455 ;
        RECT 86.655 -111.800 91.380 -109.200 ;
        RECT 134.420 -109.205 145.890 -106.465 ;
        RECT 134.420 -109.240 137.465 -109.205 ;
        RECT 140.565 -109.240 145.890 -109.205 ;
        RECT 134.420 -110.210 137.030 -109.240 ;
        RECT 141.655 -111.265 145.890 -109.240 ;
        RECT 151.615 -110.055 159.000 -105.690 ;
        RECT 176.620 -106.520 188.250 -105.550 ;
        RECT 221.065 -104.810 228.540 -103.915 ;
        RECT 267.055 -104.640 274.530 -103.745 ;
        RECT 310.825 -104.310 318.300 -103.415 ;
        RECT 356.590 -104.225 364.065 -103.330 ;
        RECT 403.410 -104.035 410.885 -103.140 ;
        RECT 403.410 -104.070 411.320 -104.035 ;
        RECT 356.590 -104.260 364.500 -104.225 ;
        RECT 310.825 -104.345 318.735 -104.310 ;
        RECT 267.055 -104.675 274.965 -104.640 ;
        RECT 221.065 -104.845 228.975 -104.810 ;
        RECT 221.065 -105.745 232.565 -104.845 ;
        RECT 267.055 -105.575 278.555 -104.675 ;
        RECT 310.825 -105.245 322.325 -104.345 ;
        RECT 356.590 -105.160 368.090 -104.260 ;
        RECT 403.410 -104.970 414.910 -104.070 ;
        RECT 176.620 -109.260 188.090 -106.520 ;
        RECT 176.620 -109.295 179.665 -109.260 ;
        RECT 182.765 -109.295 188.090 -109.260 ;
        RECT 176.620 -110.265 179.230 -109.295 ;
        RECT 183.855 -111.320 188.090 -109.295 ;
        RECT 193.815 -110.110 201.200 -105.745 ;
        RECT 220.935 -106.715 232.565 -105.745 ;
        RECT 220.935 -109.455 232.405 -106.715 ;
        RECT 220.935 -109.490 223.980 -109.455 ;
        RECT 227.080 -109.490 232.405 -109.455 ;
        RECT 220.935 -110.460 223.545 -109.490 ;
        RECT 228.170 -111.515 232.405 -109.490 ;
        RECT 238.130 -110.305 245.515 -105.940 ;
        RECT 266.925 -106.545 278.555 -105.575 ;
        RECT 266.925 -109.285 278.395 -106.545 ;
        RECT 266.925 -109.320 269.970 -109.285 ;
        RECT 273.070 -109.320 278.395 -109.285 ;
        RECT 266.925 -110.290 269.535 -109.320 ;
        RECT 274.160 -111.345 278.395 -109.320 ;
        RECT 284.120 -110.135 291.505 -105.770 ;
        RECT 310.695 -106.215 322.325 -105.245 ;
        RECT 310.695 -108.955 322.165 -106.215 ;
        RECT 310.695 -108.990 313.740 -108.955 ;
        RECT 316.840 -108.990 322.165 -108.955 ;
        RECT 310.695 -109.960 313.305 -108.990 ;
        RECT 317.930 -111.015 322.165 -108.990 ;
        RECT 327.890 -109.805 335.275 -105.440 ;
        RECT 356.460 -106.130 368.090 -105.160 ;
        RECT 356.460 -108.870 367.930 -106.130 ;
        RECT 356.460 -108.905 359.505 -108.870 ;
        RECT 362.605 -108.905 367.930 -108.870 ;
        RECT 356.460 -109.875 359.070 -108.905 ;
        RECT 363.695 -110.930 367.930 -108.905 ;
        RECT 373.655 -109.720 381.040 -105.355 ;
        RECT 403.280 -105.940 414.910 -104.970 ;
        RECT 403.280 -108.680 414.750 -105.940 ;
        RECT 403.280 -108.715 406.325 -108.680 ;
        RECT 409.425 -108.715 414.750 -108.680 ;
        RECT 403.280 -109.685 405.890 -108.715 ;
        RECT 410.515 -110.740 414.750 -108.715 ;
        RECT 420.475 -109.530 427.860 -105.165 ;
        RECT 96.280 -111.800 97.985 -111.745 ;
        RECT -36.565 -112.725 -22.885 -112.720 ;
        RECT 86.650 -114.065 123.050 -111.800 ;
        RECT 105.430 -115.410 108.095 -114.065 ;
        RECT 109.370 -114.070 123.050 -114.065 ;
        RECT -75.935 -115.665 -62.255 -115.660 ;
        RECT -75.935 -117.930 -50.625 -115.665 ;
        RECT -62.430 -117.960 -58.225 -117.930 ;
        RECT -44.480 -120.015 -40.245 -115.630 ;
        RECT -36.565 -117.000 -22.885 -116.995 ;
        RECT -36.565 -119.265 -11.255 -117.000 ;
        RECT 105.485 -118.180 108.095 -115.410 ;
        RECT -23.060 -119.295 -18.855 -119.265 ;
        RECT -113.320 -125.355 -108.595 -120.630 ;
        RECT -107.290 -124.000 -104.115 -120.595 ;
        RECT -102.765 -124.005 -99.590 -120.600 ;
        RECT -50.935 -122.900 -49.230 -122.845 ;
        RECT -95.755 -127.000 -93.145 -126.030 ;
        RECT -88.520 -127.000 -84.285 -124.975 ;
        RECT -76.000 -125.165 -46.210 -122.900 ;
        RECT -11.565 -124.235 -9.860 -124.180 ;
        RECT -8.430 -124.235 1.500 -124.150 ;
        RECT -36.630 -124.585 1.500 -124.235 ;
        RECT 6.910 -124.550 9.520 -123.580 ;
        RECT 14.935 -124.140 17.545 -123.570 ;
        RECT 14.935 -124.540 37.170 -124.140 ;
        RECT 6.475 -124.575 9.520 -124.550 ;
        RECT 14.500 -124.575 37.170 -124.540 ;
        RECT 6.475 -124.585 37.170 -124.575 ;
        RECT -76.000 -125.170 -62.320 -125.165 ;
        RECT -36.630 -126.515 37.170 -124.585 ;
        RECT 86.630 -125.335 89.805 -121.930 ;
        RECT 91.360 -125.335 94.535 -121.930 ;
        RECT 95.940 -125.390 103.220 -123.100 ;
        RECT 105.235 -125.330 108.335 -123.065 ;
        RECT 109.635 -125.370 123.265 -120.210 ;
        RECT 310.785 -120.680 314.375 -120.460 ;
        RECT 356.550 -120.595 360.140 -120.375 ;
        RECT 403.370 -120.405 406.960 -120.185 ;
        RECT 408.235 -120.405 410.845 -120.330 ;
        RECT 361.415 -120.595 364.025 -120.520 ;
        RECT 315.650 -120.680 318.260 -120.605 ;
        RECT 134.510 -120.930 138.100 -120.710 ;
        RECT 139.375 -120.930 141.985 -120.855 ;
        RECT 134.510 -121.825 141.985 -120.930 ;
        RECT 152.850 -121.085 156.440 -120.865 ;
        RECT 176.710 -120.985 180.300 -120.765 ;
        RECT 181.575 -120.985 184.185 -120.910 ;
        RECT 157.715 -121.085 160.325 -121.010 ;
        RECT 134.510 -121.860 142.420 -121.825 ;
        RECT 134.510 -122.760 146.010 -121.860 ;
        RECT 134.380 -123.730 146.010 -122.760 ;
        RECT 152.850 -121.980 160.325 -121.085 ;
        RECT 176.710 -121.880 184.185 -120.985 ;
        RECT 195.050 -121.140 198.640 -120.920 ;
        RECT 199.915 -121.140 202.525 -121.065 ;
        RECT 176.710 -121.915 184.620 -121.880 ;
        RECT 152.850 -122.015 160.760 -121.980 ;
        RECT 152.850 -122.915 164.350 -122.015 ;
        RECT 176.710 -122.815 188.210 -121.915 ;
        RECT 95.940 -125.395 103.065 -125.390 ;
        RECT 134.380 -126.470 145.850 -123.730 ;
        RECT 134.380 -126.505 137.425 -126.470 ;
        RECT 140.525 -126.505 145.850 -126.470 ;
        RECT -95.755 -127.035 -92.710 -127.000 ;
        RECT -89.610 -127.035 -84.285 -127.000 ;
        RECT -95.755 -129.775 -84.285 -127.035 ;
        RECT 68.730 -127.345 82.410 -127.340 ;
        RECT 52.620 -129.610 82.410 -127.345 ;
        RECT 134.380 -127.475 136.990 -126.505 ;
        RECT 141.615 -128.530 145.850 -126.505 ;
        RECT 152.720 -123.885 164.350 -122.915 ;
        RECT 176.580 -123.785 188.210 -122.815 ;
        RECT 195.050 -122.035 202.525 -121.140 ;
        RECT 221.025 -121.180 224.615 -120.960 ;
        RECT 267.015 -121.010 270.605 -120.790 ;
        RECT 271.880 -121.010 274.490 -120.935 ;
        RECT 225.890 -121.180 228.500 -121.105 ;
        RECT 195.050 -122.070 202.960 -122.035 ;
        RECT 195.050 -122.970 206.550 -122.070 ;
        RECT 152.720 -126.625 164.190 -123.885 ;
        RECT 152.720 -126.660 155.765 -126.625 ;
        RECT 158.865 -126.660 164.190 -126.625 ;
        RECT 152.720 -127.630 155.330 -126.660 ;
        RECT 159.955 -128.685 164.190 -126.660 ;
        RECT 176.580 -126.525 188.050 -123.785 ;
        RECT 176.580 -126.560 179.625 -126.525 ;
        RECT 182.725 -126.560 188.050 -126.525 ;
        RECT 176.580 -127.530 179.190 -126.560 ;
        RECT 183.815 -128.585 188.050 -126.560 ;
        RECT 194.920 -123.940 206.550 -122.970 ;
        RECT 221.025 -122.075 228.500 -121.180 ;
        RECT 239.365 -121.335 242.955 -121.115 ;
        RECT 244.230 -121.335 246.840 -121.260 ;
        RECT 221.025 -122.110 228.935 -122.075 ;
        RECT 221.025 -123.010 232.525 -122.110 ;
        RECT 194.920 -126.680 206.390 -123.940 ;
        RECT 194.920 -126.715 197.965 -126.680 ;
        RECT 201.065 -126.715 206.390 -126.680 ;
        RECT 194.920 -127.685 197.530 -126.715 ;
        RECT 202.155 -128.740 206.390 -126.715 ;
        RECT 220.895 -123.980 232.525 -123.010 ;
        RECT 239.365 -122.230 246.840 -121.335 ;
        RECT 267.015 -121.905 274.490 -121.010 ;
        RECT 285.355 -121.165 288.945 -120.945 ;
        RECT 290.220 -121.165 292.830 -121.090 ;
        RECT 267.015 -121.940 274.925 -121.905 ;
        RECT 239.365 -122.265 247.275 -122.230 ;
        RECT 239.365 -123.165 250.865 -122.265 ;
        RECT 267.015 -122.840 278.515 -121.940 ;
        RECT 220.895 -126.720 232.365 -123.980 ;
        RECT 220.895 -126.755 223.940 -126.720 ;
        RECT 227.040 -126.755 232.365 -126.720 ;
        RECT 220.895 -127.725 223.505 -126.755 ;
        RECT 228.130 -128.780 232.365 -126.755 ;
        RECT 239.235 -124.135 250.865 -123.165 ;
        RECT 266.885 -123.810 278.515 -122.840 ;
        RECT 285.355 -122.060 292.830 -121.165 ;
        RECT 310.785 -121.575 318.260 -120.680 ;
        RECT 329.125 -120.835 332.715 -120.615 ;
        RECT 333.990 -120.835 336.600 -120.760 ;
        RECT 310.785 -121.610 318.695 -121.575 ;
        RECT 285.355 -122.095 293.265 -122.060 ;
        RECT 285.355 -122.995 296.855 -122.095 ;
        RECT 310.785 -122.510 322.285 -121.610 ;
        RECT 239.235 -126.875 250.705 -124.135 ;
        RECT 239.235 -126.910 242.280 -126.875 ;
        RECT 245.380 -126.910 250.705 -126.875 ;
        RECT 239.235 -127.880 241.845 -126.910 ;
        RECT 246.470 -128.935 250.705 -126.910 ;
        RECT 266.885 -126.550 278.355 -123.810 ;
        RECT 266.885 -126.585 269.930 -126.550 ;
        RECT 273.030 -126.585 278.355 -126.550 ;
        RECT 266.885 -127.555 269.495 -126.585 ;
        RECT 274.120 -128.610 278.355 -126.585 ;
        RECT 285.225 -123.965 296.855 -122.995 ;
        RECT 310.655 -123.480 322.285 -122.510 ;
        RECT 329.125 -121.730 336.600 -120.835 ;
        RECT 356.550 -121.490 364.025 -120.595 ;
        RECT 374.890 -120.750 378.480 -120.530 ;
        RECT 379.755 -120.750 382.365 -120.675 ;
        RECT 356.550 -121.525 364.460 -121.490 ;
        RECT 329.125 -121.765 337.035 -121.730 ;
        RECT 329.125 -122.665 340.625 -121.765 ;
        RECT 356.550 -122.425 368.050 -121.525 ;
        RECT 285.225 -126.705 296.695 -123.965 ;
        RECT 285.225 -126.740 288.270 -126.705 ;
        RECT 291.370 -126.740 296.695 -126.705 ;
        RECT 285.225 -127.710 287.835 -126.740 ;
        RECT 292.460 -128.765 296.695 -126.740 ;
        RECT 310.655 -126.220 322.125 -123.480 ;
        RECT 310.655 -126.255 313.700 -126.220 ;
        RECT 316.800 -126.255 322.125 -126.220 ;
        RECT 310.655 -127.225 313.265 -126.255 ;
        RECT 317.890 -128.280 322.125 -126.255 ;
        RECT 328.995 -123.635 340.625 -122.665 ;
        RECT 356.420 -123.395 368.050 -122.425 ;
        RECT 374.890 -121.645 382.365 -120.750 ;
        RECT 403.370 -121.300 410.845 -120.405 ;
        RECT 421.710 -120.560 425.300 -120.340 ;
        RECT 426.575 -120.560 429.185 -120.485 ;
        RECT 403.370 -121.335 411.280 -121.300 ;
        RECT 374.890 -121.680 382.800 -121.645 ;
        RECT 374.890 -122.580 386.390 -121.680 ;
        RECT 403.370 -122.235 414.870 -121.335 ;
        RECT 328.995 -126.375 340.465 -123.635 ;
        RECT 328.995 -126.410 332.040 -126.375 ;
        RECT 335.140 -126.410 340.465 -126.375 ;
        RECT 328.995 -127.380 331.605 -126.410 ;
        RECT 336.230 -128.435 340.465 -126.410 ;
        RECT 356.420 -126.135 367.890 -123.395 ;
        RECT 356.420 -126.170 359.465 -126.135 ;
        RECT 362.565 -126.170 367.890 -126.135 ;
        RECT 356.420 -127.140 359.030 -126.170 ;
        RECT 363.655 -128.195 367.890 -126.170 ;
        RECT 374.760 -123.550 386.390 -122.580 ;
        RECT 403.240 -123.205 414.870 -122.235 ;
        RECT 421.710 -121.455 429.185 -120.560 ;
        RECT 421.710 -121.490 429.620 -121.455 ;
        RECT 421.710 -122.390 433.210 -121.490 ;
        RECT 374.760 -126.290 386.230 -123.550 ;
        RECT 374.760 -126.325 377.805 -126.290 ;
        RECT 380.905 -126.325 386.230 -126.290 ;
        RECT 374.760 -127.295 377.370 -126.325 ;
        RECT 381.995 -128.350 386.230 -126.325 ;
        RECT 403.240 -125.945 414.710 -123.205 ;
        RECT 403.240 -125.980 406.285 -125.945 ;
        RECT 409.385 -125.980 414.710 -125.945 ;
        RECT 403.240 -126.950 405.850 -125.980 ;
        RECT 410.475 -128.005 414.710 -125.980 ;
        RECT 421.580 -123.360 433.210 -122.390 ;
        RECT 421.580 -126.100 433.050 -123.360 ;
        RECT 421.580 -126.135 424.625 -126.100 ;
        RECT 427.725 -126.135 433.050 -126.100 ;
        RECT 421.580 -127.105 424.190 -126.135 ;
        RECT 428.815 -128.160 433.050 -126.135 ;
        RECT 55.640 -129.665 57.345 -129.610 ;
        RECT -95.755 -130.745 -84.125 -129.775 ;
        RECT -95.625 -131.645 -84.125 -130.745 ;
        RECT -95.625 -131.680 -87.715 -131.645 ;
        RECT -95.625 -132.575 -88.150 -131.680 ;
        RECT -95.625 -132.795 -92.035 -132.575 ;
        RECT -90.760 -132.650 -88.150 -132.575 ;
        RECT 64.635 -134.580 68.840 -134.550 ;
        RECT -37.465 -135.760 -27.880 -135.395 ;
        RECT -24.965 -135.760 -15.380 -135.395 ;
        RECT -12.465 -135.760 -2.880 -135.395 ;
        RECT 0.035 -135.760 9.620 -135.395 ;
        RECT 12.535 -135.760 22.120 -135.395 ;
        RECT 27.535 -135.760 37.120 -135.395 ;
        RECT -115.005 -138.115 -107.725 -135.825 ;
        RECT -37.470 -137.770 -27.880 -135.760 ;
        RECT -24.970 -137.770 -15.380 -135.760 ;
        RECT -12.470 -137.770 -2.880 -135.760 ;
        RECT 0.030 -137.770 9.620 -135.760 ;
        RECT 12.530 -137.770 22.120 -135.760 ;
        RECT 27.530 -137.770 37.120 -135.760 ;
        RECT 57.035 -136.845 82.345 -134.580 ;
        RECT 68.665 -136.850 82.345 -136.845 ;
        RECT -114.850 -138.120 -107.725 -138.115 ;
        RECT -130.370 -207.855 -126.525 -169.855 ;
        RECT -72.445 -173.985 -58.765 -173.980 ;
        RECT -72.445 -176.250 -47.135 -173.985 ;
        RECT -58.940 -176.280 -54.735 -176.250 ;
        RECT -110.440 -177.895 -103.315 -177.890 ;
        RECT -110.440 -180.185 -103.160 -177.895 ;
        RECT -41.125 -178.300 -36.890 -173.915 ;
        RECT -33.980 -176.915 -24.390 -174.905 ;
        RECT -21.480 -176.915 -11.890 -174.905 ;
        RECT -8.980 -176.915 0.610 -174.905 ;
        RECT 3.520 -176.915 13.110 -174.905 ;
        RECT 16.020 -176.915 25.610 -174.905 ;
        RECT 31.020 -176.915 40.610 -174.905 ;
        RECT -33.975 -177.280 -24.390 -176.915 ;
        RECT -21.475 -177.280 -11.890 -176.915 ;
        RECT -8.975 -177.280 0.610 -176.915 ;
        RECT 3.525 -177.280 13.110 -176.915 ;
        RECT 16.025 -177.280 25.610 -176.915 ;
        RECT 31.025 -177.280 40.610 -176.915 ;
        RECT -100.445 -180.290 -93.810 -178.420 ;
        RECT -100.445 -180.325 -97.400 -180.290 ;
        RECT -100.445 -181.295 -97.835 -180.325 ;
        RECT -47.445 -181.220 -45.740 -181.165 ;
        RECT -92.265 -184.955 -89.655 -183.985 ;
        RECT -85.030 -184.955 -80.795 -182.930 ;
        RECT -72.510 -183.485 -42.720 -181.220 ;
        RECT -72.510 -183.490 -58.830 -183.485 ;
        RECT -31.790 -184.570 -28.690 -182.305 ;
        RECT -92.265 -184.990 -89.220 -184.955 ;
        RECT -86.120 -184.990 -80.795 -184.955 ;
        RECT -101.290 -187.575 -94.165 -187.570 ;
        RECT -110.155 -189.835 -103.520 -187.965 ;
        RECT -110.155 -189.870 -107.110 -189.835 ;
        RECT -101.290 -189.865 -94.010 -187.575 ;
        RECT -92.265 -187.730 -80.795 -184.990 ;
        RECT -92.265 -188.700 -80.635 -187.730 ;
        RECT -92.135 -189.600 -80.635 -188.700 ;
        RECT -92.135 -189.635 -84.225 -189.600 ;
        RECT -110.155 -190.840 -107.545 -189.870 ;
        RECT -92.135 -190.530 -84.660 -189.635 ;
        RECT -92.135 -190.750 -88.545 -190.530 ;
        RECT -87.270 -190.605 -84.660 -190.530 ;
        RECT -67.320 -189.835 -64.710 -188.865 ;
        RECT -60.085 -189.835 -55.850 -187.810 ;
        RECT -33.140 -188.090 40.660 -186.160 ;
        RECT 314.315 -186.370 317.905 -186.150 ;
        RECT 360.080 -186.285 363.670 -186.065 ;
        RECT 406.900 -186.095 410.490 -185.875 ;
        RECT 411.765 -186.095 414.375 -186.020 ;
        RECT 364.945 -186.285 367.555 -186.210 ;
        RECT 319.180 -186.370 321.790 -186.295 ;
        RECT 138.040 -186.620 141.630 -186.400 ;
        RECT 142.905 -186.620 145.515 -186.545 ;
        RECT 138.040 -187.515 145.515 -186.620 ;
        RECT 180.240 -186.675 183.830 -186.455 ;
        RECT 185.105 -186.675 187.715 -186.600 ;
        RECT 112.795 -187.520 126.475 -187.515 ;
        RECT -33.140 -188.440 4.990 -188.090 ;
        RECT 9.965 -188.100 40.660 -188.090 ;
        RECT 9.965 -188.125 13.010 -188.100 ;
        RECT -8.075 -188.495 -6.370 -188.440 ;
        RECT -4.940 -188.525 4.990 -188.440 ;
        RECT 10.400 -189.095 13.010 -188.125 ;
        RECT 17.990 -188.135 40.660 -188.100 ;
        RECT 18.425 -188.535 40.660 -188.135 ;
        RECT 18.425 -189.105 21.035 -188.535 ;
        RECT 101.165 -189.785 126.475 -187.520 ;
        RECT 138.040 -187.550 145.950 -187.515 ;
        RECT 138.040 -188.450 149.540 -187.550 ;
        RECT 137.910 -189.420 149.540 -188.450 ;
        RECT 180.240 -187.570 187.715 -186.675 ;
        RECT 224.555 -186.870 228.145 -186.650 ;
        RECT 270.545 -186.700 274.135 -186.480 ;
        RECT 275.410 -186.700 278.020 -186.625 ;
        RECT 229.420 -186.870 232.030 -186.795 ;
        RECT 180.240 -187.605 188.150 -187.570 ;
        RECT 180.240 -188.505 191.740 -187.605 ;
        RECT 108.765 -189.815 112.970 -189.785 ;
        RECT -67.320 -189.870 -64.275 -189.835 ;
        RECT -61.175 -189.870 -55.850 -189.835 ;
        RECT -67.320 -192.610 -55.850 -189.870 ;
        RECT -67.320 -193.580 -55.690 -192.610 ;
        RECT -19.570 -193.410 -15.365 -193.380 ;
        RECT -67.190 -194.480 -55.690 -193.580 ;
        RECT -67.190 -194.515 -59.280 -194.480 ;
        RECT -67.190 -195.410 -59.715 -194.515 ;
        RECT -67.190 -195.630 -63.600 -195.410 ;
        RECT -62.325 -195.485 -59.715 -195.410 ;
        RECT -33.075 -195.675 -7.765 -193.410 ;
        RECT 90.145 -194.755 94.870 -192.155 ;
        RECT 137.910 -192.160 149.380 -189.420 ;
        RECT 137.910 -192.195 140.955 -192.160 ;
        RECT 144.055 -192.195 149.380 -192.160 ;
        RECT 137.910 -193.165 140.520 -192.195 ;
        RECT 145.145 -194.220 149.380 -192.195 ;
        RECT 155.105 -193.010 162.490 -188.645 ;
        RECT 180.110 -189.475 191.740 -188.505 ;
        RECT 224.555 -187.765 232.030 -186.870 ;
        RECT 270.545 -187.595 278.020 -186.700 ;
        RECT 314.315 -187.265 321.790 -186.370 ;
        RECT 360.080 -187.180 367.555 -186.285 ;
        RECT 406.900 -186.990 414.375 -186.095 ;
        RECT 406.900 -187.025 414.810 -186.990 ;
        RECT 360.080 -187.215 367.990 -187.180 ;
        RECT 314.315 -187.300 322.225 -187.265 ;
        RECT 270.545 -187.630 278.455 -187.595 ;
        RECT 224.555 -187.800 232.465 -187.765 ;
        RECT 224.555 -188.700 236.055 -187.800 ;
        RECT 270.545 -188.530 282.045 -187.630 ;
        RECT 314.315 -188.200 325.815 -187.300 ;
        RECT 360.080 -188.115 371.580 -187.215 ;
        RECT 406.900 -187.925 418.400 -187.025 ;
        RECT 180.110 -192.215 191.580 -189.475 ;
        RECT 180.110 -192.250 183.155 -192.215 ;
        RECT 186.255 -192.250 191.580 -192.215 ;
        RECT 180.110 -193.220 182.720 -192.250 ;
        RECT 187.345 -194.275 191.580 -192.250 ;
        RECT 197.305 -193.065 204.690 -188.700 ;
        RECT 224.425 -189.670 236.055 -188.700 ;
        RECT 224.425 -192.410 235.895 -189.670 ;
        RECT 224.425 -192.445 227.470 -192.410 ;
        RECT 230.570 -192.445 235.895 -192.410 ;
        RECT 224.425 -193.415 227.035 -192.445 ;
        RECT 231.660 -194.470 235.895 -192.445 ;
        RECT 241.620 -193.260 249.005 -188.895 ;
        RECT 270.415 -189.500 282.045 -188.530 ;
        RECT 270.415 -192.240 281.885 -189.500 ;
        RECT 270.415 -192.275 273.460 -192.240 ;
        RECT 276.560 -192.275 281.885 -192.240 ;
        RECT 270.415 -193.245 273.025 -192.275 ;
        RECT 277.650 -194.300 281.885 -192.275 ;
        RECT 287.610 -193.090 294.995 -188.725 ;
        RECT 314.185 -189.170 325.815 -188.200 ;
        RECT 314.185 -191.910 325.655 -189.170 ;
        RECT 314.185 -191.945 317.230 -191.910 ;
        RECT 320.330 -191.945 325.655 -191.910 ;
        RECT 314.185 -192.915 316.795 -191.945 ;
        RECT 321.420 -193.970 325.655 -191.945 ;
        RECT 331.380 -192.760 338.765 -188.395 ;
        RECT 359.950 -189.085 371.580 -188.115 ;
        RECT 359.950 -191.825 371.420 -189.085 ;
        RECT 359.950 -191.860 362.995 -191.825 ;
        RECT 366.095 -191.860 371.420 -191.825 ;
        RECT 359.950 -192.830 362.560 -191.860 ;
        RECT 367.185 -193.885 371.420 -191.860 ;
        RECT 377.145 -192.675 384.530 -188.310 ;
        RECT 406.770 -188.895 418.400 -187.925 ;
        RECT 406.770 -191.635 418.240 -188.895 ;
        RECT 406.770 -191.670 409.815 -191.635 ;
        RECT 412.915 -191.670 418.240 -191.635 ;
        RECT 406.770 -192.640 409.380 -191.670 ;
        RECT 414.005 -193.695 418.240 -191.670 ;
        RECT 423.965 -192.485 431.350 -188.120 ;
        RECT 99.770 -194.755 101.475 -194.700 ;
        RECT -33.075 -195.680 -19.395 -195.675 ;
        RECT 90.140 -197.020 126.540 -194.755 ;
        RECT 108.920 -198.365 111.585 -197.020 ;
        RECT 112.860 -197.025 126.540 -197.020 ;
        RECT -72.445 -198.620 -58.765 -198.615 ;
        RECT -72.445 -200.885 -47.135 -198.620 ;
        RECT -58.940 -200.915 -54.735 -200.885 ;
        RECT -40.990 -202.970 -36.755 -198.585 ;
        RECT -33.075 -199.955 -19.395 -199.950 ;
        RECT -33.075 -202.220 -7.765 -199.955 ;
        RECT 108.975 -201.135 111.585 -198.365 ;
        RECT -19.570 -202.250 -15.365 -202.220 ;
        RECT -109.830 -208.310 -105.105 -203.585 ;
        RECT -103.800 -206.955 -100.625 -203.550 ;
        RECT -99.275 -206.960 -96.100 -203.555 ;
        RECT -47.445 -205.855 -45.740 -205.800 ;
        RECT -92.265 -209.955 -89.655 -208.985 ;
        RECT -85.030 -209.955 -80.795 -207.930 ;
        RECT -72.510 -208.120 -42.720 -205.855 ;
        RECT -8.075 -207.190 -6.370 -207.135 ;
        RECT -4.940 -207.190 4.990 -207.105 ;
        RECT -33.140 -207.540 4.990 -207.190 ;
        RECT 10.400 -207.505 13.010 -206.535 ;
        RECT 18.425 -207.095 21.035 -206.525 ;
        RECT 18.425 -207.495 40.660 -207.095 ;
        RECT 9.965 -207.530 13.010 -207.505 ;
        RECT 17.990 -207.530 40.660 -207.495 ;
        RECT 9.965 -207.540 40.660 -207.530 ;
        RECT -72.510 -208.125 -58.830 -208.120 ;
        RECT -33.140 -209.470 40.660 -207.540 ;
        RECT 90.120 -208.290 93.295 -204.885 ;
        RECT 94.850 -208.290 98.025 -204.885 ;
        RECT 99.430 -208.345 106.710 -206.055 ;
        RECT 108.725 -208.285 111.825 -206.020 ;
        RECT 113.125 -208.325 126.755 -203.165 ;
        RECT 314.275 -203.635 317.865 -203.415 ;
        RECT 360.040 -203.550 363.630 -203.330 ;
        RECT 406.860 -203.360 410.450 -203.140 ;
        RECT 411.725 -203.360 414.335 -203.285 ;
        RECT 364.905 -203.550 367.515 -203.475 ;
        RECT 319.140 -203.635 321.750 -203.560 ;
        RECT 138.000 -203.885 141.590 -203.665 ;
        RECT 142.865 -203.885 145.475 -203.810 ;
        RECT 138.000 -204.780 145.475 -203.885 ;
        RECT 156.340 -204.040 159.930 -203.820 ;
        RECT 180.200 -203.940 183.790 -203.720 ;
        RECT 185.065 -203.940 187.675 -203.865 ;
        RECT 161.205 -204.040 163.815 -203.965 ;
        RECT 138.000 -204.815 145.910 -204.780 ;
        RECT 138.000 -205.715 149.500 -204.815 ;
        RECT 137.870 -206.685 149.500 -205.715 ;
        RECT 156.340 -204.935 163.815 -204.040 ;
        RECT 180.200 -204.835 187.675 -203.940 ;
        RECT 198.540 -204.095 202.130 -203.875 ;
        RECT 203.405 -204.095 206.015 -204.020 ;
        RECT 180.200 -204.870 188.110 -204.835 ;
        RECT 156.340 -204.970 164.250 -204.935 ;
        RECT 156.340 -205.870 167.840 -204.970 ;
        RECT 180.200 -205.770 191.700 -204.870 ;
        RECT 99.430 -208.350 106.555 -208.345 ;
        RECT 137.870 -209.425 149.340 -206.685 ;
        RECT 137.870 -209.460 140.915 -209.425 ;
        RECT 144.015 -209.460 149.340 -209.425 ;
        RECT -92.265 -209.990 -89.220 -209.955 ;
        RECT -86.120 -209.990 -80.795 -209.955 ;
        RECT -92.265 -212.730 -80.795 -209.990 ;
        RECT 72.220 -210.300 85.900 -210.295 ;
        RECT 56.110 -212.565 85.900 -210.300 ;
        RECT 137.870 -210.430 140.480 -209.460 ;
        RECT 145.105 -211.485 149.340 -209.460 ;
        RECT 156.210 -206.840 167.840 -205.870 ;
        RECT 180.070 -206.740 191.700 -205.770 ;
        RECT 198.540 -204.990 206.015 -204.095 ;
        RECT 224.515 -204.135 228.105 -203.915 ;
        RECT 270.505 -203.965 274.095 -203.745 ;
        RECT 275.370 -203.965 277.980 -203.890 ;
        RECT 229.380 -204.135 231.990 -204.060 ;
        RECT 198.540 -205.025 206.450 -204.990 ;
        RECT 198.540 -205.925 210.040 -205.025 ;
        RECT 156.210 -209.580 167.680 -206.840 ;
        RECT 156.210 -209.615 159.255 -209.580 ;
        RECT 162.355 -209.615 167.680 -209.580 ;
        RECT 156.210 -210.585 158.820 -209.615 ;
        RECT 163.445 -211.640 167.680 -209.615 ;
        RECT 180.070 -209.480 191.540 -206.740 ;
        RECT 180.070 -209.515 183.115 -209.480 ;
        RECT 186.215 -209.515 191.540 -209.480 ;
        RECT 180.070 -210.485 182.680 -209.515 ;
        RECT 187.305 -211.540 191.540 -209.515 ;
        RECT 198.410 -206.895 210.040 -205.925 ;
        RECT 224.515 -205.030 231.990 -204.135 ;
        RECT 242.855 -204.290 246.445 -204.070 ;
        RECT 247.720 -204.290 250.330 -204.215 ;
        RECT 224.515 -205.065 232.425 -205.030 ;
        RECT 224.515 -205.965 236.015 -205.065 ;
        RECT 198.410 -209.635 209.880 -206.895 ;
        RECT 198.410 -209.670 201.455 -209.635 ;
        RECT 204.555 -209.670 209.880 -209.635 ;
        RECT 198.410 -210.640 201.020 -209.670 ;
        RECT 205.645 -211.695 209.880 -209.670 ;
        RECT 224.385 -206.935 236.015 -205.965 ;
        RECT 242.855 -205.185 250.330 -204.290 ;
        RECT 270.505 -204.860 277.980 -203.965 ;
        RECT 288.845 -204.120 292.435 -203.900 ;
        RECT 293.710 -204.120 296.320 -204.045 ;
        RECT 270.505 -204.895 278.415 -204.860 ;
        RECT 242.855 -205.220 250.765 -205.185 ;
        RECT 242.855 -206.120 254.355 -205.220 ;
        RECT 270.505 -205.795 282.005 -204.895 ;
        RECT 224.385 -209.675 235.855 -206.935 ;
        RECT 224.385 -209.710 227.430 -209.675 ;
        RECT 230.530 -209.710 235.855 -209.675 ;
        RECT 224.385 -210.680 226.995 -209.710 ;
        RECT 231.620 -211.735 235.855 -209.710 ;
        RECT 242.725 -207.090 254.355 -206.120 ;
        RECT 270.375 -206.765 282.005 -205.795 ;
        RECT 288.845 -205.015 296.320 -204.120 ;
        RECT 314.275 -204.530 321.750 -203.635 ;
        RECT 332.615 -203.790 336.205 -203.570 ;
        RECT 337.480 -203.790 340.090 -203.715 ;
        RECT 314.275 -204.565 322.185 -204.530 ;
        RECT 288.845 -205.050 296.755 -205.015 ;
        RECT 288.845 -205.950 300.345 -205.050 ;
        RECT 314.275 -205.465 325.775 -204.565 ;
        RECT 242.725 -209.830 254.195 -207.090 ;
        RECT 242.725 -209.865 245.770 -209.830 ;
        RECT 248.870 -209.865 254.195 -209.830 ;
        RECT 242.725 -210.835 245.335 -209.865 ;
        RECT 249.960 -211.890 254.195 -209.865 ;
        RECT 270.375 -209.505 281.845 -206.765 ;
        RECT 270.375 -209.540 273.420 -209.505 ;
        RECT 276.520 -209.540 281.845 -209.505 ;
        RECT 270.375 -210.510 272.985 -209.540 ;
        RECT 277.610 -211.565 281.845 -209.540 ;
        RECT 288.715 -206.920 300.345 -205.950 ;
        RECT 314.145 -206.435 325.775 -205.465 ;
        RECT 332.615 -204.685 340.090 -203.790 ;
        RECT 360.040 -204.445 367.515 -203.550 ;
        RECT 378.380 -203.705 381.970 -203.485 ;
        RECT 383.245 -203.705 385.855 -203.630 ;
        RECT 360.040 -204.480 367.950 -204.445 ;
        RECT 332.615 -204.720 340.525 -204.685 ;
        RECT 332.615 -205.620 344.115 -204.720 ;
        RECT 360.040 -205.380 371.540 -204.480 ;
        RECT 288.715 -209.660 300.185 -206.920 ;
        RECT 288.715 -209.695 291.760 -209.660 ;
        RECT 294.860 -209.695 300.185 -209.660 ;
        RECT 288.715 -210.665 291.325 -209.695 ;
        RECT 295.950 -211.720 300.185 -209.695 ;
        RECT 314.145 -209.175 325.615 -206.435 ;
        RECT 314.145 -209.210 317.190 -209.175 ;
        RECT 320.290 -209.210 325.615 -209.175 ;
        RECT 314.145 -210.180 316.755 -209.210 ;
        RECT 321.380 -211.235 325.615 -209.210 ;
        RECT 332.485 -206.590 344.115 -205.620 ;
        RECT 359.910 -206.350 371.540 -205.380 ;
        RECT 378.380 -204.600 385.855 -203.705 ;
        RECT 406.860 -204.255 414.335 -203.360 ;
        RECT 425.200 -203.515 428.790 -203.295 ;
        RECT 430.065 -203.515 432.675 -203.440 ;
        RECT 406.860 -204.290 414.770 -204.255 ;
        RECT 378.380 -204.635 386.290 -204.600 ;
        RECT 378.380 -205.535 389.880 -204.635 ;
        RECT 406.860 -205.190 418.360 -204.290 ;
        RECT 332.485 -209.330 343.955 -206.590 ;
        RECT 332.485 -209.365 335.530 -209.330 ;
        RECT 338.630 -209.365 343.955 -209.330 ;
        RECT 332.485 -210.335 335.095 -209.365 ;
        RECT 339.720 -211.390 343.955 -209.365 ;
        RECT 359.910 -209.090 371.380 -206.350 ;
        RECT 359.910 -209.125 362.955 -209.090 ;
        RECT 366.055 -209.125 371.380 -209.090 ;
        RECT 359.910 -210.095 362.520 -209.125 ;
        RECT 367.145 -211.150 371.380 -209.125 ;
        RECT 378.250 -206.505 389.880 -205.535 ;
        RECT 406.730 -206.160 418.360 -205.190 ;
        RECT 425.200 -204.410 432.675 -203.515 ;
        RECT 425.200 -204.445 433.110 -204.410 ;
        RECT 425.200 -205.345 436.700 -204.445 ;
        RECT 378.250 -209.245 389.720 -206.505 ;
        RECT 378.250 -209.280 381.295 -209.245 ;
        RECT 384.395 -209.280 389.720 -209.245 ;
        RECT 378.250 -210.250 380.860 -209.280 ;
        RECT 385.485 -211.305 389.720 -209.280 ;
        RECT 406.730 -208.900 418.200 -206.160 ;
        RECT 406.730 -208.935 409.775 -208.900 ;
        RECT 412.875 -208.935 418.200 -208.900 ;
        RECT 406.730 -209.905 409.340 -208.935 ;
        RECT 413.965 -210.960 418.200 -208.935 ;
        RECT 425.070 -206.315 436.700 -205.345 ;
        RECT 425.070 -209.055 436.540 -206.315 ;
        RECT 425.070 -209.090 428.115 -209.055 ;
        RECT 431.215 -209.090 436.540 -209.055 ;
        RECT 425.070 -210.060 427.680 -209.090 ;
        RECT 432.305 -211.115 436.540 -209.090 ;
        RECT 59.130 -212.620 60.835 -212.565 ;
        RECT -92.265 -213.700 -80.635 -212.730 ;
        RECT -92.135 -214.600 -80.635 -213.700 ;
        RECT -92.135 -214.635 -84.225 -214.600 ;
        RECT -92.135 -215.530 -84.660 -214.635 ;
        RECT -92.135 -215.750 -88.545 -215.530 ;
        RECT -87.270 -215.605 -84.660 -215.530 ;
        RECT 68.125 -217.535 72.330 -217.505 ;
        RECT -33.975 -218.715 -24.390 -218.350 ;
        RECT -21.475 -218.715 -11.890 -218.350 ;
        RECT -8.975 -218.715 0.610 -218.350 ;
        RECT 3.525 -218.715 13.110 -218.350 ;
        RECT 16.025 -218.715 25.610 -218.350 ;
        RECT 31.025 -218.715 40.610 -218.350 ;
        RECT -111.515 -221.070 -104.235 -218.780 ;
        RECT -33.980 -220.725 -24.390 -218.715 ;
        RECT -21.480 -220.725 -11.890 -218.715 ;
        RECT -8.980 -220.725 0.610 -218.715 ;
        RECT 3.520 -220.725 13.110 -218.715 ;
        RECT 16.020 -220.725 25.610 -218.715 ;
        RECT 31.020 -220.725 40.610 -218.715 ;
        RECT 60.525 -219.800 85.835 -217.535 ;
        RECT 72.155 -219.805 85.835 -219.800 ;
        RECT -111.360 -221.075 -104.235 -221.070 ;
        RECT -139.470 -298.580 -135.625 -260.580 ;
        RECT -68.930 -264.540 -55.250 -264.535 ;
        RECT -68.930 -266.805 -43.620 -264.540 ;
        RECT -55.425 -266.835 -51.220 -266.805 ;
        RECT -106.925 -268.450 -99.800 -268.445 ;
        RECT -106.925 -270.740 -99.645 -268.450 ;
        RECT -37.610 -268.855 -33.375 -264.470 ;
        RECT -30.465 -267.470 -20.875 -265.460 ;
        RECT -17.965 -267.470 -8.375 -265.460 ;
        RECT -5.465 -267.470 4.125 -265.460 ;
        RECT 7.035 -267.470 16.625 -265.460 ;
        RECT 19.535 -267.470 29.125 -265.460 ;
        RECT 34.535 -267.470 44.125 -265.460 ;
        RECT -30.460 -267.835 -20.875 -267.470 ;
        RECT -17.960 -267.835 -8.375 -267.470 ;
        RECT -5.460 -267.835 4.125 -267.470 ;
        RECT 7.040 -267.835 16.625 -267.470 ;
        RECT 19.540 -267.835 29.125 -267.470 ;
        RECT 34.540 -267.835 44.125 -267.470 ;
        RECT -96.930 -270.845 -90.295 -268.975 ;
        RECT -96.930 -270.880 -93.885 -270.845 ;
        RECT -96.930 -271.850 -94.320 -270.880 ;
        RECT -43.930 -271.775 -42.225 -271.720 ;
        RECT -88.750 -275.510 -86.140 -274.540 ;
        RECT -81.515 -275.510 -77.280 -273.485 ;
        RECT -68.995 -274.040 -39.205 -271.775 ;
        RECT -68.995 -274.045 -55.315 -274.040 ;
        RECT -28.275 -275.125 -25.175 -272.860 ;
        RECT -88.750 -275.545 -85.705 -275.510 ;
        RECT -82.605 -275.545 -77.280 -275.510 ;
        RECT -97.775 -278.130 -90.650 -278.125 ;
        RECT -106.640 -280.390 -100.005 -278.520 ;
        RECT -106.640 -280.425 -103.595 -280.390 ;
        RECT -97.775 -280.420 -90.495 -278.130 ;
        RECT -88.750 -278.285 -77.280 -275.545 ;
        RECT -88.750 -279.255 -77.120 -278.285 ;
        RECT -88.620 -280.155 -77.120 -279.255 ;
        RECT -88.620 -280.190 -80.710 -280.155 ;
        RECT -106.640 -281.395 -104.030 -280.425 ;
        RECT -88.620 -281.085 -81.145 -280.190 ;
        RECT -88.620 -281.305 -85.030 -281.085 ;
        RECT -83.755 -281.160 -81.145 -281.085 ;
        RECT -63.805 -280.390 -61.195 -279.420 ;
        RECT -56.570 -280.390 -52.335 -278.365 ;
        RECT -29.625 -278.645 44.175 -276.715 ;
        RECT 317.830 -276.925 321.420 -276.705 ;
        RECT 363.595 -276.840 367.185 -276.620 ;
        RECT 410.415 -276.650 414.005 -276.430 ;
        RECT 415.280 -276.650 417.890 -276.575 ;
        RECT 368.460 -276.840 371.070 -276.765 ;
        RECT 322.695 -276.925 325.305 -276.850 ;
        RECT 141.555 -277.175 145.145 -276.955 ;
        RECT 146.420 -277.175 149.030 -277.100 ;
        RECT 141.555 -278.070 149.030 -277.175 ;
        RECT 183.755 -277.230 187.345 -277.010 ;
        RECT 188.620 -277.230 191.230 -277.155 ;
        RECT 116.310 -278.075 129.990 -278.070 ;
        RECT -29.625 -278.995 8.505 -278.645 ;
        RECT 13.480 -278.655 44.175 -278.645 ;
        RECT 13.480 -278.680 16.525 -278.655 ;
        RECT -4.560 -279.050 -2.855 -278.995 ;
        RECT -1.425 -279.080 8.505 -278.995 ;
        RECT 13.915 -279.650 16.525 -278.680 ;
        RECT 21.505 -278.690 44.175 -278.655 ;
        RECT 21.940 -279.090 44.175 -278.690 ;
        RECT 21.940 -279.660 24.550 -279.090 ;
        RECT 104.680 -280.340 129.990 -278.075 ;
        RECT 141.555 -278.105 149.465 -278.070 ;
        RECT 141.555 -279.005 153.055 -278.105 ;
        RECT 141.425 -279.975 153.055 -279.005 ;
        RECT 183.755 -278.125 191.230 -277.230 ;
        RECT 228.070 -277.425 231.660 -277.205 ;
        RECT 274.060 -277.255 277.650 -277.035 ;
        RECT 278.925 -277.255 281.535 -277.180 ;
        RECT 232.935 -277.425 235.545 -277.350 ;
        RECT 183.755 -278.160 191.665 -278.125 ;
        RECT 183.755 -279.060 195.255 -278.160 ;
        RECT 112.280 -280.370 116.485 -280.340 ;
        RECT -63.805 -280.425 -60.760 -280.390 ;
        RECT -57.660 -280.425 -52.335 -280.390 ;
        RECT -63.805 -283.165 -52.335 -280.425 ;
        RECT -63.805 -284.135 -52.175 -283.165 ;
        RECT -16.055 -283.965 -11.850 -283.935 ;
        RECT -63.675 -285.035 -52.175 -284.135 ;
        RECT -63.675 -285.070 -55.765 -285.035 ;
        RECT -63.675 -285.965 -56.200 -285.070 ;
        RECT -63.675 -286.185 -60.085 -285.965 ;
        RECT -58.810 -286.040 -56.200 -285.965 ;
        RECT -29.560 -286.230 -4.250 -283.965 ;
        RECT 93.660 -285.310 98.385 -282.710 ;
        RECT 141.425 -282.715 152.895 -279.975 ;
        RECT 141.425 -282.750 144.470 -282.715 ;
        RECT 147.570 -282.750 152.895 -282.715 ;
        RECT 141.425 -283.720 144.035 -282.750 ;
        RECT 148.660 -284.775 152.895 -282.750 ;
        RECT 158.620 -283.565 166.005 -279.200 ;
        RECT 183.625 -280.030 195.255 -279.060 ;
        RECT 228.070 -278.320 235.545 -277.425 ;
        RECT 274.060 -278.150 281.535 -277.255 ;
        RECT 317.830 -277.820 325.305 -276.925 ;
        RECT 363.595 -277.735 371.070 -276.840 ;
        RECT 410.415 -277.545 417.890 -276.650 ;
        RECT 410.415 -277.580 418.325 -277.545 ;
        RECT 363.595 -277.770 371.505 -277.735 ;
        RECT 317.830 -277.855 325.740 -277.820 ;
        RECT 274.060 -278.185 281.970 -278.150 ;
        RECT 228.070 -278.355 235.980 -278.320 ;
        RECT 228.070 -279.255 239.570 -278.355 ;
        RECT 274.060 -279.085 285.560 -278.185 ;
        RECT 317.830 -278.755 329.330 -277.855 ;
        RECT 363.595 -278.670 375.095 -277.770 ;
        RECT 410.415 -278.480 421.915 -277.580 ;
        RECT 183.625 -282.770 195.095 -280.030 ;
        RECT 183.625 -282.805 186.670 -282.770 ;
        RECT 189.770 -282.805 195.095 -282.770 ;
        RECT 183.625 -283.775 186.235 -282.805 ;
        RECT 190.860 -284.830 195.095 -282.805 ;
        RECT 200.820 -283.620 208.205 -279.255 ;
        RECT 227.940 -280.225 239.570 -279.255 ;
        RECT 227.940 -282.965 239.410 -280.225 ;
        RECT 227.940 -283.000 230.985 -282.965 ;
        RECT 234.085 -283.000 239.410 -282.965 ;
        RECT 227.940 -283.970 230.550 -283.000 ;
        RECT 235.175 -285.025 239.410 -283.000 ;
        RECT 245.135 -283.815 252.520 -279.450 ;
        RECT 273.930 -280.055 285.560 -279.085 ;
        RECT 273.930 -282.795 285.400 -280.055 ;
        RECT 273.930 -282.830 276.975 -282.795 ;
        RECT 280.075 -282.830 285.400 -282.795 ;
        RECT 273.930 -283.800 276.540 -282.830 ;
        RECT 281.165 -284.855 285.400 -282.830 ;
        RECT 291.125 -283.645 298.510 -279.280 ;
        RECT 317.700 -279.725 329.330 -278.755 ;
        RECT 317.700 -282.465 329.170 -279.725 ;
        RECT 317.700 -282.500 320.745 -282.465 ;
        RECT 323.845 -282.500 329.170 -282.465 ;
        RECT 317.700 -283.470 320.310 -282.500 ;
        RECT 324.935 -284.525 329.170 -282.500 ;
        RECT 334.895 -283.315 342.280 -278.950 ;
        RECT 363.465 -279.640 375.095 -278.670 ;
        RECT 363.465 -282.380 374.935 -279.640 ;
        RECT 363.465 -282.415 366.510 -282.380 ;
        RECT 369.610 -282.415 374.935 -282.380 ;
        RECT 363.465 -283.385 366.075 -282.415 ;
        RECT 370.700 -284.440 374.935 -282.415 ;
        RECT 380.660 -283.230 388.045 -278.865 ;
        RECT 410.285 -279.450 421.915 -278.480 ;
        RECT 410.285 -282.190 421.755 -279.450 ;
        RECT 410.285 -282.225 413.330 -282.190 ;
        RECT 416.430 -282.225 421.755 -282.190 ;
        RECT 410.285 -283.195 412.895 -282.225 ;
        RECT 417.520 -284.250 421.755 -282.225 ;
        RECT 427.480 -283.040 434.865 -278.675 ;
        RECT 103.285 -285.310 104.990 -285.255 ;
        RECT -29.560 -286.235 -15.880 -286.230 ;
        RECT 93.655 -287.575 130.055 -285.310 ;
        RECT 112.435 -288.920 115.100 -287.575 ;
        RECT 116.375 -287.580 130.055 -287.575 ;
        RECT -68.930 -289.175 -55.250 -289.170 ;
        RECT -68.930 -291.440 -43.620 -289.175 ;
        RECT -55.425 -291.470 -51.220 -291.440 ;
        RECT -37.475 -293.525 -33.240 -289.140 ;
        RECT -29.560 -290.510 -15.880 -290.505 ;
        RECT -29.560 -292.775 -4.250 -290.510 ;
        RECT 112.490 -291.690 115.100 -288.920 ;
        RECT -16.055 -292.805 -11.850 -292.775 ;
        RECT -106.315 -298.865 -101.590 -294.140 ;
        RECT -100.285 -297.510 -97.110 -294.105 ;
        RECT -95.760 -297.515 -92.585 -294.110 ;
        RECT -43.930 -296.410 -42.225 -296.355 ;
        RECT -88.750 -300.510 -86.140 -299.540 ;
        RECT -81.515 -300.510 -77.280 -298.485 ;
        RECT -68.995 -298.675 -39.205 -296.410 ;
        RECT -4.560 -297.745 -2.855 -297.690 ;
        RECT -1.425 -297.745 8.505 -297.660 ;
        RECT -29.625 -298.095 8.505 -297.745 ;
        RECT 13.915 -298.060 16.525 -297.090 ;
        RECT 21.940 -297.650 24.550 -297.080 ;
        RECT 21.940 -298.050 44.175 -297.650 ;
        RECT 13.480 -298.085 16.525 -298.060 ;
        RECT 21.505 -298.085 44.175 -298.050 ;
        RECT 13.480 -298.095 44.175 -298.085 ;
        RECT -68.995 -298.680 -55.315 -298.675 ;
        RECT -29.625 -300.025 44.175 -298.095 ;
        RECT 93.635 -298.845 96.810 -295.440 ;
        RECT 98.365 -298.845 101.540 -295.440 ;
        RECT 102.945 -298.900 110.225 -296.610 ;
        RECT 112.240 -298.840 115.340 -296.575 ;
        RECT 116.640 -298.880 130.270 -293.720 ;
        RECT 317.790 -294.190 321.380 -293.970 ;
        RECT 363.555 -294.105 367.145 -293.885 ;
        RECT 410.375 -293.915 413.965 -293.695 ;
        RECT 415.240 -293.915 417.850 -293.840 ;
        RECT 368.420 -294.105 371.030 -294.030 ;
        RECT 322.655 -294.190 325.265 -294.115 ;
        RECT 141.515 -294.440 145.105 -294.220 ;
        RECT 146.380 -294.440 148.990 -294.365 ;
        RECT 141.515 -295.335 148.990 -294.440 ;
        RECT 159.855 -294.595 163.445 -294.375 ;
        RECT 183.715 -294.495 187.305 -294.275 ;
        RECT 188.580 -294.495 191.190 -294.420 ;
        RECT 164.720 -294.595 167.330 -294.520 ;
        RECT 141.515 -295.370 149.425 -295.335 ;
        RECT 141.515 -296.270 153.015 -295.370 ;
        RECT 141.385 -297.240 153.015 -296.270 ;
        RECT 159.855 -295.490 167.330 -294.595 ;
        RECT 183.715 -295.390 191.190 -294.495 ;
        RECT 202.055 -294.650 205.645 -294.430 ;
        RECT 206.920 -294.650 209.530 -294.575 ;
        RECT 183.715 -295.425 191.625 -295.390 ;
        RECT 159.855 -295.525 167.765 -295.490 ;
        RECT 159.855 -296.425 171.355 -295.525 ;
        RECT 183.715 -296.325 195.215 -295.425 ;
        RECT 102.945 -298.905 110.070 -298.900 ;
        RECT 141.385 -299.980 152.855 -297.240 ;
        RECT 141.385 -300.015 144.430 -299.980 ;
        RECT 147.530 -300.015 152.855 -299.980 ;
        RECT -88.750 -300.545 -85.705 -300.510 ;
        RECT -82.605 -300.545 -77.280 -300.510 ;
        RECT -88.750 -303.285 -77.280 -300.545 ;
        RECT 75.735 -300.855 89.415 -300.850 ;
        RECT 59.625 -303.120 89.415 -300.855 ;
        RECT 141.385 -300.985 143.995 -300.015 ;
        RECT 148.620 -302.040 152.855 -300.015 ;
        RECT 159.725 -297.395 171.355 -296.425 ;
        RECT 183.585 -297.295 195.215 -296.325 ;
        RECT 202.055 -295.545 209.530 -294.650 ;
        RECT 228.030 -294.690 231.620 -294.470 ;
        RECT 274.020 -294.520 277.610 -294.300 ;
        RECT 278.885 -294.520 281.495 -294.445 ;
        RECT 232.895 -294.690 235.505 -294.615 ;
        RECT 202.055 -295.580 209.965 -295.545 ;
        RECT 202.055 -296.480 213.555 -295.580 ;
        RECT 159.725 -300.135 171.195 -297.395 ;
        RECT 159.725 -300.170 162.770 -300.135 ;
        RECT 165.870 -300.170 171.195 -300.135 ;
        RECT 159.725 -301.140 162.335 -300.170 ;
        RECT 166.960 -302.195 171.195 -300.170 ;
        RECT 183.585 -300.035 195.055 -297.295 ;
        RECT 183.585 -300.070 186.630 -300.035 ;
        RECT 189.730 -300.070 195.055 -300.035 ;
        RECT 183.585 -301.040 186.195 -300.070 ;
        RECT 190.820 -302.095 195.055 -300.070 ;
        RECT 201.925 -297.450 213.555 -296.480 ;
        RECT 228.030 -295.585 235.505 -294.690 ;
        RECT 246.370 -294.845 249.960 -294.625 ;
        RECT 251.235 -294.845 253.845 -294.770 ;
        RECT 228.030 -295.620 235.940 -295.585 ;
        RECT 228.030 -296.520 239.530 -295.620 ;
        RECT 201.925 -300.190 213.395 -297.450 ;
        RECT 201.925 -300.225 204.970 -300.190 ;
        RECT 208.070 -300.225 213.395 -300.190 ;
        RECT 201.925 -301.195 204.535 -300.225 ;
        RECT 209.160 -302.250 213.395 -300.225 ;
        RECT 227.900 -297.490 239.530 -296.520 ;
        RECT 246.370 -295.740 253.845 -294.845 ;
        RECT 274.020 -295.415 281.495 -294.520 ;
        RECT 292.360 -294.675 295.950 -294.455 ;
        RECT 297.225 -294.675 299.835 -294.600 ;
        RECT 274.020 -295.450 281.930 -295.415 ;
        RECT 246.370 -295.775 254.280 -295.740 ;
        RECT 246.370 -296.675 257.870 -295.775 ;
        RECT 274.020 -296.350 285.520 -295.450 ;
        RECT 227.900 -300.230 239.370 -297.490 ;
        RECT 227.900 -300.265 230.945 -300.230 ;
        RECT 234.045 -300.265 239.370 -300.230 ;
        RECT 227.900 -301.235 230.510 -300.265 ;
        RECT 235.135 -302.290 239.370 -300.265 ;
        RECT 246.240 -297.645 257.870 -296.675 ;
        RECT 273.890 -297.320 285.520 -296.350 ;
        RECT 292.360 -295.570 299.835 -294.675 ;
        RECT 317.790 -295.085 325.265 -294.190 ;
        RECT 336.130 -294.345 339.720 -294.125 ;
        RECT 340.995 -294.345 343.605 -294.270 ;
        RECT 317.790 -295.120 325.700 -295.085 ;
        RECT 292.360 -295.605 300.270 -295.570 ;
        RECT 292.360 -296.505 303.860 -295.605 ;
        RECT 317.790 -296.020 329.290 -295.120 ;
        RECT 246.240 -300.385 257.710 -297.645 ;
        RECT 246.240 -300.420 249.285 -300.385 ;
        RECT 252.385 -300.420 257.710 -300.385 ;
        RECT 246.240 -301.390 248.850 -300.420 ;
        RECT 253.475 -302.445 257.710 -300.420 ;
        RECT 273.890 -300.060 285.360 -297.320 ;
        RECT 273.890 -300.095 276.935 -300.060 ;
        RECT 280.035 -300.095 285.360 -300.060 ;
        RECT 273.890 -301.065 276.500 -300.095 ;
        RECT 281.125 -302.120 285.360 -300.095 ;
        RECT 292.230 -297.475 303.860 -296.505 ;
        RECT 317.660 -296.990 329.290 -296.020 ;
        RECT 336.130 -295.240 343.605 -294.345 ;
        RECT 363.555 -295.000 371.030 -294.105 ;
        RECT 381.895 -294.260 385.485 -294.040 ;
        RECT 386.760 -294.260 389.370 -294.185 ;
        RECT 363.555 -295.035 371.465 -295.000 ;
        RECT 336.130 -295.275 344.040 -295.240 ;
        RECT 336.130 -296.175 347.630 -295.275 ;
        RECT 363.555 -295.935 375.055 -295.035 ;
        RECT 292.230 -300.215 303.700 -297.475 ;
        RECT 292.230 -300.250 295.275 -300.215 ;
        RECT 298.375 -300.250 303.700 -300.215 ;
        RECT 292.230 -301.220 294.840 -300.250 ;
        RECT 299.465 -302.275 303.700 -300.250 ;
        RECT 317.660 -299.730 329.130 -296.990 ;
        RECT 317.660 -299.765 320.705 -299.730 ;
        RECT 323.805 -299.765 329.130 -299.730 ;
        RECT 317.660 -300.735 320.270 -299.765 ;
        RECT 324.895 -301.790 329.130 -299.765 ;
        RECT 336.000 -297.145 347.630 -296.175 ;
        RECT 363.425 -296.905 375.055 -295.935 ;
        RECT 381.895 -295.155 389.370 -294.260 ;
        RECT 410.375 -294.810 417.850 -293.915 ;
        RECT 428.715 -294.070 432.305 -293.850 ;
        RECT 433.580 -294.070 436.190 -293.995 ;
        RECT 410.375 -294.845 418.285 -294.810 ;
        RECT 381.895 -295.190 389.805 -295.155 ;
        RECT 381.895 -296.090 393.395 -295.190 ;
        RECT 410.375 -295.745 421.875 -294.845 ;
        RECT 336.000 -299.885 347.470 -297.145 ;
        RECT 336.000 -299.920 339.045 -299.885 ;
        RECT 342.145 -299.920 347.470 -299.885 ;
        RECT 336.000 -300.890 338.610 -299.920 ;
        RECT 343.235 -301.945 347.470 -299.920 ;
        RECT 363.425 -299.645 374.895 -296.905 ;
        RECT 363.425 -299.680 366.470 -299.645 ;
        RECT 369.570 -299.680 374.895 -299.645 ;
        RECT 363.425 -300.650 366.035 -299.680 ;
        RECT 370.660 -301.705 374.895 -299.680 ;
        RECT 381.765 -297.060 393.395 -296.090 ;
        RECT 410.245 -296.715 421.875 -295.745 ;
        RECT 428.715 -294.965 436.190 -294.070 ;
        RECT 428.715 -295.000 436.625 -294.965 ;
        RECT 428.715 -295.900 440.215 -295.000 ;
        RECT 381.765 -299.800 393.235 -297.060 ;
        RECT 381.765 -299.835 384.810 -299.800 ;
        RECT 387.910 -299.835 393.235 -299.800 ;
        RECT 381.765 -300.805 384.375 -299.835 ;
        RECT 389.000 -301.860 393.235 -299.835 ;
        RECT 410.245 -299.455 421.715 -296.715 ;
        RECT 410.245 -299.490 413.290 -299.455 ;
        RECT 416.390 -299.490 421.715 -299.455 ;
        RECT 410.245 -300.460 412.855 -299.490 ;
        RECT 417.480 -301.515 421.715 -299.490 ;
        RECT 428.585 -296.870 440.215 -295.900 ;
        RECT 428.585 -299.610 440.055 -296.870 ;
        RECT 428.585 -299.645 431.630 -299.610 ;
        RECT 434.730 -299.645 440.055 -299.610 ;
        RECT 428.585 -300.615 431.195 -299.645 ;
        RECT 435.820 -301.670 440.055 -299.645 ;
        RECT 62.645 -303.175 64.350 -303.120 ;
        RECT -88.750 -304.255 -77.120 -303.285 ;
        RECT -88.620 -305.155 -77.120 -304.255 ;
        RECT -88.620 -305.190 -80.710 -305.155 ;
        RECT -88.620 -306.085 -81.145 -305.190 ;
        RECT -88.620 -306.305 -85.030 -306.085 ;
        RECT -83.755 -306.160 -81.145 -306.085 ;
        RECT 71.640 -308.090 75.845 -308.060 ;
        RECT -30.460 -309.270 -20.875 -308.905 ;
        RECT -17.960 -309.270 -8.375 -308.905 ;
        RECT -5.460 -309.270 4.125 -308.905 ;
        RECT 7.040 -309.270 16.625 -308.905 ;
        RECT 19.540 -309.270 29.125 -308.905 ;
        RECT 34.540 -309.270 44.125 -308.905 ;
        RECT -108.000 -311.625 -100.720 -309.335 ;
        RECT -30.465 -311.280 -20.875 -309.270 ;
        RECT -17.965 -311.280 -8.375 -309.270 ;
        RECT -5.465 -311.280 4.125 -309.270 ;
        RECT 7.035 -311.280 16.625 -309.270 ;
        RECT 19.535 -311.280 29.125 -309.270 ;
        RECT 34.535 -311.280 44.125 -309.270 ;
        RECT 64.040 -310.355 89.350 -308.090 ;
        RECT 75.670 -310.360 89.350 -310.355 ;
        RECT -107.845 -311.630 -100.720 -311.625 ;
      LAYER li1 ;
        RECT -56.590 601.610 -50.305 601.975 ;
        RECT -56.730 601.365 -50.305 601.610 ;
        RECT -56.730 600.915 -55.895 601.365 ;
        RECT -56.665 599.665 -55.970 600.060 ;
        RECT -56.540 599.410 -56.125 599.665 ;
        RECT -56.635 599.165 -56.125 599.410 ;
        RECT -55.450 599.535 -54.955 599.775 ;
        RECT -55.450 599.365 -54.125 599.535 ;
        RECT -50.915 599.425 -50.305 601.365 ;
        RECT -56.635 598.905 -56.305 599.165 ;
        RECT -57.255 598.890 -56.305 598.905 ;
        RECT -57.255 598.885 -55.750 598.890 ;
        RECT -60.215 598.715 -55.750 598.885 ;
        RECT -57.255 598.680 -55.750 598.715 ;
        RECT -56.635 596.795 -55.750 598.680 ;
        RECT -57.250 596.770 -55.750 596.795 ;
        RECT -60.215 596.600 -55.750 596.770 ;
        RECT -57.250 596.570 -55.750 596.600 ;
        RECT -56.635 596.415 -55.750 596.570 ;
        RECT -55.450 598.555 -54.955 599.365 ;
        RECT -50.915 598.815 -37.710 599.425 ;
        RECT -55.450 598.385 -54.125 598.555 ;
        RECT -38.320 598.430 -37.710 598.815 ;
        RECT -55.450 597.575 -54.955 598.385 ;
        RECT -55.450 597.405 -54.125 597.575 ;
        RECT -55.450 596.595 -54.955 597.405 ;
        RECT -55.450 596.425 -54.125 596.595 ;
        RECT -56.635 595.820 -55.665 596.415 ;
        RECT -57.265 595.790 -55.665 595.820 ;
        RECT -60.215 595.620 -55.665 595.790 ;
        RECT -57.265 595.595 -55.665 595.620 ;
        RECT -56.635 595.565 -55.665 595.595 ;
        RECT -56.515 595.540 -55.665 595.565 ;
        RECT -55.450 595.540 -54.955 596.425 ;
        RECT -56.515 595.510 -54.955 595.540 ;
        RECT -38.320 596.055 -12.635 598.430 ;
        RECT -56.515 595.340 -53.120 595.510 ;
        RECT -57.325 594.540 -56.830 594.780 ;
        RECT -58.155 594.370 -56.830 594.540 ;
        RECT -57.325 593.560 -56.830 594.370 ;
        RECT -58.155 593.390 -56.830 593.560 ;
        RECT -57.325 592.580 -56.830 593.390 ;
        RECT -58.155 592.410 -56.830 592.580 ;
        RECT -57.325 591.600 -56.830 592.410 ;
        RECT -58.155 591.430 -56.830 591.600 ;
        RECT -56.515 594.530 -55.205 595.340 ;
        RECT -56.515 594.360 -53.120 594.530 ;
        RECT -56.515 593.550 -55.205 594.360 ;
        RECT -38.320 594.195 -37.710 596.055 ;
        RECT -39.125 594.175 -37.710 594.195 ;
        RECT -40.585 594.005 -37.710 594.175 ;
        RECT -39.125 593.980 -37.710 594.005 ;
        RECT -56.515 593.380 -53.120 593.550 ;
        RECT -56.515 593.330 -55.205 593.380 ;
        RECT -56.515 593.325 -55.520 593.330 ;
        RECT -56.515 591.475 -55.750 593.325 ;
        RECT -38.325 593.210 -37.710 593.980 ;
        RECT -39.135 593.195 -37.710 593.210 ;
        RECT -40.585 593.025 -37.710 593.195 ;
        RECT -39.135 592.995 -37.710 593.025 ;
        RECT -38.325 592.090 -37.710 592.995 ;
        RECT -39.210 592.055 -37.710 592.090 ;
        RECT -41.585 591.885 -37.710 592.055 ;
        RECT -57.325 590.545 -56.830 591.430 ;
        RECT -57.325 590.515 -56.755 590.545 ;
        RECT -56.585 590.530 -55.750 591.475 ;
        RECT -59.160 590.345 -56.755 590.515 ;
        RECT -56.550 590.345 -55.750 590.530 ;
        RECT -57.075 589.535 -56.755 590.345 ;
        RECT -59.160 589.365 -56.755 589.535 ;
        RECT -57.075 588.555 -56.755 589.365 ;
        RECT -59.160 588.385 -56.755 588.555 ;
        RECT -57.075 588.335 -56.755 588.385 ;
        RECT -56.515 590.045 -55.750 590.345 ;
        RECT -54.800 591.625 -54.305 591.865 ;
        RECT -39.210 591.840 -37.710 591.885 ;
        RECT -54.800 591.455 -52.975 591.625 ;
        RECT -38.325 591.460 -37.710 591.840 ;
        RECT -54.800 590.645 -54.305 591.455 ;
        RECT -39.225 591.405 -37.710 591.460 ;
        RECT -41.585 591.235 -37.710 591.405 ;
        RECT -39.225 591.210 -37.710 591.235 ;
        RECT -54.800 590.475 -52.975 590.645 ;
        RECT -54.800 590.045 -54.305 590.475 ;
        RECT -56.515 589.665 -54.305 590.045 ;
        RECT -56.515 589.495 -52.975 589.665 ;
        RECT -56.515 589.185 -54.305 589.495 ;
        RECT -56.515 588.335 -55.750 589.185 ;
        RECT -54.800 588.685 -54.305 589.185 ;
        RECT -54.800 588.515 -52.975 588.685 ;
        RECT -56.250 584.660 -55.920 588.335 ;
        RECT -54.800 588.275 -54.305 588.515 ;
        RECT -38.325 588.440 -37.710 591.210 ;
        RECT -39.110 588.430 -37.710 588.440 ;
        RECT -41.585 588.260 -37.710 588.430 ;
        RECT -39.110 588.250 -37.710 588.260 ;
        RECT -38.325 587.455 -37.710 588.250 ;
        RECT -39.120 587.450 -37.710 587.455 ;
        RECT -41.585 587.280 -37.710 587.450 ;
        RECT -39.120 587.265 -37.710 587.280 ;
        RECT -38.645 586.015 -38.060 587.265 ;
        RECT -39.280 585.430 -38.060 586.015 ;
        RECT -56.250 584.330 -48.940 584.660 ;
        RECT -56.340 582.980 -55.775 582.985 ;
        RECT -49.270 582.980 -48.940 584.330 ;
        RECT -39.280 583.105 -38.695 585.430 ;
        RECT -56.340 582.650 -48.940 582.980 ;
        RECT -56.340 582.565 -55.775 582.650 ;
        RECT -39.310 582.615 -38.680 583.105 ;
        RECT -39.250 581.475 -38.780 581.785 ;
        RECT -55.295 581.195 -54.800 581.435 ;
        RECT -56.480 580.565 -56.150 581.070 ;
        RECT -57.100 580.550 -56.150 580.565 ;
        RECT -55.295 581.025 -53.970 581.195 ;
        RECT -39.180 581.110 -38.920 581.475 ;
        RECT -38.030 581.235 -37.535 581.475 ;
        RECT -57.100 580.545 -55.595 580.550 ;
        RECT -60.060 580.375 -55.595 580.545 ;
        RECT -57.100 580.340 -55.595 580.375 ;
        RECT -56.480 578.455 -55.595 580.340 ;
        RECT -57.095 578.430 -55.595 578.455 ;
        RECT -60.060 578.260 -55.595 578.430 ;
        RECT -57.095 578.230 -55.595 578.260 ;
        RECT -56.480 578.075 -55.595 578.230 ;
        RECT -55.295 580.215 -54.800 581.025 ;
        RECT -39.215 580.605 -38.885 581.110 ;
        RECT -39.835 580.590 -38.885 580.605 ;
        RECT -38.030 581.065 -36.705 581.235 ;
        RECT -39.835 580.585 -38.330 580.590 ;
        RECT -42.795 580.415 -38.330 580.585 ;
        RECT -39.835 580.380 -38.330 580.415 ;
        RECT -55.295 580.045 -53.970 580.215 ;
        RECT -55.295 579.235 -54.800 580.045 ;
        RECT -55.295 579.065 -53.970 579.235 ;
        RECT -55.295 578.255 -54.800 579.065 ;
        RECT -39.215 578.495 -38.330 580.380 ;
        RECT -39.830 578.470 -38.330 578.495 ;
        RECT -42.795 578.300 -38.330 578.470 ;
        RECT -39.830 578.270 -38.330 578.300 ;
        RECT -55.295 578.085 -53.970 578.255 ;
        RECT -39.215 578.115 -38.330 578.270 ;
        RECT -38.030 580.255 -37.535 581.065 ;
        RECT -38.030 580.085 -36.705 580.255 ;
        RECT -38.030 579.275 -37.535 580.085 ;
        RECT -38.030 579.105 -36.705 579.275 ;
        RECT -38.030 578.295 -37.535 579.105 ;
        RECT -38.030 578.125 -36.705 578.295 ;
        RECT -56.480 577.480 -55.510 578.075 ;
        RECT -57.110 577.450 -55.510 577.480 ;
        RECT -60.060 577.280 -55.510 577.450 ;
        RECT -57.110 577.255 -55.510 577.280 ;
        RECT -56.480 577.225 -55.510 577.255 ;
        RECT -56.360 577.200 -55.510 577.225 ;
        RECT -55.295 577.200 -54.800 578.085 ;
        RECT -39.215 577.520 -38.245 578.115 ;
        RECT -39.845 577.490 -38.245 577.520 ;
        RECT -42.795 577.320 -38.245 577.490 ;
        RECT -39.845 577.295 -38.245 577.320 ;
        RECT -39.215 577.265 -38.245 577.295 ;
        RECT -56.360 577.170 -54.800 577.200 ;
        RECT -39.095 577.240 -38.245 577.265 ;
        RECT -38.030 577.240 -37.535 578.125 ;
        RECT -39.095 577.210 -37.535 577.240 ;
        RECT -56.360 577.000 -52.965 577.170 ;
        RECT -39.095 577.040 -35.700 577.210 ;
        RECT -57.170 576.200 -56.675 576.440 ;
        RECT -58.000 576.030 -56.675 576.200 ;
        RECT -57.170 575.220 -56.675 576.030 ;
        RECT -58.000 575.050 -56.675 575.220 ;
        RECT -57.170 574.240 -56.675 575.050 ;
        RECT -58.000 574.070 -56.675 574.240 ;
        RECT -57.170 573.260 -56.675 574.070 ;
        RECT -58.000 573.090 -56.675 573.260 ;
        RECT -56.360 576.190 -55.050 577.000 ;
        RECT -39.905 576.240 -39.410 576.480 ;
        RECT -56.360 576.020 -52.965 576.190 ;
        RECT -40.735 576.070 -39.410 576.240 ;
        RECT -56.360 575.210 -55.050 576.020 ;
        RECT -39.905 575.260 -39.410 576.070 ;
        RECT -56.360 575.040 -52.965 575.210 ;
        RECT -40.735 575.090 -39.410 575.260 ;
        RECT -56.360 574.990 -55.050 575.040 ;
        RECT -56.360 574.985 -55.365 574.990 ;
        RECT -56.360 573.135 -55.595 574.985 ;
        RECT -39.905 574.280 -39.410 575.090 ;
        RECT -40.735 574.110 -39.410 574.280 ;
        RECT -57.170 572.205 -56.675 573.090 ;
        RECT -57.170 572.175 -56.600 572.205 ;
        RECT -56.430 572.190 -55.595 573.135 ;
        RECT -59.005 572.005 -56.600 572.175 ;
        RECT -56.395 572.005 -55.595 572.190 ;
        RECT -56.920 571.195 -56.600 572.005 ;
        RECT -59.005 571.025 -56.600 571.195 ;
        RECT -56.920 570.215 -56.600 571.025 ;
        RECT -59.005 570.045 -56.600 570.215 ;
        RECT -56.920 569.995 -56.600 570.045 ;
        RECT -56.360 571.705 -55.595 572.005 ;
        RECT -54.645 573.285 -54.150 573.525 ;
        RECT -39.905 573.300 -39.410 574.110 ;
        RECT -54.645 573.115 -52.820 573.285 ;
        RECT -40.735 573.130 -39.410 573.300 ;
        RECT -39.095 576.230 -37.785 577.040 ;
        RECT -39.095 576.060 -35.700 576.230 ;
        RECT -39.095 575.250 -37.785 576.060 ;
        RECT -39.095 575.080 -35.700 575.250 ;
        RECT -39.095 575.030 -37.785 575.080 ;
        RECT -39.095 575.025 -38.100 575.030 ;
        RECT -39.095 573.175 -38.330 575.025 ;
        RECT -54.645 572.305 -54.150 573.115 ;
        RECT -54.645 572.135 -52.820 572.305 ;
        RECT -39.905 572.245 -39.410 573.130 ;
        RECT -39.905 572.215 -39.335 572.245 ;
        RECT -39.165 572.230 -38.330 573.175 ;
        RECT -54.645 571.705 -54.150 572.135 ;
        RECT -41.740 572.045 -39.335 572.215 ;
        RECT -39.130 572.045 -38.330 572.230 ;
        RECT -56.360 571.325 -54.150 571.705 ;
        RECT -56.360 571.155 -52.820 571.325 ;
        RECT -39.655 571.235 -39.335 572.045 ;
        RECT -56.360 570.845 -54.150 571.155 ;
        RECT -41.740 571.065 -39.335 571.235 ;
        RECT -56.360 569.995 -55.595 570.845 ;
        RECT -54.645 570.345 -54.150 570.845 ;
        RECT -54.645 570.175 -52.820 570.345 ;
        RECT -39.655 570.255 -39.335 571.065 ;
        RECT -54.645 569.935 -54.150 570.175 ;
        RECT -41.740 570.085 -39.335 570.255 ;
        RECT -39.655 570.035 -39.335 570.085 ;
        RECT -39.095 571.745 -38.330 572.045 ;
        RECT -37.380 573.325 -36.885 573.565 ;
        RECT -37.380 573.155 -35.555 573.325 ;
        RECT -37.380 572.345 -36.885 573.155 ;
        RECT -37.380 572.175 -35.555 572.345 ;
        RECT -37.380 571.745 -36.885 572.175 ;
        RECT -39.095 571.365 -36.885 571.745 ;
        RECT -39.095 571.195 -35.555 571.365 ;
        RECT -39.095 570.385 -36.885 571.195 ;
        RECT -39.095 570.215 -35.555 570.385 ;
        RECT -39.095 570.035 -36.885 570.215 ;
        RECT -38.815 569.975 -36.885 570.035 ;
        RECT -56.780 554.790 -50.495 555.155 ;
        RECT -56.920 554.545 -50.495 554.790 ;
        RECT -56.920 554.095 -56.085 554.545 ;
        RECT -56.855 552.845 -56.160 553.240 ;
        RECT -56.730 552.590 -56.315 552.845 ;
        RECT -56.825 552.345 -56.315 552.590 ;
        RECT -55.640 552.715 -55.145 552.955 ;
        RECT -55.640 552.545 -54.315 552.715 ;
        RECT -51.105 552.605 -50.495 554.545 ;
        RECT -38.815 552.605 -37.105 569.975 ;
        RECT -56.825 552.085 -56.495 552.345 ;
        RECT -57.445 552.070 -56.495 552.085 ;
        RECT -57.445 552.065 -55.940 552.070 ;
        RECT -60.405 551.895 -55.940 552.065 ;
        RECT -57.445 551.860 -55.940 551.895 ;
        RECT -56.825 549.975 -55.940 551.860 ;
        RECT -57.440 549.950 -55.940 549.975 ;
        RECT -60.405 549.780 -55.940 549.950 ;
        RECT -57.440 549.750 -55.940 549.780 ;
        RECT -56.825 549.595 -55.940 549.750 ;
        RECT -55.640 551.735 -55.145 552.545 ;
        RECT -51.105 551.995 -37.105 552.605 ;
        RECT -55.640 551.565 -54.315 551.735 ;
        RECT -55.640 550.755 -55.145 551.565 ;
        RECT -55.640 550.585 -54.315 550.755 ;
        RECT -55.640 549.775 -55.145 550.585 ;
        RECT -55.640 549.605 -54.315 549.775 ;
        RECT -56.825 549.000 -55.855 549.595 ;
        RECT -57.455 548.970 -55.855 549.000 ;
        RECT -60.405 548.800 -55.855 548.970 ;
        RECT -57.455 548.775 -55.855 548.800 ;
        RECT -56.825 548.745 -55.855 548.775 ;
        RECT -56.705 548.720 -55.855 548.745 ;
        RECT -55.640 548.720 -55.145 549.605 ;
        RECT -56.705 548.690 -55.145 548.720 ;
        RECT -56.705 548.520 -53.310 548.690 ;
        RECT -57.515 547.720 -57.020 547.960 ;
        RECT -58.345 547.550 -57.020 547.720 ;
        RECT -57.515 546.740 -57.020 547.550 ;
        RECT -58.345 546.570 -57.020 546.740 ;
        RECT -57.515 545.760 -57.020 546.570 ;
        RECT -58.345 545.590 -57.020 545.760 ;
        RECT -57.515 544.780 -57.020 545.590 ;
        RECT -58.345 544.610 -57.020 544.780 ;
        RECT -56.705 547.710 -55.395 548.520 ;
        RECT -56.705 547.540 -53.310 547.710 ;
        RECT -56.705 546.730 -55.395 547.540 ;
        RECT -38.815 547.375 -37.105 551.995 ;
        RECT -39.315 547.355 -37.105 547.375 ;
        RECT -40.775 547.185 -37.105 547.355 ;
        RECT -39.315 547.180 -37.105 547.185 ;
        RECT -39.315 547.160 -37.900 547.180 ;
        RECT -56.705 546.560 -53.310 546.730 ;
        RECT -56.705 546.510 -55.395 546.560 ;
        RECT -56.705 546.505 -55.710 546.510 ;
        RECT -56.705 544.655 -55.940 546.505 ;
        RECT -38.515 546.390 -37.900 547.160 ;
        RECT -39.325 546.375 -37.900 546.390 ;
        RECT -40.775 546.205 -37.900 546.375 ;
        RECT -39.325 546.175 -37.900 546.205 ;
        RECT -38.515 545.270 -37.900 546.175 ;
        RECT -39.400 545.235 -37.900 545.270 ;
        RECT -41.775 545.065 -37.900 545.235 ;
        RECT -57.515 543.725 -57.020 544.610 ;
        RECT -57.515 543.695 -56.945 543.725 ;
        RECT -56.775 543.710 -55.940 544.655 ;
        RECT -59.350 543.525 -56.945 543.695 ;
        RECT -56.740 543.525 -55.940 543.710 ;
        RECT -57.265 542.715 -56.945 543.525 ;
        RECT -59.350 542.545 -56.945 542.715 ;
        RECT -57.265 541.735 -56.945 542.545 ;
        RECT -59.350 541.565 -56.945 541.735 ;
        RECT -57.265 541.515 -56.945 541.565 ;
        RECT -56.705 543.225 -55.940 543.525 ;
        RECT -54.990 544.805 -54.495 545.045 ;
        RECT -39.400 545.020 -37.900 545.065 ;
        RECT -54.990 544.635 -53.165 544.805 ;
        RECT -38.515 544.640 -37.900 545.020 ;
        RECT -54.990 543.825 -54.495 544.635 ;
        RECT -39.415 544.585 -37.900 544.640 ;
        RECT -41.775 544.415 -37.900 544.585 ;
        RECT -39.415 544.390 -37.900 544.415 ;
        RECT -54.990 543.655 -53.165 543.825 ;
        RECT -54.990 543.225 -54.495 543.655 ;
        RECT -56.705 542.845 -54.495 543.225 ;
        RECT -56.705 542.675 -53.165 542.845 ;
        RECT -56.705 542.365 -54.495 542.675 ;
        RECT -56.705 541.515 -55.940 542.365 ;
        RECT -54.990 541.865 -54.495 542.365 ;
        RECT -54.990 541.695 -53.165 541.865 ;
        RECT -56.440 537.840 -56.110 541.515 ;
        RECT -54.990 541.455 -54.495 541.695 ;
        RECT -38.515 541.620 -37.900 544.390 ;
        RECT -39.300 541.610 -37.900 541.620 ;
        RECT -41.775 541.440 -37.900 541.610 ;
        RECT -39.300 541.430 -37.900 541.440 ;
        RECT -38.515 540.635 -37.900 541.430 ;
        RECT -39.310 540.630 -37.900 540.635 ;
        RECT -41.775 540.460 -37.900 540.630 ;
        RECT -39.310 540.445 -37.900 540.460 ;
        RECT -38.835 539.195 -38.250 540.445 ;
        RECT -39.470 538.610 -38.250 539.195 ;
        RECT -56.440 537.510 -49.130 537.840 ;
        RECT -56.530 536.160 -55.965 536.165 ;
        RECT -49.460 536.160 -49.130 537.510 ;
        RECT -39.470 536.285 -38.885 538.610 ;
        RECT -56.530 535.830 -49.130 536.160 ;
        RECT -56.530 535.745 -55.965 535.830 ;
        RECT -39.500 535.795 -38.870 536.285 ;
        RECT -39.440 534.655 -38.970 534.965 ;
        RECT -55.485 534.375 -54.990 534.615 ;
        RECT -56.670 533.745 -56.340 534.250 ;
        RECT -57.290 533.730 -56.340 533.745 ;
        RECT -55.485 534.205 -54.160 534.375 ;
        RECT -39.370 534.290 -39.110 534.655 ;
        RECT -38.220 534.415 -37.725 534.655 ;
        RECT -57.290 533.725 -55.785 533.730 ;
        RECT -60.250 533.555 -55.785 533.725 ;
        RECT -57.290 533.520 -55.785 533.555 ;
        RECT -56.670 531.635 -55.785 533.520 ;
        RECT -57.285 531.610 -55.785 531.635 ;
        RECT -60.250 531.440 -55.785 531.610 ;
        RECT -57.285 531.410 -55.785 531.440 ;
        RECT -56.670 531.255 -55.785 531.410 ;
        RECT -55.485 533.395 -54.990 534.205 ;
        RECT -39.405 533.785 -39.075 534.290 ;
        RECT -40.025 533.770 -39.075 533.785 ;
        RECT -38.220 534.245 -36.895 534.415 ;
        RECT -40.025 533.765 -38.520 533.770 ;
        RECT -42.985 533.595 -38.520 533.765 ;
        RECT -40.025 533.560 -38.520 533.595 ;
        RECT -55.485 533.225 -54.160 533.395 ;
        RECT -55.485 532.415 -54.990 533.225 ;
        RECT -55.485 532.245 -54.160 532.415 ;
        RECT -55.485 531.435 -54.990 532.245 ;
        RECT -39.405 531.675 -38.520 533.560 ;
        RECT -40.020 531.650 -38.520 531.675 ;
        RECT -42.985 531.480 -38.520 531.650 ;
        RECT -40.020 531.450 -38.520 531.480 ;
        RECT -55.485 531.265 -54.160 531.435 ;
        RECT -39.405 531.295 -38.520 531.450 ;
        RECT -38.220 533.435 -37.725 534.245 ;
        RECT -38.220 533.265 -36.895 533.435 ;
        RECT -38.220 532.455 -37.725 533.265 ;
        RECT -38.220 532.285 -36.895 532.455 ;
        RECT -38.220 531.475 -37.725 532.285 ;
        RECT -38.220 531.305 -36.895 531.475 ;
        RECT -56.670 530.660 -55.700 531.255 ;
        RECT -57.300 530.630 -55.700 530.660 ;
        RECT -60.250 530.460 -55.700 530.630 ;
        RECT -57.300 530.435 -55.700 530.460 ;
        RECT -56.670 530.405 -55.700 530.435 ;
        RECT -56.550 530.380 -55.700 530.405 ;
        RECT -55.485 530.380 -54.990 531.265 ;
        RECT -39.405 530.700 -38.435 531.295 ;
        RECT -40.035 530.670 -38.435 530.700 ;
        RECT -42.985 530.500 -38.435 530.670 ;
        RECT -40.035 530.475 -38.435 530.500 ;
        RECT -39.405 530.445 -38.435 530.475 ;
        RECT -56.550 530.350 -54.990 530.380 ;
        RECT -39.285 530.420 -38.435 530.445 ;
        RECT -38.220 530.420 -37.725 531.305 ;
        RECT -39.285 530.390 -37.725 530.420 ;
        RECT -56.550 530.180 -53.155 530.350 ;
        RECT -39.285 530.220 -35.890 530.390 ;
        RECT -57.360 529.380 -56.865 529.620 ;
        RECT -58.190 529.210 -56.865 529.380 ;
        RECT -57.360 528.400 -56.865 529.210 ;
        RECT -58.190 528.230 -56.865 528.400 ;
        RECT -57.360 527.420 -56.865 528.230 ;
        RECT -58.190 527.250 -56.865 527.420 ;
        RECT -57.360 526.440 -56.865 527.250 ;
        RECT -58.190 526.270 -56.865 526.440 ;
        RECT -56.550 529.370 -55.240 530.180 ;
        RECT -40.095 529.420 -39.600 529.660 ;
        RECT -56.550 529.200 -53.155 529.370 ;
        RECT -40.925 529.250 -39.600 529.420 ;
        RECT -56.550 528.390 -55.240 529.200 ;
        RECT -40.095 528.440 -39.600 529.250 ;
        RECT -56.550 528.220 -53.155 528.390 ;
        RECT -40.925 528.270 -39.600 528.440 ;
        RECT -56.550 528.170 -55.240 528.220 ;
        RECT -56.550 528.165 -55.555 528.170 ;
        RECT -56.550 526.315 -55.785 528.165 ;
        RECT -40.095 527.460 -39.600 528.270 ;
        RECT -40.925 527.290 -39.600 527.460 ;
        RECT -57.360 525.385 -56.865 526.270 ;
        RECT -57.360 525.355 -56.790 525.385 ;
        RECT -56.620 525.370 -55.785 526.315 ;
        RECT -59.195 525.185 -56.790 525.355 ;
        RECT -56.585 525.185 -55.785 525.370 ;
        RECT -57.110 524.375 -56.790 525.185 ;
        RECT -59.195 524.205 -56.790 524.375 ;
        RECT -57.110 523.395 -56.790 524.205 ;
        RECT -59.195 523.225 -56.790 523.395 ;
        RECT -57.110 523.175 -56.790 523.225 ;
        RECT -56.550 524.885 -55.785 525.185 ;
        RECT -54.835 526.465 -54.340 526.705 ;
        RECT -40.095 526.480 -39.600 527.290 ;
        RECT -54.835 526.295 -53.010 526.465 ;
        RECT -40.925 526.310 -39.600 526.480 ;
        RECT -39.285 529.410 -37.975 530.220 ;
        RECT -39.285 529.240 -35.890 529.410 ;
        RECT -39.285 528.430 -37.975 529.240 ;
        RECT -39.285 528.260 -35.890 528.430 ;
        RECT -39.285 528.210 -37.975 528.260 ;
        RECT -39.285 528.205 -38.290 528.210 ;
        RECT -39.285 526.355 -38.520 528.205 ;
        RECT -54.835 525.485 -54.340 526.295 ;
        RECT -54.835 525.315 -53.010 525.485 ;
        RECT -40.095 525.425 -39.600 526.310 ;
        RECT -40.095 525.395 -39.525 525.425 ;
        RECT -39.355 525.410 -38.520 526.355 ;
        RECT -54.835 524.885 -54.340 525.315 ;
        RECT -41.930 525.225 -39.525 525.395 ;
        RECT -39.320 525.225 -38.520 525.410 ;
        RECT -56.550 524.505 -54.340 524.885 ;
        RECT -56.550 524.335 -53.010 524.505 ;
        RECT -39.845 524.415 -39.525 525.225 ;
        RECT -56.550 524.025 -54.340 524.335 ;
        RECT -41.930 524.245 -39.525 524.415 ;
        RECT -56.550 523.175 -55.785 524.025 ;
        RECT -54.835 523.525 -54.340 524.025 ;
        RECT -54.835 523.355 -53.010 523.525 ;
        RECT -39.845 523.435 -39.525 524.245 ;
        RECT -54.835 523.115 -54.340 523.355 ;
        RECT -41.930 523.265 -39.525 523.435 ;
        RECT -39.845 523.215 -39.525 523.265 ;
        RECT -39.285 524.925 -38.520 525.225 ;
        RECT -37.570 526.505 -37.075 526.745 ;
        RECT -37.570 526.335 -35.745 526.505 ;
        RECT -37.570 525.525 -37.075 526.335 ;
        RECT -37.570 525.355 -35.745 525.525 ;
        RECT -37.570 524.925 -37.075 525.355 ;
        RECT -39.285 524.545 -37.075 524.925 ;
        RECT -39.285 524.375 -35.745 524.545 ;
        RECT -39.285 523.565 -37.075 524.375 ;
        RECT -39.285 523.395 -35.745 523.565 ;
        RECT -39.285 523.215 -37.075 523.395 ;
        RECT -38.770 523.155 -37.075 523.215 ;
        RECT -56.865 509.025 -50.580 509.390 ;
        RECT -57.005 508.780 -50.580 509.025 ;
        RECT -57.005 508.330 -56.170 508.780 ;
        RECT -56.940 507.080 -56.245 507.475 ;
        RECT -56.815 506.825 -56.400 507.080 ;
        RECT -56.910 506.580 -56.400 506.825 ;
        RECT -55.725 506.950 -55.230 507.190 ;
        RECT -55.725 506.780 -54.400 506.950 ;
        RECT -51.190 506.840 -50.580 508.780 ;
        RECT -38.770 506.840 -37.450 523.155 ;
        RECT -56.910 506.320 -56.580 506.580 ;
        RECT -57.530 506.305 -56.580 506.320 ;
        RECT -57.530 506.300 -56.025 506.305 ;
        RECT -60.490 506.130 -56.025 506.300 ;
        RECT -57.530 506.095 -56.025 506.130 ;
        RECT -56.910 504.210 -56.025 506.095 ;
        RECT -57.525 504.185 -56.025 504.210 ;
        RECT -60.490 504.015 -56.025 504.185 ;
        RECT -57.525 503.985 -56.025 504.015 ;
        RECT -56.910 503.830 -56.025 503.985 ;
        RECT -55.725 505.970 -55.230 506.780 ;
        RECT -51.190 506.230 -37.450 506.840 ;
        RECT -55.725 505.800 -54.400 505.970 ;
        RECT -55.725 504.990 -55.230 505.800 ;
        RECT -55.725 504.820 -54.400 504.990 ;
        RECT -55.725 504.010 -55.230 504.820 ;
        RECT -55.725 503.840 -54.400 504.010 ;
        RECT -56.910 503.235 -55.940 503.830 ;
        RECT -57.540 503.205 -55.940 503.235 ;
        RECT -60.490 503.035 -55.940 503.205 ;
        RECT -57.540 503.010 -55.940 503.035 ;
        RECT -56.910 502.980 -55.940 503.010 ;
        RECT -56.790 502.955 -55.940 502.980 ;
        RECT -55.725 502.955 -55.230 503.840 ;
        RECT -56.790 502.925 -55.230 502.955 ;
        RECT -56.790 502.755 -53.395 502.925 ;
        RECT -57.600 501.955 -57.105 502.195 ;
        RECT -58.430 501.785 -57.105 501.955 ;
        RECT -57.600 500.975 -57.105 501.785 ;
        RECT -58.430 500.805 -57.105 500.975 ;
        RECT -57.600 499.995 -57.105 500.805 ;
        RECT -58.430 499.825 -57.105 499.995 ;
        RECT -57.600 499.015 -57.105 499.825 ;
        RECT -58.430 498.845 -57.105 499.015 ;
        RECT -56.790 501.945 -55.480 502.755 ;
        RECT -56.790 501.775 -53.395 501.945 ;
        RECT -56.790 500.965 -55.480 501.775 ;
        RECT -38.770 501.610 -37.450 506.230 ;
        RECT -39.400 501.590 -37.450 501.610 ;
        RECT -40.860 501.420 -37.450 501.590 ;
        RECT -39.400 501.395 -37.450 501.420 ;
        RECT -38.770 501.370 -37.450 501.395 ;
        RECT -56.790 500.795 -53.395 500.965 ;
        RECT -56.790 500.745 -55.480 500.795 ;
        RECT -56.790 500.740 -55.795 500.745 ;
        RECT -56.790 498.890 -56.025 500.740 ;
        RECT -38.600 500.625 -37.985 501.370 ;
        RECT -39.410 500.610 -37.985 500.625 ;
        RECT -40.860 500.440 -37.985 500.610 ;
        RECT -39.410 500.410 -37.985 500.440 ;
        RECT -38.600 499.505 -37.985 500.410 ;
        RECT -39.485 499.470 -37.985 499.505 ;
        RECT -41.860 499.300 -37.985 499.470 ;
        RECT -57.600 497.960 -57.105 498.845 ;
        RECT -57.600 497.930 -57.030 497.960 ;
        RECT -56.860 497.945 -56.025 498.890 ;
        RECT -59.435 497.760 -57.030 497.930 ;
        RECT -56.825 497.760 -56.025 497.945 ;
        RECT -57.350 496.950 -57.030 497.760 ;
        RECT -59.435 496.780 -57.030 496.950 ;
        RECT -57.350 495.970 -57.030 496.780 ;
        RECT -59.435 495.800 -57.030 495.970 ;
        RECT -57.350 495.750 -57.030 495.800 ;
        RECT -56.790 497.460 -56.025 497.760 ;
        RECT -55.075 499.040 -54.580 499.280 ;
        RECT -39.485 499.255 -37.985 499.300 ;
        RECT -55.075 498.870 -53.250 499.040 ;
        RECT -38.600 498.875 -37.985 499.255 ;
        RECT -55.075 498.060 -54.580 498.870 ;
        RECT -39.500 498.820 -37.985 498.875 ;
        RECT -41.860 498.650 -37.985 498.820 ;
        RECT -39.500 498.625 -37.985 498.650 ;
        RECT -55.075 497.890 -53.250 498.060 ;
        RECT -55.075 497.460 -54.580 497.890 ;
        RECT -56.790 497.080 -54.580 497.460 ;
        RECT -56.790 496.910 -53.250 497.080 ;
        RECT -56.790 496.600 -54.580 496.910 ;
        RECT -56.790 495.750 -56.025 496.600 ;
        RECT -55.075 496.100 -54.580 496.600 ;
        RECT -55.075 495.930 -53.250 496.100 ;
        RECT -56.525 492.075 -56.195 495.750 ;
        RECT -55.075 495.690 -54.580 495.930 ;
        RECT -38.600 495.855 -37.985 498.625 ;
        RECT -39.385 495.845 -37.985 495.855 ;
        RECT -41.860 495.675 -37.985 495.845 ;
        RECT -39.385 495.665 -37.985 495.675 ;
        RECT -38.600 494.870 -37.985 495.665 ;
        RECT -39.395 494.865 -37.985 494.870 ;
        RECT -41.860 494.695 -37.985 494.865 ;
        RECT -39.395 494.680 -37.985 494.695 ;
        RECT -38.920 493.430 -38.335 494.680 ;
        RECT -39.555 492.845 -38.335 493.430 ;
        RECT -56.525 491.745 -49.215 492.075 ;
        RECT -56.615 490.395 -56.050 490.400 ;
        RECT -49.545 490.395 -49.215 491.745 ;
        RECT -39.555 490.520 -38.970 492.845 ;
        RECT -56.615 490.065 -49.215 490.395 ;
        RECT -56.615 489.980 -56.050 490.065 ;
        RECT -39.585 490.030 -38.955 490.520 ;
        RECT -39.525 488.890 -39.055 489.200 ;
        RECT -55.570 488.610 -55.075 488.850 ;
        RECT -56.755 487.980 -56.425 488.485 ;
        RECT -57.375 487.965 -56.425 487.980 ;
        RECT -55.570 488.440 -54.245 488.610 ;
        RECT -39.455 488.525 -39.195 488.890 ;
        RECT -38.305 488.650 -37.810 488.890 ;
        RECT -57.375 487.960 -55.870 487.965 ;
        RECT -60.335 487.790 -55.870 487.960 ;
        RECT -57.375 487.755 -55.870 487.790 ;
        RECT -56.755 485.870 -55.870 487.755 ;
        RECT -57.370 485.845 -55.870 485.870 ;
        RECT -60.335 485.675 -55.870 485.845 ;
        RECT -57.370 485.645 -55.870 485.675 ;
        RECT -56.755 485.490 -55.870 485.645 ;
        RECT -55.570 487.630 -55.075 488.440 ;
        RECT -39.490 488.020 -39.160 488.525 ;
        RECT -40.110 488.005 -39.160 488.020 ;
        RECT -38.305 488.480 -36.980 488.650 ;
        RECT -40.110 488.000 -38.605 488.005 ;
        RECT -43.070 487.830 -38.605 488.000 ;
        RECT -40.110 487.795 -38.605 487.830 ;
        RECT -55.570 487.460 -54.245 487.630 ;
        RECT -55.570 486.650 -55.075 487.460 ;
        RECT -55.570 486.480 -54.245 486.650 ;
        RECT -55.570 485.670 -55.075 486.480 ;
        RECT -39.490 485.910 -38.605 487.795 ;
        RECT -40.105 485.885 -38.605 485.910 ;
        RECT -43.070 485.715 -38.605 485.885 ;
        RECT -40.105 485.685 -38.605 485.715 ;
        RECT -55.570 485.500 -54.245 485.670 ;
        RECT -39.490 485.530 -38.605 485.685 ;
        RECT -38.305 487.670 -37.810 488.480 ;
        RECT -38.305 487.500 -36.980 487.670 ;
        RECT -38.305 486.690 -37.810 487.500 ;
        RECT -38.305 486.520 -36.980 486.690 ;
        RECT -38.305 485.710 -37.810 486.520 ;
        RECT -38.305 485.540 -36.980 485.710 ;
        RECT -56.755 484.895 -55.785 485.490 ;
        RECT -57.385 484.865 -55.785 484.895 ;
        RECT -60.335 484.695 -55.785 484.865 ;
        RECT -57.385 484.670 -55.785 484.695 ;
        RECT -56.755 484.640 -55.785 484.670 ;
        RECT -56.635 484.615 -55.785 484.640 ;
        RECT -55.570 484.615 -55.075 485.500 ;
        RECT -39.490 484.935 -38.520 485.530 ;
        RECT -40.120 484.905 -38.520 484.935 ;
        RECT -43.070 484.735 -38.520 484.905 ;
        RECT -40.120 484.710 -38.520 484.735 ;
        RECT -39.490 484.680 -38.520 484.710 ;
        RECT -56.635 484.585 -55.075 484.615 ;
        RECT -39.370 484.655 -38.520 484.680 ;
        RECT -38.305 484.655 -37.810 485.540 ;
        RECT -39.370 484.625 -37.810 484.655 ;
        RECT -56.635 484.415 -53.240 484.585 ;
        RECT -39.370 484.455 -35.975 484.625 ;
        RECT -57.445 483.615 -56.950 483.855 ;
        RECT -58.275 483.445 -56.950 483.615 ;
        RECT -57.445 482.635 -56.950 483.445 ;
        RECT -58.275 482.465 -56.950 482.635 ;
        RECT -57.445 481.655 -56.950 482.465 ;
        RECT -58.275 481.485 -56.950 481.655 ;
        RECT -57.445 480.675 -56.950 481.485 ;
        RECT -58.275 480.505 -56.950 480.675 ;
        RECT -56.635 483.605 -55.325 484.415 ;
        RECT -40.180 483.655 -39.685 483.895 ;
        RECT -56.635 483.435 -53.240 483.605 ;
        RECT -41.010 483.485 -39.685 483.655 ;
        RECT -56.635 482.625 -55.325 483.435 ;
        RECT -40.180 482.675 -39.685 483.485 ;
        RECT -56.635 482.455 -53.240 482.625 ;
        RECT -41.010 482.505 -39.685 482.675 ;
        RECT -56.635 482.405 -55.325 482.455 ;
        RECT -56.635 482.400 -55.640 482.405 ;
        RECT -56.635 480.550 -55.870 482.400 ;
        RECT -40.180 481.695 -39.685 482.505 ;
        RECT -41.010 481.525 -39.685 481.695 ;
        RECT -57.445 479.620 -56.950 480.505 ;
        RECT -57.445 479.590 -56.875 479.620 ;
        RECT -56.705 479.605 -55.870 480.550 ;
        RECT -59.280 479.420 -56.875 479.590 ;
        RECT -56.670 479.420 -55.870 479.605 ;
        RECT -57.195 478.610 -56.875 479.420 ;
        RECT -59.280 478.440 -56.875 478.610 ;
        RECT -57.195 477.630 -56.875 478.440 ;
        RECT -59.280 477.460 -56.875 477.630 ;
        RECT -57.195 477.410 -56.875 477.460 ;
        RECT -56.635 479.120 -55.870 479.420 ;
        RECT -54.920 480.700 -54.425 480.940 ;
        RECT -40.180 480.715 -39.685 481.525 ;
        RECT -54.920 480.530 -53.095 480.700 ;
        RECT -41.010 480.545 -39.685 480.715 ;
        RECT -39.370 483.645 -38.060 484.455 ;
        RECT -39.370 483.475 -35.975 483.645 ;
        RECT -39.370 482.665 -38.060 483.475 ;
        RECT -39.370 482.495 -35.975 482.665 ;
        RECT -39.370 482.445 -38.060 482.495 ;
        RECT -39.370 482.440 -38.375 482.445 ;
        RECT -39.370 480.590 -38.605 482.440 ;
        RECT -54.920 479.720 -54.425 480.530 ;
        RECT -54.920 479.550 -53.095 479.720 ;
        RECT -40.180 479.660 -39.685 480.545 ;
        RECT -40.180 479.630 -39.610 479.660 ;
        RECT -39.440 479.645 -38.605 480.590 ;
        RECT -54.920 479.120 -54.425 479.550 ;
        RECT -42.015 479.460 -39.610 479.630 ;
        RECT -39.405 479.460 -38.605 479.645 ;
        RECT -56.635 478.740 -54.425 479.120 ;
        RECT -56.635 478.570 -53.095 478.740 ;
        RECT -39.930 478.650 -39.610 479.460 ;
        RECT -56.635 478.260 -54.425 478.570 ;
        RECT -42.015 478.480 -39.610 478.650 ;
        RECT -56.635 477.410 -55.870 478.260 ;
        RECT -54.920 477.760 -54.425 478.260 ;
        RECT -54.920 477.590 -53.095 477.760 ;
        RECT -39.930 477.670 -39.610 478.480 ;
        RECT -54.920 477.350 -54.425 477.590 ;
        RECT -42.015 477.500 -39.610 477.670 ;
        RECT -39.930 477.450 -39.610 477.500 ;
        RECT -39.370 479.160 -38.605 479.460 ;
        RECT -37.655 480.740 -37.160 480.980 ;
        RECT -37.655 480.570 -35.830 480.740 ;
        RECT -37.655 479.760 -37.160 480.570 ;
        RECT -37.655 479.590 -35.830 479.760 ;
        RECT -37.655 479.160 -37.160 479.590 ;
        RECT -39.370 478.780 -37.160 479.160 ;
        RECT -39.370 478.610 -35.830 478.780 ;
        RECT -39.370 477.800 -37.160 478.610 ;
        RECT -39.370 477.630 -35.830 477.800 ;
        RECT -39.370 477.450 -37.160 477.630 ;
        RECT -39.240 477.390 -37.160 477.450 ;
        RECT -57.195 465.255 -50.910 465.620 ;
        RECT -57.335 465.010 -50.910 465.255 ;
        RECT -57.335 464.560 -56.500 465.010 ;
        RECT -57.270 463.310 -56.575 463.705 ;
        RECT -57.145 463.055 -56.730 463.310 ;
        RECT -57.240 462.810 -56.730 463.055 ;
        RECT -56.055 463.180 -55.560 463.420 ;
        RECT -56.055 463.010 -54.730 463.180 ;
        RECT -51.520 463.070 -50.910 465.010 ;
        RECT -39.240 463.070 -37.345 477.390 ;
        RECT -57.240 462.550 -56.910 462.810 ;
        RECT -57.860 462.535 -56.910 462.550 ;
        RECT -57.860 462.530 -56.355 462.535 ;
        RECT -60.820 462.360 -56.355 462.530 ;
        RECT -57.860 462.325 -56.355 462.360 ;
        RECT -57.240 460.440 -56.355 462.325 ;
        RECT -57.855 460.415 -56.355 460.440 ;
        RECT -60.820 460.245 -56.355 460.415 ;
        RECT -57.855 460.215 -56.355 460.245 ;
        RECT -57.240 460.060 -56.355 460.215 ;
        RECT -56.055 462.200 -55.560 463.010 ;
        RECT -51.520 462.460 -37.345 463.070 ;
        RECT -56.055 462.030 -54.730 462.200 ;
        RECT -56.055 461.220 -55.560 462.030 ;
        RECT -56.055 461.050 -54.730 461.220 ;
        RECT -56.055 460.240 -55.560 461.050 ;
        RECT -56.055 460.070 -54.730 460.240 ;
        RECT -57.240 459.465 -56.270 460.060 ;
        RECT -57.870 459.435 -56.270 459.465 ;
        RECT -60.820 459.265 -56.270 459.435 ;
        RECT -57.870 459.240 -56.270 459.265 ;
        RECT -57.240 459.210 -56.270 459.240 ;
        RECT -57.120 459.185 -56.270 459.210 ;
        RECT -56.055 459.185 -55.560 460.070 ;
        RECT -57.120 459.155 -55.560 459.185 ;
        RECT -57.120 458.985 -53.725 459.155 ;
        RECT -57.930 458.185 -57.435 458.425 ;
        RECT -58.760 458.015 -57.435 458.185 ;
        RECT -57.930 457.205 -57.435 458.015 ;
        RECT -58.760 457.035 -57.435 457.205 ;
        RECT -57.930 456.225 -57.435 457.035 ;
        RECT -58.760 456.055 -57.435 456.225 ;
        RECT -57.930 455.245 -57.435 456.055 ;
        RECT -58.760 455.075 -57.435 455.245 ;
        RECT -57.120 458.175 -55.810 458.985 ;
        RECT -57.120 458.005 -53.725 458.175 ;
        RECT -57.120 457.195 -55.810 458.005 ;
        RECT -39.240 457.840 -37.345 462.460 ;
        RECT -39.730 457.820 -37.345 457.840 ;
        RECT -41.190 457.650 -37.345 457.820 ;
        RECT -39.730 457.635 -37.345 457.650 ;
        RECT -39.730 457.625 -38.315 457.635 ;
        RECT -57.120 457.025 -53.725 457.195 ;
        RECT -57.120 456.975 -55.810 457.025 ;
        RECT -57.120 456.970 -56.125 456.975 ;
        RECT -57.120 455.120 -56.355 456.970 ;
        RECT -38.930 456.855 -38.315 457.625 ;
        RECT -39.740 456.840 -38.315 456.855 ;
        RECT -41.190 456.670 -38.315 456.840 ;
        RECT -39.740 456.640 -38.315 456.670 ;
        RECT -38.930 455.735 -38.315 456.640 ;
        RECT -39.815 455.700 -38.315 455.735 ;
        RECT -42.190 455.530 -38.315 455.700 ;
        RECT -57.930 454.190 -57.435 455.075 ;
        RECT -57.930 454.160 -57.360 454.190 ;
        RECT -57.190 454.175 -56.355 455.120 ;
        RECT -59.765 453.990 -57.360 454.160 ;
        RECT -57.155 453.990 -56.355 454.175 ;
        RECT -57.680 453.180 -57.360 453.990 ;
        RECT -59.765 453.010 -57.360 453.180 ;
        RECT -57.680 452.200 -57.360 453.010 ;
        RECT -59.765 452.030 -57.360 452.200 ;
        RECT -57.680 451.980 -57.360 452.030 ;
        RECT -57.120 453.690 -56.355 453.990 ;
        RECT -55.405 455.270 -54.910 455.510 ;
        RECT -39.815 455.485 -38.315 455.530 ;
        RECT -55.405 455.100 -53.580 455.270 ;
        RECT -38.930 455.105 -38.315 455.485 ;
        RECT -55.405 454.290 -54.910 455.100 ;
        RECT -39.830 455.050 -38.315 455.105 ;
        RECT -42.190 454.880 -38.315 455.050 ;
        RECT -39.830 454.855 -38.315 454.880 ;
        RECT -55.405 454.120 -53.580 454.290 ;
        RECT -55.405 453.690 -54.910 454.120 ;
        RECT -57.120 453.310 -54.910 453.690 ;
        RECT -57.120 453.140 -53.580 453.310 ;
        RECT -57.120 452.830 -54.910 453.140 ;
        RECT -57.120 451.980 -56.355 452.830 ;
        RECT -55.405 452.330 -54.910 452.830 ;
        RECT -55.405 452.160 -53.580 452.330 ;
        RECT -56.855 448.305 -56.525 451.980 ;
        RECT -55.405 451.920 -54.910 452.160 ;
        RECT -38.930 452.085 -38.315 454.855 ;
        RECT -39.715 452.075 -38.315 452.085 ;
        RECT -42.190 451.905 -38.315 452.075 ;
        RECT -39.715 451.895 -38.315 451.905 ;
        RECT -38.930 451.100 -38.315 451.895 ;
        RECT -39.725 451.095 -38.315 451.100 ;
        RECT -42.190 450.925 -38.315 451.095 ;
        RECT -39.725 450.910 -38.315 450.925 ;
        RECT -39.250 449.660 -38.665 450.910 ;
        RECT -39.885 449.075 -38.665 449.660 ;
        RECT -56.855 447.975 -49.545 448.305 ;
        RECT -56.945 446.625 -56.380 446.630 ;
        RECT -49.875 446.625 -49.545 447.975 ;
        RECT -39.885 446.750 -39.300 449.075 ;
        RECT -56.945 446.295 -49.545 446.625 ;
        RECT -56.945 446.210 -56.380 446.295 ;
        RECT -39.915 446.260 -39.285 446.750 ;
        RECT -39.855 445.120 -39.385 445.430 ;
        RECT -55.900 444.840 -55.405 445.080 ;
        RECT -57.085 444.210 -56.755 444.715 ;
        RECT -57.705 444.195 -56.755 444.210 ;
        RECT -55.900 444.670 -54.575 444.840 ;
        RECT -39.785 444.755 -39.525 445.120 ;
        RECT -38.635 444.880 -38.140 445.120 ;
        RECT -57.705 444.190 -56.200 444.195 ;
        RECT -60.665 444.020 -56.200 444.190 ;
        RECT -57.705 443.985 -56.200 444.020 ;
        RECT -57.085 442.100 -56.200 443.985 ;
        RECT -57.700 442.075 -56.200 442.100 ;
        RECT -60.665 441.905 -56.200 442.075 ;
        RECT -57.700 441.875 -56.200 441.905 ;
        RECT -57.085 441.720 -56.200 441.875 ;
        RECT -55.900 443.860 -55.405 444.670 ;
        RECT -39.820 444.250 -39.490 444.755 ;
        RECT -40.440 444.235 -39.490 444.250 ;
        RECT -38.635 444.710 -37.310 444.880 ;
        RECT -40.440 444.230 -38.935 444.235 ;
        RECT -43.400 444.060 -38.935 444.230 ;
        RECT -40.440 444.025 -38.935 444.060 ;
        RECT -55.900 443.690 -54.575 443.860 ;
        RECT -55.900 442.880 -55.405 443.690 ;
        RECT -55.900 442.710 -54.575 442.880 ;
        RECT -55.900 441.900 -55.405 442.710 ;
        RECT -39.820 442.140 -38.935 444.025 ;
        RECT -40.435 442.115 -38.935 442.140 ;
        RECT -43.400 441.945 -38.935 442.115 ;
        RECT -40.435 441.915 -38.935 441.945 ;
        RECT -55.900 441.730 -54.575 441.900 ;
        RECT -39.820 441.760 -38.935 441.915 ;
        RECT -38.635 443.900 -38.140 444.710 ;
        RECT -38.635 443.730 -37.310 443.900 ;
        RECT -38.635 442.920 -38.140 443.730 ;
        RECT -38.635 442.750 -37.310 442.920 ;
        RECT -38.635 441.940 -38.140 442.750 ;
        RECT -38.635 441.770 -37.310 441.940 ;
        RECT -57.085 441.125 -56.115 441.720 ;
        RECT -57.715 441.095 -56.115 441.125 ;
        RECT -60.665 440.925 -56.115 441.095 ;
        RECT -57.715 440.900 -56.115 440.925 ;
        RECT -57.085 440.870 -56.115 440.900 ;
        RECT -56.965 440.845 -56.115 440.870 ;
        RECT -55.900 440.845 -55.405 441.730 ;
        RECT -39.820 441.165 -38.850 441.760 ;
        RECT -40.450 441.135 -38.850 441.165 ;
        RECT -43.400 440.965 -38.850 441.135 ;
        RECT -40.450 440.940 -38.850 440.965 ;
        RECT -39.820 440.910 -38.850 440.940 ;
        RECT -56.965 440.815 -55.405 440.845 ;
        RECT -39.700 440.885 -38.850 440.910 ;
        RECT -38.635 440.885 -38.140 441.770 ;
        RECT -39.700 440.855 -38.140 440.885 ;
        RECT -56.965 440.645 -53.570 440.815 ;
        RECT -39.700 440.685 -36.305 440.855 ;
        RECT -57.775 439.845 -57.280 440.085 ;
        RECT -58.605 439.675 -57.280 439.845 ;
        RECT -57.775 438.865 -57.280 439.675 ;
        RECT -58.605 438.695 -57.280 438.865 ;
        RECT -57.775 437.885 -57.280 438.695 ;
        RECT -58.605 437.715 -57.280 437.885 ;
        RECT -57.775 436.905 -57.280 437.715 ;
        RECT -58.605 436.735 -57.280 436.905 ;
        RECT -56.965 439.835 -55.655 440.645 ;
        RECT -40.510 439.885 -40.015 440.125 ;
        RECT -56.965 439.665 -53.570 439.835 ;
        RECT -41.340 439.715 -40.015 439.885 ;
        RECT -56.965 438.855 -55.655 439.665 ;
        RECT -40.510 438.905 -40.015 439.715 ;
        RECT -56.965 438.685 -53.570 438.855 ;
        RECT -41.340 438.735 -40.015 438.905 ;
        RECT -56.965 438.635 -55.655 438.685 ;
        RECT -56.965 438.630 -55.970 438.635 ;
        RECT -56.965 436.780 -56.200 438.630 ;
        RECT -40.510 437.925 -40.015 438.735 ;
        RECT -41.340 437.755 -40.015 437.925 ;
        RECT -57.775 435.850 -57.280 436.735 ;
        RECT -57.775 435.820 -57.205 435.850 ;
        RECT -57.035 435.835 -56.200 436.780 ;
        RECT -59.610 435.650 -57.205 435.820 ;
        RECT -57.000 435.650 -56.200 435.835 ;
        RECT -57.525 434.840 -57.205 435.650 ;
        RECT -59.610 434.670 -57.205 434.840 ;
        RECT -57.525 433.860 -57.205 434.670 ;
        RECT -59.610 433.690 -57.205 433.860 ;
        RECT -57.525 433.640 -57.205 433.690 ;
        RECT -56.965 435.350 -56.200 435.650 ;
        RECT -55.250 436.930 -54.755 437.170 ;
        RECT -40.510 436.945 -40.015 437.755 ;
        RECT -55.250 436.760 -53.425 436.930 ;
        RECT -41.340 436.775 -40.015 436.945 ;
        RECT -39.700 439.875 -38.390 440.685 ;
        RECT -39.700 439.705 -36.305 439.875 ;
        RECT -39.700 438.895 -38.390 439.705 ;
        RECT -39.700 438.725 -36.305 438.895 ;
        RECT -39.700 438.675 -38.390 438.725 ;
        RECT -39.700 438.670 -38.705 438.675 ;
        RECT -39.700 436.820 -38.935 438.670 ;
        RECT -55.250 435.950 -54.755 436.760 ;
        RECT -55.250 435.780 -53.425 435.950 ;
        RECT -40.510 435.890 -40.015 436.775 ;
        RECT -40.510 435.860 -39.940 435.890 ;
        RECT -39.770 435.875 -38.935 436.820 ;
        RECT -55.250 435.350 -54.755 435.780 ;
        RECT -42.345 435.690 -39.940 435.860 ;
        RECT -39.735 435.690 -38.935 435.875 ;
        RECT -56.965 434.970 -54.755 435.350 ;
        RECT -56.965 434.800 -53.425 434.970 ;
        RECT -40.260 434.880 -39.940 435.690 ;
        RECT -56.965 434.490 -54.755 434.800 ;
        RECT -42.345 434.710 -39.940 434.880 ;
        RECT -56.965 433.640 -56.200 434.490 ;
        RECT -55.250 433.990 -54.755 434.490 ;
        RECT -55.250 433.820 -53.425 433.990 ;
        RECT -40.260 433.900 -39.940 434.710 ;
        RECT -55.250 433.580 -54.755 433.820 ;
        RECT -42.345 433.730 -39.940 433.900 ;
        RECT -40.260 433.680 -39.940 433.730 ;
        RECT -39.700 435.390 -38.935 435.690 ;
        RECT -37.985 436.970 -37.490 437.210 ;
        RECT -37.985 436.800 -36.160 436.970 ;
        RECT -37.985 435.990 -37.490 436.800 ;
        RECT -37.985 435.820 -36.160 435.990 ;
        RECT -37.985 435.390 -37.490 435.820 ;
        RECT -39.700 435.010 -37.490 435.390 ;
        RECT -39.700 434.840 -36.160 435.010 ;
        RECT -39.700 434.030 -37.490 434.840 ;
        RECT -39.700 433.860 -36.160 434.030 ;
        RECT -39.700 433.680 -37.490 433.860 ;
        RECT -39.400 433.620 -37.490 433.680 ;
        RECT -57.365 419.265 -51.080 419.630 ;
        RECT -57.505 419.020 -51.080 419.265 ;
        RECT -57.505 418.570 -56.670 419.020 ;
        RECT -57.440 417.320 -56.745 417.715 ;
        RECT -57.315 417.065 -56.900 417.320 ;
        RECT -57.410 416.820 -56.900 417.065 ;
        RECT -56.225 417.190 -55.730 417.430 ;
        RECT -56.225 417.020 -54.900 417.190 ;
        RECT -51.690 417.080 -51.080 419.020 ;
        RECT -39.400 417.080 -37.830 433.620 ;
        RECT -57.410 416.560 -57.080 416.820 ;
        RECT -58.030 416.545 -57.080 416.560 ;
        RECT -58.030 416.540 -56.525 416.545 ;
        RECT -60.990 416.370 -56.525 416.540 ;
        RECT -58.030 416.335 -56.525 416.370 ;
        RECT -57.410 414.450 -56.525 416.335 ;
        RECT -58.025 414.425 -56.525 414.450 ;
        RECT -60.990 414.255 -56.525 414.425 ;
        RECT -58.025 414.225 -56.525 414.255 ;
        RECT -57.410 414.070 -56.525 414.225 ;
        RECT -56.225 416.210 -55.730 417.020 ;
        RECT -51.690 416.470 -37.830 417.080 ;
        RECT -56.225 416.040 -54.900 416.210 ;
        RECT -56.225 415.230 -55.730 416.040 ;
        RECT -56.225 415.060 -54.900 415.230 ;
        RECT -56.225 414.250 -55.730 415.060 ;
        RECT -56.225 414.080 -54.900 414.250 ;
        RECT -57.410 413.475 -56.440 414.070 ;
        RECT -58.040 413.445 -56.440 413.475 ;
        RECT -60.990 413.275 -56.440 413.445 ;
        RECT -58.040 413.250 -56.440 413.275 ;
        RECT -57.410 413.220 -56.440 413.250 ;
        RECT -57.290 413.195 -56.440 413.220 ;
        RECT -56.225 413.195 -55.730 414.080 ;
        RECT -57.290 413.165 -55.730 413.195 ;
        RECT -57.290 412.995 -53.895 413.165 ;
        RECT -58.100 412.195 -57.605 412.435 ;
        RECT -58.930 412.025 -57.605 412.195 ;
        RECT -58.100 411.215 -57.605 412.025 ;
        RECT -58.930 411.045 -57.605 411.215 ;
        RECT -58.100 410.235 -57.605 411.045 ;
        RECT -58.930 410.065 -57.605 410.235 ;
        RECT -58.100 409.255 -57.605 410.065 ;
        RECT -58.930 409.085 -57.605 409.255 ;
        RECT -57.290 412.185 -55.980 412.995 ;
        RECT -57.290 412.015 -53.895 412.185 ;
        RECT -57.290 411.205 -55.980 412.015 ;
        RECT -39.400 411.850 -37.830 416.470 ;
        RECT -39.900 411.830 -37.830 411.850 ;
        RECT -41.360 411.720 -37.830 411.830 ;
        RECT -41.360 411.660 -38.485 411.720 ;
        RECT -39.900 411.635 -38.485 411.660 ;
        RECT -57.290 411.035 -53.895 411.205 ;
        RECT -57.290 410.985 -55.980 411.035 ;
        RECT -57.290 410.980 -56.295 410.985 ;
        RECT -57.290 409.130 -56.525 410.980 ;
        RECT -39.100 410.865 -38.485 411.635 ;
        RECT -39.910 410.850 -38.485 410.865 ;
        RECT -41.360 410.680 -38.485 410.850 ;
        RECT -39.910 410.650 -38.485 410.680 ;
        RECT -39.100 409.745 -38.485 410.650 ;
        RECT -39.985 409.710 -38.485 409.745 ;
        RECT -42.360 409.540 -38.485 409.710 ;
        RECT -58.100 408.200 -57.605 409.085 ;
        RECT -58.100 408.170 -57.530 408.200 ;
        RECT -57.360 408.185 -56.525 409.130 ;
        RECT -59.935 408.000 -57.530 408.170 ;
        RECT -57.325 408.000 -56.525 408.185 ;
        RECT -57.850 407.190 -57.530 408.000 ;
        RECT -59.935 407.020 -57.530 407.190 ;
        RECT -57.850 406.210 -57.530 407.020 ;
        RECT -59.935 406.040 -57.530 406.210 ;
        RECT -57.850 405.990 -57.530 406.040 ;
        RECT -57.290 407.700 -56.525 408.000 ;
        RECT -55.575 409.280 -55.080 409.520 ;
        RECT -39.985 409.495 -38.485 409.540 ;
        RECT -55.575 409.110 -53.750 409.280 ;
        RECT -39.100 409.115 -38.485 409.495 ;
        RECT -55.575 408.300 -55.080 409.110 ;
        RECT -40.000 409.060 -38.485 409.115 ;
        RECT -42.360 408.890 -38.485 409.060 ;
        RECT -40.000 408.865 -38.485 408.890 ;
        RECT -55.575 408.130 -53.750 408.300 ;
        RECT -55.575 407.700 -55.080 408.130 ;
        RECT -57.290 407.320 -55.080 407.700 ;
        RECT -57.290 407.150 -53.750 407.320 ;
        RECT -57.290 406.840 -55.080 407.150 ;
        RECT -57.290 405.990 -56.525 406.840 ;
        RECT -55.575 406.340 -55.080 406.840 ;
        RECT -55.575 406.170 -53.750 406.340 ;
        RECT -57.025 402.315 -56.695 405.990 ;
        RECT -55.575 405.930 -55.080 406.170 ;
        RECT -39.100 406.095 -38.485 408.865 ;
        RECT -39.885 406.085 -38.485 406.095 ;
        RECT -42.360 405.915 -38.485 406.085 ;
        RECT -39.885 405.905 -38.485 405.915 ;
        RECT -39.100 405.110 -38.485 405.905 ;
        RECT -39.895 405.105 -38.485 405.110 ;
        RECT -42.360 404.935 -38.485 405.105 ;
        RECT -39.895 404.920 -38.485 404.935 ;
        RECT -39.420 403.670 -38.835 404.920 ;
        RECT -40.055 403.085 -38.835 403.670 ;
        RECT -57.025 401.985 -49.715 402.315 ;
        RECT -57.115 400.635 -56.550 400.640 ;
        RECT -50.045 400.635 -49.715 401.985 ;
        RECT -40.055 400.760 -39.470 403.085 ;
        RECT -57.115 400.305 -49.715 400.635 ;
        RECT -57.115 400.220 -56.550 400.305 ;
        RECT -40.085 400.270 -39.455 400.760 ;
        RECT -40.025 399.130 -39.555 399.440 ;
        RECT -56.070 398.850 -55.575 399.090 ;
        RECT -57.255 398.220 -56.925 398.725 ;
        RECT -57.875 398.205 -56.925 398.220 ;
        RECT -56.070 398.680 -54.745 398.850 ;
        RECT -39.955 398.765 -39.695 399.130 ;
        RECT -38.805 398.890 -38.310 399.130 ;
        RECT -57.875 398.200 -56.370 398.205 ;
        RECT -60.835 398.030 -56.370 398.200 ;
        RECT -57.875 397.995 -56.370 398.030 ;
        RECT -57.255 396.110 -56.370 397.995 ;
        RECT -57.870 396.085 -56.370 396.110 ;
        RECT -60.835 395.915 -56.370 396.085 ;
        RECT -57.870 395.885 -56.370 395.915 ;
        RECT -57.255 395.730 -56.370 395.885 ;
        RECT -56.070 397.870 -55.575 398.680 ;
        RECT -39.990 398.260 -39.660 398.765 ;
        RECT -40.610 398.245 -39.660 398.260 ;
        RECT -38.805 398.720 -37.480 398.890 ;
        RECT -40.610 398.240 -39.105 398.245 ;
        RECT -43.570 398.070 -39.105 398.240 ;
        RECT -40.610 398.035 -39.105 398.070 ;
        RECT -56.070 397.700 -54.745 397.870 ;
        RECT -56.070 396.890 -55.575 397.700 ;
        RECT -56.070 396.720 -54.745 396.890 ;
        RECT -56.070 395.910 -55.575 396.720 ;
        RECT -39.990 396.150 -39.105 398.035 ;
        RECT -40.605 396.125 -39.105 396.150 ;
        RECT -43.570 395.955 -39.105 396.125 ;
        RECT -40.605 395.925 -39.105 395.955 ;
        RECT -56.070 395.740 -54.745 395.910 ;
        RECT -39.990 395.770 -39.105 395.925 ;
        RECT -38.805 397.910 -38.310 398.720 ;
        RECT -38.805 397.740 -37.480 397.910 ;
        RECT -38.805 396.930 -38.310 397.740 ;
        RECT -38.805 396.760 -37.480 396.930 ;
        RECT -38.805 395.950 -38.310 396.760 ;
        RECT -38.805 395.780 -37.480 395.950 ;
        RECT -57.255 395.135 -56.285 395.730 ;
        RECT -57.885 395.105 -56.285 395.135 ;
        RECT -60.835 394.935 -56.285 395.105 ;
        RECT -57.885 394.910 -56.285 394.935 ;
        RECT -57.255 394.880 -56.285 394.910 ;
        RECT -57.135 394.855 -56.285 394.880 ;
        RECT -56.070 394.855 -55.575 395.740 ;
        RECT -39.990 395.175 -39.020 395.770 ;
        RECT -40.620 395.145 -39.020 395.175 ;
        RECT -43.570 394.975 -39.020 395.145 ;
        RECT -40.620 394.950 -39.020 394.975 ;
        RECT -39.990 394.920 -39.020 394.950 ;
        RECT -57.135 394.825 -55.575 394.855 ;
        RECT -39.870 394.895 -39.020 394.920 ;
        RECT -38.805 394.895 -38.310 395.780 ;
        RECT -39.870 394.865 -38.310 394.895 ;
        RECT -57.135 394.655 -53.740 394.825 ;
        RECT -39.870 394.695 -36.475 394.865 ;
        RECT -57.945 393.855 -57.450 394.095 ;
        RECT -58.775 393.685 -57.450 393.855 ;
        RECT -57.945 392.875 -57.450 393.685 ;
        RECT -58.775 392.705 -57.450 392.875 ;
        RECT -57.945 391.895 -57.450 392.705 ;
        RECT -58.775 391.725 -57.450 391.895 ;
        RECT -57.945 390.915 -57.450 391.725 ;
        RECT -58.775 390.745 -57.450 390.915 ;
        RECT -57.135 393.845 -55.825 394.655 ;
        RECT -40.680 393.895 -40.185 394.135 ;
        RECT -57.135 393.675 -53.740 393.845 ;
        RECT -41.510 393.725 -40.185 393.895 ;
        RECT -57.135 392.865 -55.825 393.675 ;
        RECT -40.680 392.915 -40.185 393.725 ;
        RECT -57.135 392.695 -53.740 392.865 ;
        RECT -41.510 392.745 -40.185 392.915 ;
        RECT -57.135 392.645 -55.825 392.695 ;
        RECT -57.135 392.640 -56.140 392.645 ;
        RECT -57.135 390.790 -56.370 392.640 ;
        RECT -40.680 391.935 -40.185 392.745 ;
        RECT -41.510 391.765 -40.185 391.935 ;
        RECT -57.945 389.860 -57.450 390.745 ;
        RECT -57.945 389.830 -57.375 389.860 ;
        RECT -57.205 389.845 -56.370 390.790 ;
        RECT -59.780 389.660 -57.375 389.830 ;
        RECT -57.170 389.660 -56.370 389.845 ;
        RECT -57.695 388.850 -57.375 389.660 ;
        RECT -59.780 388.680 -57.375 388.850 ;
        RECT -57.695 387.870 -57.375 388.680 ;
        RECT -59.780 387.700 -57.375 387.870 ;
        RECT -57.695 387.650 -57.375 387.700 ;
        RECT -57.135 389.360 -56.370 389.660 ;
        RECT -55.420 390.940 -54.925 391.180 ;
        RECT -40.680 390.955 -40.185 391.765 ;
        RECT -55.420 390.770 -53.595 390.940 ;
        RECT -41.510 390.785 -40.185 390.955 ;
        RECT -39.870 393.885 -38.560 394.695 ;
        RECT -39.870 393.715 -36.475 393.885 ;
        RECT -39.870 392.905 -38.560 393.715 ;
        RECT -39.870 392.735 -36.475 392.905 ;
        RECT -39.870 392.685 -38.560 392.735 ;
        RECT -39.870 392.680 -38.875 392.685 ;
        RECT -39.870 390.830 -39.105 392.680 ;
        RECT -55.420 389.960 -54.925 390.770 ;
        RECT -55.420 389.790 -53.595 389.960 ;
        RECT -40.680 389.900 -40.185 390.785 ;
        RECT -40.680 389.870 -40.110 389.900 ;
        RECT -39.940 389.885 -39.105 390.830 ;
        RECT -55.420 389.360 -54.925 389.790 ;
        RECT -42.515 389.700 -40.110 389.870 ;
        RECT -39.905 389.700 -39.105 389.885 ;
        RECT -57.135 388.980 -54.925 389.360 ;
        RECT -57.135 388.810 -53.595 388.980 ;
        RECT -40.430 388.890 -40.110 389.700 ;
        RECT -57.135 388.500 -54.925 388.810 ;
        RECT -42.515 388.720 -40.110 388.890 ;
        RECT -57.135 387.650 -56.370 388.500 ;
        RECT -55.420 388.000 -54.925 388.500 ;
        RECT -55.420 387.830 -53.595 388.000 ;
        RECT -40.430 387.910 -40.110 388.720 ;
        RECT -55.420 387.590 -54.925 387.830 ;
        RECT -42.515 387.740 -40.110 387.910 ;
        RECT -40.430 387.690 -40.110 387.740 ;
        RECT -39.870 389.400 -39.105 389.700 ;
        RECT -38.155 390.980 -37.660 391.220 ;
        RECT -38.155 390.810 -36.330 390.980 ;
        RECT -38.155 390.000 -37.660 390.810 ;
        RECT -38.155 389.830 -36.330 390.000 ;
        RECT -38.155 389.400 -37.660 389.830 ;
        RECT -39.870 389.020 -37.660 389.400 ;
        RECT -39.870 388.850 -36.330 389.020 ;
        RECT -39.870 388.040 -37.660 388.850 ;
        RECT -39.870 387.870 -36.330 388.040 ;
        RECT -39.870 387.690 -37.660 387.870 ;
        RECT -39.350 387.630 -37.660 387.690 ;
        RECT -57.170 374.950 -50.885 375.315 ;
        RECT -57.310 374.705 -50.885 374.950 ;
        RECT -57.310 374.255 -56.475 374.705 ;
        RECT -57.245 373.005 -56.550 373.400 ;
        RECT -57.120 372.750 -56.705 373.005 ;
        RECT -57.215 372.505 -56.705 372.750 ;
        RECT -56.030 372.875 -55.535 373.115 ;
        RECT -56.030 372.705 -54.705 372.875 ;
        RECT -51.495 372.765 -50.885 374.705 ;
        RECT -39.350 372.765 -38.080 387.630 ;
        RECT -57.215 372.245 -56.885 372.505 ;
        RECT -57.835 372.230 -56.885 372.245 ;
        RECT -57.835 372.225 -56.330 372.230 ;
        RECT -60.795 372.055 -56.330 372.225 ;
        RECT -57.835 372.020 -56.330 372.055 ;
        RECT -57.215 370.135 -56.330 372.020 ;
        RECT -57.830 370.110 -56.330 370.135 ;
        RECT -60.795 369.940 -56.330 370.110 ;
        RECT -57.830 369.910 -56.330 369.940 ;
        RECT -57.215 369.755 -56.330 369.910 ;
        RECT -56.030 371.895 -55.535 372.705 ;
        RECT -51.495 372.155 -38.080 372.765 ;
        RECT -56.030 371.725 -54.705 371.895 ;
        RECT -56.030 370.915 -55.535 371.725 ;
        RECT -56.030 370.745 -54.705 370.915 ;
        RECT -56.030 369.935 -55.535 370.745 ;
        RECT -56.030 369.765 -54.705 369.935 ;
        RECT -57.215 369.160 -56.245 369.755 ;
        RECT -57.845 369.130 -56.245 369.160 ;
        RECT -60.795 368.960 -56.245 369.130 ;
        RECT -57.845 368.935 -56.245 368.960 ;
        RECT -57.215 368.905 -56.245 368.935 ;
        RECT -57.095 368.880 -56.245 368.905 ;
        RECT -56.030 368.880 -55.535 369.765 ;
        RECT -57.095 368.850 -55.535 368.880 ;
        RECT -57.095 368.680 -53.700 368.850 ;
        RECT -57.905 367.880 -57.410 368.120 ;
        RECT -58.735 367.710 -57.410 367.880 ;
        RECT -57.905 366.900 -57.410 367.710 ;
        RECT -58.735 366.730 -57.410 366.900 ;
        RECT -57.905 365.920 -57.410 366.730 ;
        RECT -58.735 365.750 -57.410 365.920 ;
        RECT -57.905 364.940 -57.410 365.750 ;
        RECT -58.735 364.770 -57.410 364.940 ;
        RECT -57.095 367.870 -55.785 368.680 ;
        RECT -57.095 367.700 -53.700 367.870 ;
        RECT -57.095 366.890 -55.785 367.700 ;
        RECT -39.350 367.535 -38.080 372.155 ;
        RECT -39.705 367.515 -38.080 367.535 ;
        RECT -41.165 367.465 -38.080 367.515 ;
        RECT -41.165 367.345 -38.290 367.465 ;
        RECT -39.705 367.320 -38.290 367.345 ;
        RECT -57.095 366.720 -53.700 366.890 ;
        RECT -57.095 366.670 -55.785 366.720 ;
        RECT -57.095 366.665 -56.100 366.670 ;
        RECT -57.095 364.815 -56.330 366.665 ;
        RECT -38.905 366.550 -38.290 367.320 ;
        RECT -39.715 366.535 -38.290 366.550 ;
        RECT -41.165 366.365 -38.290 366.535 ;
        RECT -39.715 366.335 -38.290 366.365 ;
        RECT -38.905 365.430 -38.290 366.335 ;
        RECT -39.790 365.395 -38.290 365.430 ;
        RECT -42.165 365.225 -38.290 365.395 ;
        RECT -57.905 363.885 -57.410 364.770 ;
        RECT -57.905 363.855 -57.335 363.885 ;
        RECT -57.165 363.870 -56.330 364.815 ;
        RECT -59.740 363.685 -57.335 363.855 ;
        RECT -57.130 363.685 -56.330 363.870 ;
        RECT -57.655 362.875 -57.335 363.685 ;
        RECT -59.740 362.705 -57.335 362.875 ;
        RECT -57.655 361.895 -57.335 362.705 ;
        RECT -59.740 361.725 -57.335 361.895 ;
        RECT -57.655 361.675 -57.335 361.725 ;
        RECT -57.095 363.385 -56.330 363.685 ;
        RECT -55.380 364.965 -54.885 365.205 ;
        RECT -39.790 365.180 -38.290 365.225 ;
        RECT -55.380 364.795 -53.555 364.965 ;
        RECT -38.905 364.800 -38.290 365.180 ;
        RECT -55.380 363.985 -54.885 364.795 ;
        RECT -39.805 364.745 -38.290 364.800 ;
        RECT -42.165 364.575 -38.290 364.745 ;
        RECT -39.805 364.550 -38.290 364.575 ;
        RECT -55.380 363.815 -53.555 363.985 ;
        RECT -55.380 363.385 -54.885 363.815 ;
        RECT -57.095 363.005 -54.885 363.385 ;
        RECT -57.095 362.835 -53.555 363.005 ;
        RECT -57.095 362.525 -54.885 362.835 ;
        RECT -57.095 361.675 -56.330 362.525 ;
        RECT -55.380 362.025 -54.885 362.525 ;
        RECT -55.380 361.855 -53.555 362.025 ;
        RECT -56.830 358.000 -56.500 361.675 ;
        RECT -55.380 361.615 -54.885 361.855 ;
        RECT -38.905 361.780 -38.290 364.550 ;
        RECT -39.690 361.770 -38.290 361.780 ;
        RECT -42.165 361.600 -38.290 361.770 ;
        RECT -39.690 361.590 -38.290 361.600 ;
        RECT -38.905 360.795 -38.290 361.590 ;
        RECT -39.700 360.790 -38.290 360.795 ;
        RECT -42.165 360.620 -38.290 360.790 ;
        RECT -39.700 360.605 -38.290 360.620 ;
        RECT -39.225 359.355 -38.640 360.605 ;
        RECT -39.860 358.770 -38.640 359.355 ;
        RECT -56.830 357.670 -49.520 358.000 ;
        RECT -56.920 356.320 -56.355 356.325 ;
        RECT -49.850 356.320 -49.520 357.670 ;
        RECT -39.860 356.445 -39.275 358.770 ;
        RECT -56.920 355.990 -49.520 356.320 ;
        RECT -56.920 355.905 -56.355 355.990 ;
        RECT -39.890 355.955 -39.260 356.445 ;
        RECT -39.830 354.815 -39.360 355.125 ;
        RECT -55.875 354.535 -55.380 354.775 ;
        RECT -57.060 353.905 -56.730 354.410 ;
        RECT -57.680 353.890 -56.730 353.905 ;
        RECT -55.875 354.365 -54.550 354.535 ;
        RECT -39.760 354.450 -39.500 354.815 ;
        RECT -38.610 354.575 -38.115 354.815 ;
        RECT -57.680 353.885 -56.175 353.890 ;
        RECT -60.640 353.715 -56.175 353.885 ;
        RECT -57.680 353.680 -56.175 353.715 ;
        RECT -57.060 351.795 -56.175 353.680 ;
        RECT -57.675 351.770 -56.175 351.795 ;
        RECT -60.640 351.600 -56.175 351.770 ;
        RECT -57.675 351.570 -56.175 351.600 ;
        RECT -57.060 351.415 -56.175 351.570 ;
        RECT -55.875 353.555 -55.380 354.365 ;
        RECT -39.795 353.945 -39.465 354.450 ;
        RECT -40.415 353.930 -39.465 353.945 ;
        RECT -38.610 354.405 -37.285 354.575 ;
        RECT -40.415 353.925 -38.910 353.930 ;
        RECT -43.375 353.755 -38.910 353.925 ;
        RECT -40.415 353.720 -38.910 353.755 ;
        RECT -55.875 353.385 -54.550 353.555 ;
        RECT -55.875 352.575 -55.380 353.385 ;
        RECT -55.875 352.405 -54.550 352.575 ;
        RECT -55.875 351.595 -55.380 352.405 ;
        RECT -39.795 351.835 -38.910 353.720 ;
        RECT -40.410 351.810 -38.910 351.835 ;
        RECT -43.375 351.640 -38.910 351.810 ;
        RECT -40.410 351.610 -38.910 351.640 ;
        RECT -55.875 351.425 -54.550 351.595 ;
        RECT -39.795 351.455 -38.910 351.610 ;
        RECT -38.610 353.595 -38.115 354.405 ;
        RECT -38.610 353.425 -37.285 353.595 ;
        RECT -38.610 352.615 -38.115 353.425 ;
        RECT -38.610 352.445 -37.285 352.615 ;
        RECT -38.610 351.635 -38.115 352.445 ;
        RECT -38.610 351.465 -37.285 351.635 ;
        RECT -57.060 350.820 -56.090 351.415 ;
        RECT -57.690 350.790 -56.090 350.820 ;
        RECT -60.640 350.620 -56.090 350.790 ;
        RECT -57.690 350.595 -56.090 350.620 ;
        RECT -57.060 350.565 -56.090 350.595 ;
        RECT -56.940 350.540 -56.090 350.565 ;
        RECT -55.875 350.540 -55.380 351.425 ;
        RECT -39.795 350.860 -38.825 351.455 ;
        RECT -40.425 350.830 -38.825 350.860 ;
        RECT -43.375 350.660 -38.825 350.830 ;
        RECT -40.425 350.635 -38.825 350.660 ;
        RECT -39.795 350.605 -38.825 350.635 ;
        RECT -56.940 350.510 -55.380 350.540 ;
        RECT -39.675 350.580 -38.825 350.605 ;
        RECT -38.610 350.580 -38.115 351.465 ;
        RECT -39.675 350.550 -38.115 350.580 ;
        RECT -56.940 350.340 -53.545 350.510 ;
        RECT -39.675 350.380 -36.280 350.550 ;
        RECT -57.750 349.540 -57.255 349.780 ;
        RECT -58.580 349.370 -57.255 349.540 ;
        RECT -57.750 348.560 -57.255 349.370 ;
        RECT -58.580 348.390 -57.255 348.560 ;
        RECT -57.750 347.580 -57.255 348.390 ;
        RECT -58.580 347.410 -57.255 347.580 ;
        RECT -57.750 346.600 -57.255 347.410 ;
        RECT -58.580 346.430 -57.255 346.600 ;
        RECT -56.940 349.530 -55.630 350.340 ;
        RECT -40.485 349.580 -39.990 349.820 ;
        RECT -56.940 349.360 -53.545 349.530 ;
        RECT -41.315 349.410 -39.990 349.580 ;
        RECT -56.940 348.550 -55.630 349.360 ;
        RECT -40.485 348.600 -39.990 349.410 ;
        RECT -56.940 348.380 -53.545 348.550 ;
        RECT -41.315 348.430 -39.990 348.600 ;
        RECT -56.940 348.330 -55.630 348.380 ;
        RECT -56.940 348.325 -55.945 348.330 ;
        RECT -56.940 346.475 -56.175 348.325 ;
        RECT -40.485 347.620 -39.990 348.430 ;
        RECT -41.315 347.450 -39.990 347.620 ;
        RECT -57.750 345.545 -57.255 346.430 ;
        RECT -57.750 345.515 -57.180 345.545 ;
        RECT -57.010 345.530 -56.175 346.475 ;
        RECT -59.585 345.345 -57.180 345.515 ;
        RECT -56.975 345.345 -56.175 345.530 ;
        RECT -57.500 344.535 -57.180 345.345 ;
        RECT -59.585 344.365 -57.180 344.535 ;
        RECT -57.500 343.555 -57.180 344.365 ;
        RECT -59.585 343.385 -57.180 343.555 ;
        RECT -57.500 343.335 -57.180 343.385 ;
        RECT -56.940 345.045 -56.175 345.345 ;
        RECT -55.225 346.625 -54.730 346.865 ;
        RECT -40.485 346.640 -39.990 347.450 ;
        RECT -55.225 346.455 -53.400 346.625 ;
        RECT -41.315 346.470 -39.990 346.640 ;
        RECT -39.675 349.570 -38.365 350.380 ;
        RECT -39.675 349.400 -36.280 349.570 ;
        RECT -39.675 348.590 -38.365 349.400 ;
        RECT -39.675 348.420 -36.280 348.590 ;
        RECT -39.675 348.370 -38.365 348.420 ;
        RECT -39.675 348.365 -38.680 348.370 ;
        RECT -39.675 346.515 -38.910 348.365 ;
        RECT -55.225 345.645 -54.730 346.455 ;
        RECT -55.225 345.475 -53.400 345.645 ;
        RECT -40.485 345.585 -39.990 346.470 ;
        RECT -40.485 345.555 -39.915 345.585 ;
        RECT -39.745 345.570 -38.910 346.515 ;
        RECT -55.225 345.045 -54.730 345.475 ;
        RECT -42.320 345.385 -39.915 345.555 ;
        RECT -39.710 345.385 -38.910 345.570 ;
        RECT -56.940 344.665 -54.730 345.045 ;
        RECT -56.940 344.495 -53.400 344.665 ;
        RECT -40.235 344.575 -39.915 345.385 ;
        RECT -56.940 344.185 -54.730 344.495 ;
        RECT -42.320 344.405 -39.915 344.575 ;
        RECT -56.940 343.335 -56.175 344.185 ;
        RECT -55.225 343.685 -54.730 344.185 ;
        RECT -55.225 343.515 -53.400 343.685 ;
        RECT -40.235 343.595 -39.915 344.405 ;
        RECT -55.225 343.275 -54.730 343.515 ;
        RECT -42.320 343.425 -39.915 343.595 ;
        RECT -40.235 343.375 -39.915 343.425 ;
        RECT -39.675 345.085 -38.910 345.385 ;
        RECT -37.960 346.665 -37.465 346.905 ;
        RECT -37.960 346.495 -36.135 346.665 ;
        RECT -37.960 345.685 -37.465 346.495 ;
        RECT -37.960 345.515 -36.135 345.685 ;
        RECT -37.960 345.085 -37.465 345.515 ;
        RECT -39.675 344.705 -37.465 345.085 ;
        RECT -39.675 344.535 -36.135 344.705 ;
        RECT -39.675 344.225 -37.465 344.535 ;
        RECT -57.115 332.750 -50.830 333.115 ;
        RECT -57.255 332.505 -50.830 332.750 ;
        RECT -57.255 332.055 -56.420 332.505 ;
        RECT -57.190 330.805 -56.495 331.200 ;
        RECT -57.065 330.550 -56.650 330.805 ;
        RECT -57.160 330.305 -56.650 330.550 ;
        RECT -55.975 330.675 -55.480 330.915 ;
        RECT -55.975 330.505 -54.650 330.675 ;
        RECT -51.440 330.565 -50.830 332.505 ;
        RECT -39.675 330.565 -38.910 344.225 ;
        RECT -37.960 343.725 -37.465 344.225 ;
        RECT -37.960 343.555 -36.135 343.725 ;
        RECT -37.960 343.315 -37.465 343.555 ;
        RECT -57.160 330.045 -56.830 330.305 ;
        RECT -57.780 330.030 -56.830 330.045 ;
        RECT -57.780 330.025 -56.275 330.030 ;
        RECT -60.740 329.855 -56.275 330.025 ;
        RECT -57.780 329.820 -56.275 329.855 ;
        RECT -57.160 327.935 -56.275 329.820 ;
        RECT -57.775 327.910 -56.275 327.935 ;
        RECT -60.740 327.740 -56.275 327.910 ;
        RECT -57.775 327.710 -56.275 327.740 ;
        RECT -57.160 327.555 -56.275 327.710 ;
        RECT -55.975 329.695 -55.480 330.505 ;
        RECT -51.440 329.955 -38.235 330.565 ;
        RECT -55.975 329.525 -54.650 329.695 ;
        RECT -55.975 328.715 -55.480 329.525 ;
        RECT -55.975 328.545 -54.650 328.715 ;
        RECT -55.975 327.735 -55.480 328.545 ;
        RECT -55.975 327.565 -54.650 327.735 ;
        RECT -57.160 326.960 -56.190 327.555 ;
        RECT -57.790 326.930 -56.190 326.960 ;
        RECT -60.740 326.760 -56.190 326.930 ;
        RECT -57.790 326.735 -56.190 326.760 ;
        RECT -57.160 326.705 -56.190 326.735 ;
        RECT -57.040 326.680 -56.190 326.705 ;
        RECT -55.975 326.680 -55.480 327.565 ;
        RECT -57.040 326.650 -55.480 326.680 ;
        RECT -57.040 326.480 -53.645 326.650 ;
        RECT -57.850 325.680 -57.355 325.920 ;
        RECT -58.680 325.510 -57.355 325.680 ;
        RECT -57.850 324.700 -57.355 325.510 ;
        RECT -58.680 324.530 -57.355 324.700 ;
        RECT -57.850 323.720 -57.355 324.530 ;
        RECT -58.680 323.550 -57.355 323.720 ;
        RECT -57.850 322.740 -57.355 323.550 ;
        RECT -58.680 322.570 -57.355 322.740 ;
        RECT -57.040 325.670 -55.730 326.480 ;
        RECT -57.040 325.500 -53.645 325.670 ;
        RECT -57.040 324.690 -55.730 325.500 ;
        RECT -38.845 325.335 -38.235 329.955 ;
        RECT -39.650 325.315 -38.235 325.335 ;
        RECT -41.110 325.145 -38.235 325.315 ;
        RECT -39.650 325.120 -38.235 325.145 ;
        RECT -57.040 324.520 -53.645 324.690 ;
        RECT -57.040 324.470 -55.730 324.520 ;
        RECT -57.040 324.465 -56.045 324.470 ;
        RECT -57.040 322.615 -56.275 324.465 ;
        RECT -38.850 324.350 -38.235 325.120 ;
        RECT -39.660 324.335 -38.235 324.350 ;
        RECT -41.110 324.165 -38.235 324.335 ;
        RECT -39.660 324.135 -38.235 324.165 ;
        RECT -38.850 323.230 -38.235 324.135 ;
        RECT -39.735 323.195 -38.235 323.230 ;
        RECT -42.110 323.025 -38.235 323.195 ;
        RECT -57.850 321.685 -57.355 322.570 ;
        RECT -57.850 321.655 -57.280 321.685 ;
        RECT -57.110 321.670 -56.275 322.615 ;
        RECT -59.685 321.485 -57.280 321.655 ;
        RECT -57.075 321.485 -56.275 321.670 ;
        RECT -57.600 320.675 -57.280 321.485 ;
        RECT -59.685 320.505 -57.280 320.675 ;
        RECT -57.600 319.695 -57.280 320.505 ;
        RECT -59.685 319.525 -57.280 319.695 ;
        RECT -57.600 319.475 -57.280 319.525 ;
        RECT -57.040 321.185 -56.275 321.485 ;
        RECT -55.325 322.765 -54.830 323.005 ;
        RECT -39.735 322.980 -38.235 323.025 ;
        RECT -55.325 322.595 -53.500 322.765 ;
        RECT -38.850 322.600 -38.235 322.980 ;
        RECT -55.325 321.785 -54.830 322.595 ;
        RECT -39.750 322.545 -38.235 322.600 ;
        RECT -42.110 322.375 -38.235 322.545 ;
        RECT -39.750 322.350 -38.235 322.375 ;
        RECT -55.325 321.615 -53.500 321.785 ;
        RECT -55.325 321.185 -54.830 321.615 ;
        RECT -57.040 320.805 -54.830 321.185 ;
        RECT -57.040 320.635 -53.500 320.805 ;
        RECT -57.040 320.325 -54.830 320.635 ;
        RECT -57.040 319.475 -56.275 320.325 ;
        RECT -55.325 319.825 -54.830 320.325 ;
        RECT -55.325 319.655 -53.500 319.825 ;
        RECT -56.775 315.800 -56.445 319.475 ;
        RECT -55.325 319.415 -54.830 319.655 ;
        RECT -38.850 319.580 -38.235 322.350 ;
        RECT -39.635 319.570 -38.235 319.580 ;
        RECT -42.110 319.400 -38.235 319.570 ;
        RECT -39.635 319.390 -38.235 319.400 ;
        RECT -38.850 318.595 -38.235 319.390 ;
        RECT -39.645 318.590 -38.235 318.595 ;
        RECT -42.110 318.420 -38.235 318.590 ;
        RECT -39.645 318.405 -38.235 318.420 ;
        RECT -39.170 317.155 -38.585 318.405 ;
        RECT -39.805 316.570 -38.585 317.155 ;
        RECT -56.775 315.470 -49.465 315.800 ;
        RECT -56.865 314.120 -56.300 314.125 ;
        RECT -49.795 314.120 -49.465 315.470 ;
        RECT -39.805 314.245 -39.220 316.570 ;
        RECT -56.865 313.790 -49.465 314.120 ;
        RECT -56.865 313.705 -56.300 313.790 ;
        RECT -39.835 313.755 -39.205 314.245 ;
        RECT -39.775 312.615 -39.305 312.925 ;
        RECT -55.820 312.335 -55.325 312.575 ;
        RECT -57.005 311.705 -56.675 312.210 ;
        RECT -57.625 311.690 -56.675 311.705 ;
        RECT -55.820 312.165 -54.495 312.335 ;
        RECT -39.705 312.250 -39.445 312.615 ;
        RECT -38.555 312.375 -38.060 312.615 ;
        RECT -57.625 311.685 -56.120 311.690 ;
        RECT -60.585 311.515 -56.120 311.685 ;
        RECT -57.625 311.480 -56.120 311.515 ;
        RECT -57.005 309.595 -56.120 311.480 ;
        RECT -57.620 309.570 -56.120 309.595 ;
        RECT -60.585 309.400 -56.120 309.570 ;
        RECT -57.620 309.370 -56.120 309.400 ;
        RECT -57.005 309.215 -56.120 309.370 ;
        RECT -55.820 311.355 -55.325 312.165 ;
        RECT -39.740 311.745 -39.410 312.250 ;
        RECT -40.360 311.730 -39.410 311.745 ;
        RECT -38.555 312.205 -37.230 312.375 ;
        RECT -40.360 311.725 -38.855 311.730 ;
        RECT -43.320 311.555 -38.855 311.725 ;
        RECT -40.360 311.520 -38.855 311.555 ;
        RECT -55.820 311.185 -54.495 311.355 ;
        RECT -55.820 310.375 -55.325 311.185 ;
        RECT -55.820 310.205 -54.495 310.375 ;
        RECT -55.820 309.395 -55.325 310.205 ;
        RECT -39.740 309.635 -38.855 311.520 ;
        RECT -40.355 309.610 -38.855 309.635 ;
        RECT -43.320 309.440 -38.855 309.610 ;
        RECT -40.355 309.410 -38.855 309.440 ;
        RECT -55.820 309.225 -54.495 309.395 ;
        RECT -39.740 309.255 -38.855 309.410 ;
        RECT -38.555 311.395 -38.060 312.205 ;
        RECT -38.555 311.225 -37.230 311.395 ;
        RECT -38.555 310.415 -38.060 311.225 ;
        RECT -38.555 310.245 -37.230 310.415 ;
        RECT -38.555 309.435 -38.060 310.245 ;
        RECT -38.555 309.265 -37.230 309.435 ;
        RECT -57.005 308.620 -56.035 309.215 ;
        RECT -57.635 308.590 -56.035 308.620 ;
        RECT -60.585 308.420 -56.035 308.590 ;
        RECT -57.635 308.395 -56.035 308.420 ;
        RECT -57.005 308.365 -56.035 308.395 ;
        RECT -56.885 308.340 -56.035 308.365 ;
        RECT -55.820 308.340 -55.325 309.225 ;
        RECT -39.740 308.660 -38.770 309.255 ;
        RECT -40.370 308.630 -38.770 308.660 ;
        RECT -43.320 308.460 -38.770 308.630 ;
        RECT -40.370 308.435 -38.770 308.460 ;
        RECT -39.740 308.405 -38.770 308.435 ;
        RECT -56.885 308.310 -55.325 308.340 ;
        RECT -39.620 308.380 -38.770 308.405 ;
        RECT -38.555 308.380 -38.060 309.265 ;
        RECT -39.620 308.350 -38.060 308.380 ;
        RECT -56.885 308.140 -53.490 308.310 ;
        RECT -39.620 308.180 -36.225 308.350 ;
        RECT -57.695 307.340 -57.200 307.580 ;
        RECT -58.525 307.170 -57.200 307.340 ;
        RECT -57.695 306.360 -57.200 307.170 ;
        RECT -58.525 306.190 -57.200 306.360 ;
        RECT -57.695 305.380 -57.200 306.190 ;
        RECT -58.525 305.210 -57.200 305.380 ;
        RECT -57.695 304.400 -57.200 305.210 ;
        RECT -58.525 304.230 -57.200 304.400 ;
        RECT -56.885 307.330 -55.575 308.140 ;
        RECT -40.430 307.380 -39.935 307.620 ;
        RECT -56.885 307.160 -53.490 307.330 ;
        RECT -41.260 307.210 -39.935 307.380 ;
        RECT -56.885 306.350 -55.575 307.160 ;
        RECT -40.430 306.400 -39.935 307.210 ;
        RECT -56.885 306.180 -53.490 306.350 ;
        RECT -41.260 306.230 -39.935 306.400 ;
        RECT -56.885 306.130 -55.575 306.180 ;
        RECT -56.885 306.125 -55.890 306.130 ;
        RECT -56.885 304.275 -56.120 306.125 ;
        RECT -40.430 305.420 -39.935 306.230 ;
        RECT -41.260 305.250 -39.935 305.420 ;
        RECT -57.695 303.345 -57.200 304.230 ;
        RECT -57.695 303.315 -57.125 303.345 ;
        RECT -56.955 303.330 -56.120 304.275 ;
        RECT -59.530 303.145 -57.125 303.315 ;
        RECT -56.920 303.145 -56.120 303.330 ;
        RECT -57.445 302.335 -57.125 303.145 ;
        RECT -59.530 302.165 -57.125 302.335 ;
        RECT -57.445 301.355 -57.125 302.165 ;
        RECT -59.530 301.185 -57.125 301.355 ;
        RECT -57.445 301.135 -57.125 301.185 ;
        RECT -56.885 302.845 -56.120 303.145 ;
        RECT -55.170 304.425 -54.675 304.665 ;
        RECT -40.430 304.440 -39.935 305.250 ;
        RECT -55.170 304.255 -53.345 304.425 ;
        RECT -41.260 304.270 -39.935 304.440 ;
        RECT -39.620 307.370 -38.310 308.180 ;
        RECT -39.620 307.200 -36.225 307.370 ;
        RECT -39.620 306.390 -38.310 307.200 ;
        RECT -39.620 306.220 -36.225 306.390 ;
        RECT -39.620 306.170 -38.310 306.220 ;
        RECT -39.620 306.165 -38.625 306.170 ;
        RECT -39.620 304.315 -38.855 306.165 ;
        RECT -55.170 303.445 -54.675 304.255 ;
        RECT -55.170 303.275 -53.345 303.445 ;
        RECT -40.430 303.385 -39.935 304.270 ;
        RECT -40.430 303.355 -39.860 303.385 ;
        RECT -39.690 303.370 -38.855 304.315 ;
        RECT -55.170 302.845 -54.675 303.275 ;
        RECT -42.265 303.185 -39.860 303.355 ;
        RECT -39.655 303.185 -38.855 303.370 ;
        RECT -56.885 302.465 -54.675 302.845 ;
        RECT -56.885 302.295 -53.345 302.465 ;
        RECT -40.180 302.375 -39.860 303.185 ;
        RECT -56.885 301.985 -54.675 302.295 ;
        RECT -42.265 302.205 -39.860 302.375 ;
        RECT -56.885 301.135 -56.120 301.985 ;
        RECT -55.170 301.485 -54.675 301.985 ;
        RECT -55.170 301.315 -53.345 301.485 ;
        RECT -40.180 301.395 -39.860 302.205 ;
        RECT -55.170 301.075 -54.675 301.315 ;
        RECT -42.265 301.225 -39.860 301.395 ;
        RECT -40.180 301.175 -39.860 301.225 ;
        RECT -39.620 302.885 -38.855 303.185 ;
        RECT -37.905 304.465 -37.410 304.705 ;
        RECT -37.905 304.295 -36.080 304.465 ;
        RECT -37.905 303.485 -37.410 304.295 ;
        RECT -37.905 303.315 -36.080 303.485 ;
        RECT -37.905 302.885 -37.410 303.315 ;
        RECT -39.620 302.505 -37.410 302.885 ;
        RECT -39.620 302.335 -36.080 302.505 ;
        RECT -39.620 301.525 -37.410 302.335 ;
        RECT -39.620 301.355 -36.080 301.525 ;
        RECT -39.620 301.175 -37.410 301.355 ;
        RECT -39.200 301.115 -37.410 301.175 ;
        RECT -39.200 290.555 -37.730 301.115 ;
        RECT -18.150 298.205 -12.635 596.055 ;
        RECT -25.095 292.690 -12.635 298.205 ;
        RECT -57.535 290.110 -37.090 290.555 ;
        RECT -57.535 289.590 -57.020 290.110 ;
        RECT -57.535 289.420 -52.845 289.590 ;
        RECT -57.535 288.610 -57.020 289.420 ;
        RECT -46.245 289.120 -45.905 290.110 ;
        RECT -37.430 289.310 -37.090 290.110 ;
        RECT -38.885 289.140 -37.090 289.310 ;
        RECT -46.245 288.820 -45.890 289.120 ;
        RECT -46.245 288.650 -44.435 288.820 ;
        RECT -57.535 288.440 -52.845 288.610 ;
        RECT -57.535 287.590 -57.020 288.440 ;
        RECT -46.245 287.840 -45.890 288.650 ;
        RECT -37.430 288.330 -37.090 289.140 ;
        RECT -38.885 288.160 -37.090 288.330 ;
        RECT -46.245 287.670 -44.435 287.840 ;
        RECT -57.535 287.420 -52.845 287.590 ;
        RECT -57.535 286.610 -57.020 287.420 ;
        RECT -46.245 286.860 -45.890 287.670 ;
        RECT -37.430 287.350 -37.090 288.160 ;
        RECT -38.885 287.180 -37.090 287.350 ;
        RECT -46.245 286.690 -44.435 286.860 ;
        RECT -46.245 286.645 -45.890 286.690 ;
        RECT -57.535 286.440 -52.845 286.610 ;
        RECT -57.535 284.590 -57.020 286.440 ;
        RECT -46.245 285.035 -45.905 286.645 ;
        RECT -37.430 285.125 -37.090 287.180 ;
        RECT -57.535 284.420 -52.845 284.590 ;
        RECT -57.535 283.610 -57.020 284.420 ;
        RECT -57.535 283.440 -52.845 283.610 ;
        RECT -57.535 282.590 -57.020 283.440 ;
        RECT -57.535 282.420 -52.845 282.590 ;
        RECT -57.535 281.610 -57.020 282.420 ;
        RECT -57.535 281.440 -52.845 281.610 ;
        RECT -57.535 279.590 -57.020 281.440 ;
        RECT -46.230 280.410 -45.915 285.035 ;
        RECT -38.885 284.955 -37.090 285.125 ;
        RECT -37.430 284.145 -37.090 284.955 ;
        RECT -38.885 283.975 -37.090 284.145 ;
        RECT -37.430 283.165 -37.090 283.975 ;
        RECT -38.885 282.995 -37.090 283.165 ;
        RECT -37.430 282.690 -37.090 282.995 ;
        RECT -46.230 280.105 -45.890 280.410 ;
        RECT -46.230 279.935 -44.435 280.105 ;
        RECT -57.535 279.420 -52.845 279.590 ;
        RECT -57.535 278.610 -57.020 279.420 ;
        RECT -46.230 279.125 -45.890 279.935 ;
        RECT -46.230 278.955 -44.435 279.125 ;
        RECT -57.535 278.440 -52.845 278.610 ;
        RECT -57.535 277.590 -57.020 278.440 ;
        RECT -46.230 278.145 -45.890 278.955 ;
        RECT -37.405 278.200 -37.090 282.690 ;
        RECT -46.230 277.975 -44.435 278.145 ;
        RECT -57.535 277.420 -52.845 277.590 ;
        RECT -57.535 276.610 -57.020 277.420 ;
        RECT -57.535 276.440 -52.845 276.610 ;
        RECT -57.535 274.170 -57.020 276.440 ;
        RECT -46.230 275.320 -45.890 277.975 ;
        RECT -37.430 275.810 -37.090 278.200 ;
        RECT -38.885 275.640 -37.090 275.810 ;
        RECT -46.230 275.150 -44.435 275.320 ;
        RECT -47.650 274.420 -47.330 274.450 ;
        RECT -50.235 274.250 -47.330 274.420 ;
        RECT -57.535 274.110 -55.700 274.170 ;
        RECT -57.495 274.000 -55.700 274.110 ;
        RECT -57.495 273.190 -57.155 274.000 ;
        RECT -47.650 273.690 -47.330 274.250 ;
        RECT -46.230 274.340 -45.890 275.150 ;
        RECT -37.430 274.830 -37.090 275.640 ;
        RECT -38.885 274.660 -37.090 274.830 ;
        RECT -46.230 274.170 -44.435 274.340 ;
        RECT -46.230 273.945 -45.890 274.170 ;
        RECT -46.235 273.690 -45.890 273.945 ;
        RECT -37.430 273.850 -37.090 274.660 ;
        RECT -47.650 273.440 -45.890 273.690 ;
        RECT -38.885 273.680 -37.090 273.850 ;
        RECT -50.235 273.360 -45.890 273.440 ;
        RECT -50.235 273.270 -44.435 273.360 ;
        RECT -47.650 273.190 -44.435 273.270 ;
        RECT -57.495 273.020 -55.700 273.190 ;
        RECT -47.650 273.145 -45.890 273.190 ;
        RECT -57.495 272.210 -57.155 273.020 ;
        RECT -47.650 272.530 -45.895 273.145 ;
        RECT -47.650 272.460 -47.330 272.530 ;
        RECT -50.235 272.290 -47.330 272.460 ;
        RECT -47.650 272.240 -47.330 272.290 ;
        RECT -57.495 272.040 -55.700 272.210 ;
        RECT -57.495 270.895 -57.155 272.040 ;
        RECT -46.235 271.580 -45.895 272.530 ;
        RECT -37.430 271.625 -37.090 273.680 ;
        RECT -57.560 270.525 -57.125 270.895 ;
        RECT -57.530 269.545 -57.195 270.525 ;
        RECT -57.530 269.375 -55.735 269.545 ;
        RECT -57.530 268.565 -57.195 269.375 ;
        RECT -57.530 268.395 -55.735 268.565 ;
        RECT -57.530 267.435 -57.195 268.395 ;
        RECT -57.615 267.120 -57.125 267.435 ;
        RECT -57.560 265.855 -57.215 267.120 ;
        RECT -46.230 266.910 -45.915 271.580 ;
        RECT -38.885 271.455 -37.090 271.625 ;
        RECT -37.430 270.645 -37.090 271.455 ;
        RECT -38.885 270.475 -37.090 270.645 ;
        RECT -37.430 269.665 -37.090 270.475 ;
        RECT -38.885 269.495 -37.090 269.665 ;
        RECT -37.430 269.190 -37.090 269.495 ;
        RECT -46.230 266.605 -45.890 266.910 ;
        RECT -46.230 266.435 -44.435 266.605 ;
        RECT -57.560 265.685 -55.735 265.855 ;
        RECT -57.560 264.875 -57.215 265.685 ;
        RECT -46.230 265.625 -45.890 266.435 ;
        RECT -46.230 265.455 -44.435 265.625 ;
        RECT -57.560 264.705 -55.735 264.875 ;
        RECT -57.560 263.895 -57.215 264.705 ;
        RECT -46.230 264.645 -45.890 265.455 ;
        RECT -46.230 264.475 -44.435 264.645 ;
        RECT -57.560 263.725 -55.735 263.895 ;
        RECT -57.560 262.915 -57.215 263.725 ;
        RECT -57.560 262.745 -55.735 262.915 ;
        RECT -57.560 261.950 -57.215 262.745 ;
        RECT -46.230 262.195 -45.890 264.475 ;
        RECT -37.405 264.430 -37.090 269.190 ;
        RECT -46.230 262.025 -44.435 262.195 ;
        RECT -57.580 261.520 -57.115 261.950 ;
        RECT -57.500 259.355 -57.155 261.520 ;
        RECT -46.230 261.215 -45.890 262.025 ;
        RECT -46.230 261.045 -44.435 261.215 ;
        RECT -46.230 260.235 -45.890 261.045 ;
        RECT -46.230 260.065 -44.435 260.235 ;
        RECT -46.230 260.020 -45.890 260.065 ;
        RECT -57.500 259.315 -56.490 259.355 ;
        RECT -57.500 259.145 -54.565 259.315 ;
        RECT -57.500 259.115 -56.490 259.145 ;
        RECT -57.500 258.370 -57.155 259.115 ;
        RECT -57.500 258.335 -56.520 258.370 ;
        RECT -57.500 258.165 -54.565 258.335 ;
        RECT -57.500 258.130 -56.520 258.165 ;
        RECT -57.500 254.625 -57.155 258.130 ;
        RECT -46.060 254.660 -45.395 257.755 ;
        RECT -57.500 254.585 -56.490 254.625 ;
        RECT -46.060 254.610 -44.755 254.660 ;
        RECT -57.500 254.415 -54.565 254.585 ;
        RECT -46.060 254.440 -41.835 254.610 ;
        RECT -57.500 254.385 -56.490 254.415 ;
        RECT -46.060 254.395 -44.755 254.440 ;
        RECT -57.500 253.640 -57.155 254.385 ;
        RECT -46.060 253.680 -45.395 254.395 ;
        RECT -57.500 253.605 -56.520 253.640 ;
        RECT -46.060 253.630 -44.835 253.680 ;
        RECT -57.500 253.435 -54.565 253.605 ;
        RECT -46.060 253.460 -41.835 253.630 ;
        RECT -57.500 253.400 -56.520 253.435 ;
        RECT -46.060 253.415 -44.835 253.460 ;
        RECT -57.500 249.915 -57.155 253.400 ;
        RECT -69.010 249.470 -57.155 249.915 ;
        RECT -69.010 248.670 -68.670 249.470 ;
        RECT -60.195 249.285 -57.155 249.470 ;
        RECT -69.010 248.500 -67.215 248.670 ;
        RECT -69.010 247.690 -68.670 248.500 ;
        RECT -60.195 248.480 -59.855 249.285 ;
        RECT -60.210 248.180 -59.855 248.480 ;
        RECT -61.665 248.010 -59.855 248.180 ;
        RECT -69.010 247.520 -67.215 247.690 ;
        RECT -69.010 246.710 -68.670 247.520 ;
        RECT -60.210 247.200 -59.855 248.010 ;
        RECT -61.665 247.030 -59.855 247.200 ;
        RECT -69.010 246.540 -67.215 246.710 ;
        RECT -69.010 244.485 -68.670 246.540 ;
        RECT -60.210 246.220 -59.855 247.030 ;
        RECT -61.665 246.050 -59.855 246.220 ;
        RECT -60.210 246.005 -59.855 246.050 ;
        RECT -69.010 244.315 -67.215 244.485 ;
        RECT -60.195 244.395 -59.855 246.005 ;
        RECT -69.010 243.505 -68.670 244.315 ;
        RECT -69.010 243.335 -67.215 243.505 ;
        RECT -69.010 242.525 -68.670 243.335 ;
        RECT -69.010 242.355 -67.215 242.525 ;
        RECT -69.010 242.050 -68.670 242.355 ;
        RECT -69.010 237.560 -68.695 242.050 ;
        RECT -60.185 239.770 -59.870 244.395 ;
        RECT -60.210 239.465 -59.870 239.770 ;
        RECT -61.665 239.295 -59.870 239.465 ;
        RECT -60.210 238.485 -59.870 239.295 ;
        RECT -61.665 238.315 -59.870 238.485 ;
        RECT -69.010 235.170 -68.670 237.560 ;
        RECT -60.210 237.505 -59.870 238.315 ;
        RECT -61.665 237.335 -59.870 237.505 ;
        RECT -69.010 235.000 -67.215 235.170 ;
        RECT -69.010 234.190 -68.670 235.000 ;
        RECT -60.210 234.680 -59.870 237.335 ;
        RECT -61.665 234.510 -59.870 234.680 ;
        RECT -69.010 234.020 -67.215 234.190 ;
        RECT -69.010 233.210 -68.670 234.020 ;
        RECT -60.210 233.700 -59.870 234.510 ;
        RECT -61.665 233.530 -59.870 233.700 ;
        RECT -60.210 233.305 -59.870 233.530 ;
        RECT -69.010 233.040 -67.215 233.210 ;
        RECT -69.010 230.985 -68.670 233.040 ;
        RECT -60.210 232.720 -59.865 233.305 ;
        RECT -61.665 232.550 -59.865 232.720 ;
        RECT -60.210 232.505 -59.865 232.550 ;
        RECT -69.010 230.815 -67.215 230.985 ;
        RECT -60.205 230.940 -59.865 232.505 ;
        RECT -69.010 230.005 -68.670 230.815 ;
        RECT -69.010 229.835 -67.215 230.005 ;
        RECT -69.010 229.025 -68.670 229.835 ;
        RECT -69.010 228.855 -67.215 229.025 ;
        RECT -69.010 228.550 -68.670 228.855 ;
        RECT -69.010 223.790 -68.695 228.550 ;
        RECT -60.185 226.270 -59.870 230.940 ;
        RECT -60.210 225.965 -59.870 226.270 ;
        RECT -61.665 225.795 -59.870 225.965 ;
        RECT -60.210 224.985 -59.870 225.795 ;
        RECT -61.665 224.815 -59.870 224.985 ;
        RECT -60.210 224.005 -59.870 224.815 ;
        RECT -61.665 223.835 -59.870 224.005 ;
        RECT -60.210 221.555 -59.870 223.835 ;
        RECT -61.665 221.385 -59.870 221.555 ;
        RECT -60.210 220.575 -59.870 221.385 ;
        RECT -61.665 220.405 -59.870 220.575 ;
        RECT -60.210 219.595 -59.870 220.405 ;
        RECT -61.665 219.425 -59.870 219.595 ;
        RECT -60.210 219.380 -59.870 219.425 ;
        RECT -71.090 203.480 -70.125 203.705 ;
        RECT -58.680 203.495 -57.725 203.530 ;
        RECT -36.685 203.495 -35.730 203.530 ;
        RECT -71.090 203.445 -68.980 203.480 ;
        RECT -71.090 203.275 -68.030 203.445 ;
        RECT -58.680 203.325 -56.775 203.495 ;
        RECT -37.635 203.325 -35.730 203.495 ;
        RECT -24.285 203.480 -23.320 203.705 ;
        RECT -25.430 203.445 -23.320 203.480 ;
        RECT -58.680 203.300 -57.725 203.325 ;
        RECT -36.685 203.300 -35.730 203.325 ;
        RECT -71.090 203.250 -68.980 203.275 ;
        RECT -71.090 202.495 -69.590 203.250 ;
        RECT -58.680 202.545 -58.335 203.300 ;
        RECT -36.075 202.545 -35.730 203.300 ;
        RECT -26.380 203.275 -23.320 203.445 ;
        RECT -25.430 203.250 -23.320 203.275 ;
        RECT -58.680 202.515 -57.665 202.545 ;
        RECT -36.745 202.515 -35.730 202.545 ;
        RECT -71.090 202.465 -68.920 202.495 ;
        RECT -71.090 202.295 -68.030 202.465 ;
        RECT -58.680 202.345 -56.775 202.515 ;
        RECT -37.635 202.345 -35.730 202.515 ;
        RECT -24.820 202.495 -23.320 203.250 ;
        RECT -17.550 202.855 -13.740 292.690 ;
        RECT -25.490 202.465 -23.320 202.495 ;
        RECT -58.680 202.315 -57.665 202.345 ;
        RECT -36.745 202.315 -35.730 202.345 ;
        RECT -71.090 202.265 -68.920 202.295 ;
        RECT -71.090 201.930 -69.590 202.265 ;
        RECT -58.680 201.980 -58.335 202.315 ;
        RECT -36.075 201.980 -35.730 202.315 ;
        RECT -26.380 202.295 -23.320 202.465 ;
        RECT -25.490 202.265 -23.320 202.295 ;
        RECT -58.680 201.950 -57.715 201.980 ;
        RECT -36.695 201.950 -35.730 201.980 ;
        RECT -71.090 201.900 -68.970 201.930 ;
        RECT -71.090 201.730 -68.030 201.900 ;
        RECT -58.680 201.780 -56.775 201.950 ;
        RECT -37.635 201.780 -35.730 201.950 ;
        RECT -24.820 201.930 -23.320 202.265 ;
        RECT -25.440 201.900 -23.320 201.930 ;
        RECT -58.680 201.750 -57.715 201.780 ;
        RECT -36.695 201.750 -35.730 201.780 ;
        RECT -71.090 201.700 -68.970 201.730 ;
        RECT -71.090 200.950 -69.590 201.700 ;
        RECT -58.680 201.000 -58.335 201.750 ;
        RECT -36.075 201.000 -35.730 201.750 ;
        RECT -26.380 201.730 -23.320 201.900 ;
        RECT -25.440 201.700 -23.320 201.730 ;
        RECT -58.680 200.970 -57.690 201.000 ;
        RECT -36.720 200.970 -35.730 201.000 ;
        RECT -71.090 200.920 -68.945 200.950 ;
        RECT -71.090 200.750 -68.030 200.920 ;
        RECT -58.680 200.800 -56.775 200.970 ;
        RECT -37.635 200.800 -35.730 200.970 ;
        RECT -24.820 201.360 -23.320 201.700 ;
        RECT -18.710 201.360 -12.635 202.855 ;
        RECT -24.820 200.950 -12.635 201.360 ;
        RECT -25.465 200.920 -12.635 200.950 ;
        RECT -58.680 200.770 -57.690 200.800 ;
        RECT -36.720 200.770 -35.730 200.800 ;
        RECT -71.090 200.720 -68.945 200.750 ;
        RECT -71.090 200.385 -69.590 200.720 ;
        RECT -58.680 200.435 -58.335 200.770 ;
        RECT -36.075 200.435 -35.730 200.770 ;
        RECT -26.380 200.750 -12.635 200.920 ;
        RECT -25.465 200.720 -12.635 200.750 ;
        RECT -58.680 200.400 -57.710 200.435 ;
        RECT -36.700 200.400 -35.730 200.435 ;
        RECT -71.090 200.350 -68.965 200.385 ;
        RECT -71.090 200.180 -68.030 200.350 ;
        RECT -58.680 200.230 -56.775 200.400 ;
        RECT -37.635 200.230 -35.730 200.400 ;
        RECT -24.820 200.385 -12.635 200.720 ;
        RECT -25.445 200.350 -12.635 200.385 ;
        RECT -58.680 200.205 -57.710 200.230 ;
        RECT -36.700 200.205 -35.730 200.230 ;
        RECT -71.090 200.155 -68.965 200.180 ;
        RECT -71.090 199.395 -69.590 200.155 ;
        RECT -58.680 199.445 -58.335 200.205 ;
        RECT -36.075 199.445 -35.730 200.205 ;
        RECT -26.380 200.180 -12.635 200.350 ;
        RECT -25.445 200.155 -12.635 200.180 ;
        RECT -58.680 199.420 -57.690 199.445 ;
        RECT -36.720 199.420 -35.730 199.445 ;
        RECT -71.090 199.370 -68.945 199.395 ;
        RECT -71.090 199.200 -68.030 199.370 ;
        RECT -58.680 199.250 -56.775 199.420 ;
        RECT -37.635 199.250 -35.730 199.420 ;
        RECT -24.820 199.395 -12.635 200.155 ;
        RECT -25.465 199.370 -12.635 199.395 ;
        RECT -58.680 199.215 -57.690 199.250 ;
        RECT -36.720 199.215 -35.730 199.250 ;
        RECT -71.090 199.165 -68.945 199.200 ;
        RECT -71.090 198.420 -69.590 199.165 ;
        RECT -58.680 198.880 -58.335 199.215 ;
        RECT -36.075 198.880 -35.730 199.215 ;
        RECT -26.380 199.200 -12.635 199.370 ;
        RECT -25.465 199.165 -12.635 199.200 ;
        RECT -58.815 198.470 -58.135 198.880 ;
        RECT -36.275 198.470 -35.595 198.880 ;
        RECT -58.815 198.440 -57.690 198.470 ;
        RECT -36.720 198.440 -35.595 198.470 ;
        RECT -71.090 198.390 -68.945 198.420 ;
        RECT -71.090 198.220 -68.030 198.390 ;
        RECT -58.815 198.270 -56.775 198.440 ;
        RECT -37.635 198.270 -35.595 198.440 ;
        RECT -24.820 198.420 -12.635 199.165 ;
        RECT -25.465 198.390 -12.635 198.420 ;
        RECT -58.815 198.265 -58.135 198.270 ;
        RECT -36.275 198.265 -35.595 198.270 ;
        RECT -26.380 198.220 -12.635 198.390 ;
        RECT -71.090 187.570 -70.125 198.220 ;
        RECT -24.285 197.550 -12.635 198.220 ;
        RECT -58.820 192.635 -58.140 192.800 ;
        RECT -36.270 192.635 -35.590 192.800 ;
        RECT -58.820 192.465 -56.830 192.635 ;
        RECT -37.580 192.465 -35.590 192.635 ;
        RECT -58.820 192.185 -58.140 192.465 ;
        RECT -36.270 192.185 -35.590 192.465 ;
        RECT -58.655 191.655 -58.310 192.185 ;
        RECT -36.100 191.655 -35.755 192.185 ;
        RECT -58.655 191.485 -56.830 191.655 ;
        RECT -37.580 191.485 -35.755 191.655 ;
        RECT -58.655 190.675 -58.310 191.485 ;
        RECT -36.100 190.675 -35.755 191.485 ;
        RECT -58.655 190.505 -56.830 190.675 ;
        RECT -37.580 190.505 -35.755 190.675 ;
        RECT -58.655 189.885 -58.310 190.505 ;
        RECT -58.680 189.695 -58.310 189.885 ;
        RECT -36.100 189.885 -35.755 190.505 ;
        RECT -36.100 189.695 -35.730 189.885 ;
        RECT -58.680 189.525 -56.830 189.695 ;
        RECT -37.580 189.525 -35.730 189.695 ;
        RECT -69.935 188.445 -68.980 188.480 ;
        RECT -69.935 188.275 -68.030 188.445 ;
        RECT -69.935 188.250 -68.980 188.275 ;
        RECT -69.935 187.570 -69.590 188.250 ;
        RECT -71.090 187.495 -69.590 187.570 ;
        RECT -71.090 187.465 -68.920 187.495 ;
        RECT -71.090 187.295 -68.030 187.465 ;
        RECT -71.090 187.265 -68.920 187.295 ;
        RECT -71.090 186.930 -69.590 187.265 ;
        RECT -58.680 187.010 -58.315 189.525 ;
        RECT -36.095 187.010 -35.730 189.525 ;
        RECT -25.430 188.445 -24.475 188.480 ;
        RECT -26.380 188.275 -24.475 188.445 ;
        RECT -25.430 188.250 -24.475 188.275 ;
        RECT -24.820 187.570 -24.475 188.250 ;
        RECT -24.285 187.570 -23.320 197.550 ;
        RECT -18.710 196.780 -12.635 197.550 ;
        RECT -24.820 187.495 -23.320 187.570 ;
        RECT -25.490 187.465 -23.320 187.495 ;
        RECT -26.380 187.295 -23.320 187.465 ;
        RECT -25.490 187.265 -23.320 187.295 ;
        RECT -58.680 186.985 -58.290 187.010 ;
        RECT -36.120 186.985 -35.730 187.010 ;
        RECT -71.090 186.900 -68.970 186.930 ;
        RECT -71.090 186.730 -68.030 186.900 ;
        RECT -58.680 186.815 -56.830 186.985 ;
        RECT -37.580 186.815 -35.730 186.985 ;
        RECT -24.820 186.930 -23.320 187.265 ;
        RECT -25.440 186.900 -23.320 186.930 ;
        RECT -71.090 186.700 -68.970 186.730 ;
        RECT -71.090 185.950 -69.590 186.700 ;
        RECT -58.680 186.020 -58.290 186.815 ;
        RECT -36.120 186.020 -35.730 186.815 ;
        RECT -26.380 186.730 -23.320 186.900 ;
        RECT -25.440 186.700 -23.320 186.730 ;
        RECT -58.845 186.005 -58.165 186.020 ;
        RECT -36.245 186.005 -35.565 186.020 ;
        RECT -71.090 185.920 -68.945 185.950 ;
        RECT -71.090 185.750 -68.030 185.920 ;
        RECT -58.845 185.835 -56.830 186.005 ;
        RECT -37.580 185.835 -35.565 186.005 ;
        RECT -24.820 185.950 -23.320 186.700 ;
        RECT -25.465 185.920 -23.320 185.950 ;
        RECT -71.090 185.720 -68.945 185.750 ;
        RECT -71.090 185.385 -69.590 185.720 ;
        RECT -58.845 185.405 -58.165 185.835 ;
        RECT -36.245 185.405 -35.565 185.835 ;
        RECT -26.380 185.750 -23.320 185.920 ;
        RECT -25.465 185.720 -23.320 185.750 ;
        RECT -24.820 185.385 -23.320 185.720 ;
        RECT -71.090 185.350 -68.965 185.385 ;
        RECT -25.445 185.350 -23.320 185.385 ;
        RECT -71.090 185.180 -68.030 185.350 ;
        RECT -26.380 185.180 -23.320 185.350 ;
        RECT -71.090 185.155 -68.965 185.180 ;
        RECT -25.445 185.155 -23.320 185.180 ;
        RECT -71.090 184.605 -69.590 185.155 ;
        RECT -71.090 175.505 -70.125 184.605 ;
        RECT -69.935 184.395 -69.590 184.605 ;
        RECT -24.820 184.605 -23.320 185.155 ;
        RECT -24.820 184.395 -24.475 184.605 ;
        RECT -69.935 184.370 -68.945 184.395 ;
        RECT -25.465 184.370 -24.475 184.395 ;
        RECT -69.935 184.200 -68.030 184.370 ;
        RECT -26.380 184.200 -24.475 184.370 ;
        RECT -69.935 184.165 -68.945 184.200 ;
        RECT -25.465 184.165 -24.475 184.200 ;
        RECT -69.935 183.420 -69.590 184.165 ;
        RECT -58.835 183.870 -58.155 184.015 ;
        RECT -36.255 183.870 -35.575 184.015 ;
        RECT -58.835 183.700 -56.205 183.870 ;
        RECT -38.205 183.700 -35.575 183.870 ;
        RECT -69.935 183.390 -68.945 183.420 ;
        RECT -58.835 183.400 -58.155 183.700 ;
        RECT -36.255 183.400 -35.575 183.700 ;
        RECT -24.820 183.420 -24.475 184.165 ;
        RECT -69.935 183.220 -68.030 183.390 ;
        RECT -58.610 182.890 -58.290 183.400 ;
        RECT -36.120 182.890 -35.800 183.400 ;
        RECT -25.465 183.390 -24.475 183.420 ;
        RECT -26.380 183.220 -24.475 183.390 ;
        RECT -58.610 182.720 -56.205 182.890 ;
        RECT -38.205 182.720 -35.800 182.890 ;
        RECT -58.610 181.910 -58.290 182.720 ;
        RECT -36.120 181.910 -35.800 182.720 ;
        RECT -58.610 181.740 -56.205 181.910 ;
        RECT -38.205 181.740 -35.800 181.910 ;
        RECT -58.610 181.710 -58.040 181.740 ;
        RECT -58.535 180.825 -58.040 181.710 ;
        RECT -36.370 181.710 -35.800 181.740 ;
        RECT -36.370 180.825 -35.875 181.710 ;
        RECT -58.535 180.655 -57.210 180.825 ;
        RECT -37.200 180.655 -35.875 180.825 ;
        RECT -58.535 179.845 -58.040 180.655 ;
        RECT -36.370 179.845 -35.875 180.655 ;
        RECT -58.535 179.675 -57.210 179.845 ;
        RECT -37.200 179.675 -35.875 179.845 ;
        RECT -58.535 178.865 -58.040 179.675 ;
        RECT -36.370 178.865 -35.875 179.675 ;
        RECT -58.535 178.695 -57.210 178.865 ;
        RECT -37.200 178.695 -35.875 178.865 ;
        RECT -58.535 177.885 -58.040 178.695 ;
        RECT -36.370 177.885 -35.875 178.695 ;
        RECT -58.535 177.875 -57.210 177.885 ;
        RECT -58.720 177.715 -57.210 177.875 ;
        RECT -37.200 177.875 -35.875 177.885 ;
        RECT -37.200 177.715 -35.690 177.875 ;
        RECT -58.720 177.260 -58.040 177.715 ;
        RECT -36.370 177.260 -35.690 177.715 ;
        RECT -69.935 175.945 -68.980 175.980 ;
        RECT -25.430 175.945 -24.475 175.980 ;
        RECT -69.935 175.775 -68.030 175.945 ;
        RECT -58.715 175.845 -58.035 175.930 ;
        RECT -36.375 175.845 -35.695 175.930 ;
        RECT -69.935 175.750 -68.980 175.775 ;
        RECT -69.935 175.505 -69.590 175.750 ;
        RECT -71.090 174.995 -69.590 175.505 ;
        RECT -58.715 175.675 -56.215 175.845 ;
        RECT -38.195 175.675 -35.695 175.845 ;
        RECT -26.380 175.775 -24.475 175.945 ;
        RECT -25.430 175.750 -24.475 175.775 ;
        RECT -58.715 175.315 -58.035 175.675 ;
        RECT -36.375 175.315 -35.695 175.675 ;
        RECT -24.820 175.505 -24.475 175.750 ;
        RECT -24.285 175.505 -23.320 184.605 ;
        RECT -71.090 174.965 -68.920 174.995 ;
        RECT -71.090 174.795 -68.030 174.965 ;
        RECT -58.645 174.865 -58.250 175.315 ;
        RECT -36.160 174.865 -35.765 175.315 ;
        RECT -24.820 174.995 -23.320 175.505 ;
        RECT -25.490 174.965 -23.320 174.995 ;
        RECT -71.090 174.765 -68.920 174.795 ;
        RECT -71.090 174.430 -69.590 174.765 ;
        RECT -58.645 174.695 -56.215 174.865 ;
        RECT -38.195 174.695 -35.765 174.865 ;
        RECT -26.380 174.795 -23.320 174.965 ;
        RECT -25.490 174.765 -23.320 174.795 ;
        RECT -71.090 174.400 -68.970 174.430 ;
        RECT -71.090 174.230 -68.030 174.400 ;
        RECT -71.090 174.200 -68.970 174.230 ;
        RECT -71.090 173.450 -69.590 174.200 ;
        RECT -58.645 173.885 -58.250 174.695 ;
        RECT -36.160 173.885 -35.765 174.695 ;
        RECT -24.820 174.430 -23.320 174.765 ;
        RECT -25.440 174.400 -23.320 174.430 ;
        RECT -26.380 174.230 -23.320 174.400 ;
        RECT -25.440 174.200 -23.320 174.230 ;
        RECT -58.645 173.715 -56.215 173.885 ;
        RECT -38.195 173.715 -35.765 173.885 ;
        RECT -71.090 173.420 -68.945 173.450 ;
        RECT -71.090 173.250 -68.030 173.420 ;
        RECT -71.090 173.220 -68.945 173.250 ;
        RECT -71.090 172.885 -69.590 173.220 ;
        RECT -71.090 172.850 -68.965 172.885 ;
        RECT -71.090 172.680 -68.030 172.850 ;
        RECT -58.645 172.800 -58.050 173.715 ;
        RECT -36.360 172.800 -35.765 173.715 ;
        RECT -24.820 173.450 -23.320 174.200 ;
        RECT -25.465 173.420 -23.320 173.450 ;
        RECT -26.380 173.250 -23.320 173.420 ;
        RECT -25.465 173.220 -23.320 173.250 ;
        RECT -24.820 172.885 -23.320 173.220 ;
        RECT -25.445 172.850 -23.320 172.885 ;
        RECT -71.090 172.655 -68.965 172.680 ;
        RECT -71.090 172.540 -69.590 172.655 ;
        RECT -71.090 165.680 -70.125 172.540 ;
        RECT -69.935 171.895 -69.590 172.540 ;
        RECT -58.645 172.630 -57.220 172.800 ;
        RECT -37.190 172.630 -35.765 172.800 ;
        RECT -26.380 172.680 -23.320 172.850 ;
        RECT -25.445 172.655 -23.320 172.680 ;
        RECT -69.935 171.870 -68.945 171.895 ;
        RECT -69.935 171.700 -68.030 171.870 ;
        RECT -58.645 171.820 -58.050 172.630 ;
        RECT -36.360 171.820 -35.765 172.630 ;
        RECT -24.820 172.540 -23.320 172.655 ;
        RECT -24.820 171.895 -24.475 172.540 ;
        RECT -25.465 171.870 -24.475 171.895 ;
        RECT -69.935 171.665 -68.945 171.700 ;
        RECT -69.935 170.920 -69.590 171.665 ;
        RECT -58.645 171.650 -57.220 171.820 ;
        RECT -37.190 171.650 -35.765 171.820 ;
        RECT -26.380 171.700 -24.475 171.870 ;
        RECT -25.465 171.665 -24.475 171.700 ;
        RECT -69.935 170.890 -68.945 170.920 ;
        RECT -69.935 170.720 -68.030 170.890 ;
        RECT -58.645 170.840 -58.050 171.650 ;
        RECT -36.360 170.840 -35.765 171.650 ;
        RECT -24.820 170.920 -24.475 171.665 ;
        RECT -25.465 170.890 -24.475 170.920 ;
        RECT -58.645 170.670 -57.220 170.840 ;
        RECT -37.190 170.670 -35.765 170.840 ;
        RECT -26.380 170.720 -24.475 170.890 ;
        RECT -58.645 169.860 -58.050 170.670 ;
        RECT -36.360 169.860 -35.765 170.670 ;
        RECT -58.645 169.690 -57.220 169.860 ;
        RECT -37.190 169.690 -35.765 169.860 ;
        RECT -58.645 169.450 -58.050 169.690 ;
        RECT -36.360 169.450 -35.765 169.690 ;
        RECT -58.645 167.825 -58.250 169.450 ;
        RECT -36.160 167.825 -35.765 169.450 ;
        RECT -58.645 167.655 -56.785 167.825 ;
        RECT -37.625 167.655 -35.765 167.825 ;
        RECT -58.645 166.845 -58.250 167.655 ;
        RECT -36.160 166.845 -35.765 167.655 ;
        RECT -58.645 166.675 -56.785 166.845 ;
        RECT -37.625 166.675 -35.765 166.845 ;
        RECT -65.765 165.680 -65.085 165.695 ;
        RECT -62.995 165.690 -62.685 166.605 ;
        RECT -71.090 165.105 -65.085 165.680 ;
        RECT -71.090 162.835 -70.125 165.105 ;
        RECT -65.765 165.080 -65.085 165.105 ;
        RECT -63.000 165.675 -62.685 165.690 ;
        RECT -58.645 165.865 -58.250 166.675 ;
        RECT -36.160 165.865 -35.765 166.675 ;
        RECT -58.645 165.695 -56.785 165.865 ;
        RECT -37.625 165.695 -35.765 165.865 ;
        RECT -58.645 165.675 -58.250 165.695 ;
        RECT -63.000 165.100 -58.250 165.675 ;
        RECT -63.000 165.075 -62.685 165.100 ;
        RECT -58.645 164.885 -58.250 165.100 ;
        RECT -36.160 165.675 -35.765 165.695 ;
        RECT -31.725 165.690 -31.415 166.605 ;
        RECT -31.725 165.675 -31.410 165.690 ;
        RECT -36.160 165.100 -31.410 165.675 ;
        RECT -36.160 164.885 -35.765 165.100 ;
        RECT -31.725 165.075 -31.410 165.100 ;
        RECT -29.325 165.680 -28.645 165.695 ;
        RECT -24.285 165.680 -23.320 172.540 ;
        RECT -29.325 165.105 -23.320 165.680 ;
        RECT -29.325 165.080 -28.645 165.105 ;
        RECT -58.645 164.715 -56.785 164.885 ;
        RECT -37.625 164.715 -35.765 164.885 ;
        RECT -69.935 163.445 -68.980 163.480 ;
        RECT -69.935 163.275 -68.030 163.445 ;
        RECT -69.935 163.250 -68.980 163.275 ;
        RECT -69.935 162.835 -69.590 163.250 ;
        RECT -71.090 162.495 -69.590 162.835 ;
        RECT -71.090 162.465 -68.920 162.495 ;
        RECT -71.090 162.295 -68.030 162.465 ;
        RECT -71.090 162.265 -68.920 162.295 ;
        RECT -71.090 161.930 -69.590 162.265 ;
        RECT -58.645 162.200 -58.250 164.715 ;
        RECT -36.160 162.200 -35.765 164.715 ;
        RECT -25.430 163.445 -24.475 163.480 ;
        RECT -26.380 163.275 -24.475 163.445 ;
        RECT -25.430 163.250 -24.475 163.275 ;
        RECT -24.820 162.835 -24.475 163.250 ;
        RECT -24.285 162.835 -23.320 165.105 ;
        RECT -24.820 162.495 -23.320 162.835 ;
        RECT -25.490 162.465 -23.320 162.495 ;
        RECT -26.380 162.295 -23.320 162.465 ;
        RECT -25.490 162.265 -23.320 162.295 ;
        RECT -58.645 162.175 -58.245 162.200 ;
        RECT -36.165 162.175 -35.765 162.200 ;
        RECT -58.645 162.005 -56.785 162.175 ;
        RECT -37.625 162.005 -35.765 162.175 ;
        RECT -71.090 161.900 -68.970 161.930 ;
        RECT -71.090 161.730 -68.030 161.900 ;
        RECT -71.090 161.700 -68.970 161.730 ;
        RECT -71.090 160.950 -69.590 161.700 ;
        RECT -58.645 161.195 -58.245 162.005 ;
        RECT -36.165 161.195 -35.765 162.005 ;
        RECT -24.820 161.930 -23.320 162.265 ;
        RECT -25.440 161.900 -23.320 161.930 ;
        RECT -26.380 161.730 -23.320 161.900 ;
        RECT -25.440 161.700 -23.320 161.730 ;
        RECT -58.645 161.040 -56.785 161.195 ;
        RECT -58.780 161.025 -56.785 161.040 ;
        RECT -37.625 161.040 -35.765 161.195 ;
        RECT -37.625 161.025 -35.630 161.040 ;
        RECT -71.090 160.920 -68.945 160.950 ;
        RECT -71.090 160.750 -68.030 160.920 ;
        RECT -71.090 160.720 -68.945 160.750 ;
        RECT -71.090 160.385 -69.590 160.720 ;
        RECT -58.780 160.425 -58.100 161.025 ;
        RECT -36.310 160.425 -35.630 161.025 ;
        RECT -24.820 160.950 -23.320 161.700 ;
        RECT -25.465 160.920 -23.320 160.950 ;
        RECT -26.380 160.750 -23.320 160.920 ;
        RECT -25.465 160.720 -23.320 160.750 ;
        RECT -24.820 160.385 -23.320 160.720 ;
        RECT -71.090 160.350 -68.965 160.385 ;
        RECT -25.445 160.350 -23.320 160.385 ;
        RECT -71.090 160.180 -68.030 160.350 ;
        RECT -26.380 160.180 -23.320 160.350 ;
        RECT -71.090 160.155 -68.965 160.180 ;
        RECT -25.445 160.155 -23.320 160.180 ;
        RECT -71.090 159.870 -69.590 160.155 ;
        RECT -71.090 153.265 -70.125 159.870 ;
        RECT -69.935 159.395 -69.590 159.870 ;
        RECT -24.820 159.870 -23.320 160.155 ;
        RECT -58.775 159.485 -58.095 159.570 ;
        RECT -36.315 159.485 -35.635 159.570 ;
        RECT -69.935 159.370 -68.945 159.395 ;
        RECT -69.935 159.200 -68.030 159.370 ;
        RECT -58.775 159.315 -56.870 159.485 ;
        RECT -37.540 159.315 -35.635 159.485 ;
        RECT -24.820 159.395 -24.475 159.870 ;
        RECT -25.465 159.370 -24.475 159.395 ;
        RECT -69.935 159.165 -68.945 159.200 ;
        RECT -69.935 158.420 -69.590 159.165 ;
        RECT -58.775 158.955 -58.095 159.315 ;
        RECT -36.315 158.955 -35.635 159.315 ;
        RECT -26.380 159.200 -24.475 159.370 ;
        RECT -25.465 159.165 -24.475 159.200 ;
        RECT -58.665 158.505 -58.325 158.955 ;
        RECT -36.085 158.505 -35.745 158.955 ;
        RECT -69.935 158.390 -68.945 158.420 ;
        RECT -69.935 158.220 -68.030 158.390 ;
        RECT -58.665 158.335 -56.870 158.505 ;
        RECT -37.540 158.335 -35.745 158.505 ;
        RECT -24.820 158.420 -24.475 159.165 ;
        RECT -25.465 158.390 -24.475 158.420 ;
        RECT -58.665 157.525 -58.325 158.335 ;
        RECT -36.085 157.525 -35.745 158.335 ;
        RECT -26.380 158.220 -24.475 158.390 ;
        RECT -58.665 157.355 -56.870 157.525 ;
        RECT -37.540 157.355 -35.745 157.525 ;
        RECT -58.665 155.075 -58.325 157.355 ;
        RECT -58.665 154.905 -56.870 155.075 ;
        RECT -58.665 154.095 -58.325 154.905 ;
        RECT -58.665 153.925 -56.870 154.095 ;
        RECT -65.765 153.265 -65.085 153.280 ;
        RECT -71.090 152.695 -65.085 153.265 ;
        RECT -71.090 150.255 -70.125 152.695 ;
        RECT -65.765 152.665 -65.085 152.695 ;
        RECT -62.825 153.255 -62.145 153.275 ;
        RECT -58.665 153.255 -58.325 153.925 ;
        RECT -62.825 153.115 -58.325 153.255 ;
        RECT -62.825 152.945 -56.870 153.115 ;
        RECT -62.825 152.680 -58.325 152.945 ;
        RECT -62.825 152.660 -62.145 152.680 ;
        RECT -58.665 152.640 -58.325 152.680 ;
        RECT -49.840 152.875 -49.525 155.120 ;
        RECT -44.885 152.875 -44.570 155.120 ;
        RECT -36.085 155.075 -35.745 157.355 ;
        RECT -37.540 154.905 -35.745 155.075 ;
        RECT -36.085 154.095 -35.745 154.905 ;
        RECT -37.540 153.925 -35.745 154.095 ;
        RECT -36.085 153.255 -35.745 153.925 ;
        RECT -32.265 153.255 -31.585 153.275 ;
        RECT -36.085 153.115 -31.585 153.255 ;
        RECT -37.540 152.945 -31.585 153.115 ;
        RECT -69.935 150.945 -68.980 150.980 ;
        RECT -69.935 150.775 -68.030 150.945 ;
        RECT -69.935 150.750 -68.980 150.775 ;
        RECT -69.935 150.255 -69.590 150.750 ;
        RECT -71.090 149.995 -69.590 150.255 ;
        RECT -71.090 149.965 -68.920 149.995 ;
        RECT -71.090 149.795 -68.030 149.965 ;
        RECT -71.090 149.765 -68.920 149.795 ;
        RECT -71.090 149.430 -69.590 149.765 ;
        RECT -71.090 149.400 -68.970 149.430 ;
        RECT -71.090 149.230 -68.030 149.400 ;
        RECT -71.090 149.200 -68.970 149.230 ;
        RECT -71.090 148.450 -69.590 149.200 ;
        RECT -71.090 148.420 -68.945 148.450 ;
        RECT -71.090 148.250 -68.030 148.420 ;
        RECT -71.090 148.220 -68.945 148.250 ;
        RECT -71.090 147.885 -69.590 148.220 ;
        RECT -58.665 147.970 -58.350 152.640 ;
        RECT -49.840 151.530 -44.570 152.875 ;
        RECT -36.085 152.680 -31.585 152.945 ;
        RECT -36.085 152.640 -35.745 152.680 ;
        RECT -32.265 152.660 -31.585 152.680 ;
        RECT -29.325 153.265 -28.645 153.280 ;
        RECT -24.285 153.265 -23.320 159.870 ;
        RECT -29.325 152.695 -23.320 153.265 ;
        RECT -29.325 152.665 -28.645 152.695 ;
        RECT -49.840 150.360 -49.525 151.530 ;
        RECT -49.865 150.055 -49.525 150.360 ;
        RECT -51.320 149.885 -49.525 150.055 ;
        RECT -49.865 149.075 -49.525 149.885 ;
        RECT -51.320 148.905 -49.525 149.075 ;
        RECT -49.865 148.095 -49.525 148.905 ;
        RECT -71.090 147.850 -68.965 147.885 ;
        RECT -71.090 147.680 -68.030 147.850 ;
        RECT -71.090 147.655 -68.965 147.680 ;
        RECT -71.090 147.290 -69.590 147.655 ;
        RECT -71.090 140.430 -70.125 147.290 ;
        RECT -69.935 146.895 -69.590 147.290 ;
        RECT -69.935 146.870 -68.945 146.895 ;
        RECT -69.935 146.700 -68.030 146.870 ;
        RECT -69.935 146.665 -68.945 146.700 ;
        RECT -69.935 145.920 -69.590 146.665 ;
        RECT -58.670 146.405 -58.330 147.970 ;
        RECT -51.320 147.925 -49.525 148.095 ;
        RECT -49.865 147.720 -49.525 147.925 ;
        RECT -44.885 150.360 -44.570 151.530 ;
        RECT -44.885 150.055 -44.545 150.360 ;
        RECT -44.885 149.885 -43.090 150.055 ;
        RECT -44.885 149.075 -44.545 149.885 ;
        RECT -44.885 148.905 -43.090 149.075 ;
        RECT -44.885 148.095 -44.545 148.905 ;
        RECT -44.885 147.925 -43.090 148.095 ;
        RECT -36.060 147.970 -35.745 152.640 ;
        RECT -25.430 150.945 -24.475 150.980 ;
        RECT -26.380 150.775 -24.475 150.945 ;
        RECT -25.430 150.750 -24.475 150.775 ;
        RECT -24.820 150.255 -24.475 150.750 ;
        RECT -24.285 150.255 -23.320 152.695 ;
        RECT -24.820 149.995 -23.320 150.255 ;
        RECT -25.490 149.965 -23.320 149.995 ;
        RECT -26.380 149.795 -23.320 149.965 ;
        RECT -25.490 149.765 -23.320 149.795 ;
        RECT -24.820 149.430 -23.320 149.765 ;
        RECT -25.440 149.400 -23.320 149.430 ;
        RECT -26.380 149.230 -23.320 149.400 ;
        RECT -25.440 149.200 -23.320 149.230 ;
        RECT -24.820 148.450 -23.320 149.200 ;
        RECT -25.465 148.420 -23.320 148.450 ;
        RECT -26.380 148.250 -23.320 148.420 ;
        RECT -25.465 148.220 -23.320 148.250 ;
        RECT -44.885 147.720 -44.545 147.925 ;
        RECT -58.670 146.360 -58.325 146.405 ;
        RECT -49.865 146.375 -44.545 147.720 ;
        RECT -36.080 146.405 -35.740 147.970 ;
        RECT -24.820 147.885 -23.320 148.220 ;
        RECT -25.445 147.850 -23.320 147.885 ;
        RECT -26.380 147.680 -23.320 147.850 ;
        RECT -25.445 147.655 -23.320 147.680 ;
        RECT -24.820 147.290 -23.320 147.655 ;
        RECT -24.820 146.895 -24.475 147.290 ;
        RECT -25.465 146.870 -24.475 146.895 ;
        RECT -26.380 146.700 -24.475 146.870 ;
        RECT -25.465 146.665 -24.475 146.700 ;
        RECT -58.670 146.190 -56.870 146.360 ;
        RECT -69.935 145.890 -68.945 145.920 ;
        RECT -69.935 145.720 -68.030 145.890 ;
        RECT -58.670 145.605 -58.325 146.190 ;
        RECT -49.865 145.870 -49.525 146.375 ;
        RECT -51.320 145.700 -49.525 145.870 ;
        RECT -58.665 145.380 -58.325 145.605 ;
        RECT -58.665 145.210 -56.870 145.380 ;
        RECT -58.665 144.400 -58.325 145.210 ;
        RECT -49.865 144.890 -49.525 145.700 ;
        RECT -51.320 144.720 -49.525 144.890 ;
        RECT -58.665 144.230 -56.870 144.400 ;
        RECT -58.665 141.575 -58.325 144.230 ;
        RECT -49.865 143.910 -49.525 144.720 ;
        RECT -51.320 143.740 -49.525 143.910 ;
        RECT -49.865 143.205 -49.525 143.740 ;
        RECT -44.885 145.870 -44.545 146.375 ;
        RECT -36.085 146.360 -35.740 146.405 ;
        RECT -37.540 146.190 -35.740 146.360 ;
        RECT -44.885 145.700 -43.090 145.870 ;
        RECT -44.885 144.890 -44.545 145.700 ;
        RECT -36.085 145.605 -35.740 146.190 ;
        RECT -24.820 145.920 -24.475 146.665 ;
        RECT -25.465 145.890 -24.475 145.920 ;
        RECT -26.380 145.720 -24.475 145.890 ;
        RECT -36.085 145.380 -35.745 145.605 ;
        RECT -37.540 145.210 -35.745 145.380 ;
        RECT -44.885 144.720 -43.090 144.890 ;
        RECT -44.885 143.910 -44.545 144.720 ;
        RECT -36.085 144.400 -35.745 145.210 ;
        RECT -37.540 144.230 -35.745 144.400 ;
        RECT -44.885 143.740 -43.090 143.910 ;
        RECT -44.885 143.205 -44.545 143.740 ;
        RECT -49.865 141.860 -44.545 143.205 ;
        RECT -58.665 141.405 -56.870 141.575 ;
        RECT -58.665 140.595 -58.325 141.405 ;
        RECT -49.865 141.350 -49.525 141.860 ;
        RECT -65.940 140.430 -65.260 140.445 ;
        RECT -71.090 139.855 -65.260 140.430 ;
        RECT -71.090 138.480 -70.125 139.855 ;
        RECT -65.940 139.830 -65.260 139.855 ;
        RECT -62.105 140.425 -61.425 140.440 ;
        RECT -58.665 140.425 -56.870 140.595 ;
        RECT -62.105 139.850 -58.325 140.425 ;
        RECT -62.105 139.825 -61.425 139.850 ;
        RECT -58.665 139.615 -58.325 139.850 ;
        RECT -58.665 139.445 -56.870 139.615 ;
        RECT -58.665 139.140 -58.325 139.445 ;
        RECT -71.090 138.445 -68.980 138.480 ;
        RECT -71.090 138.275 -68.030 138.445 ;
        RECT -71.090 138.250 -68.980 138.275 ;
        RECT -71.090 137.495 -69.590 138.250 ;
        RECT -71.090 137.465 -68.920 137.495 ;
        RECT -71.090 137.295 -68.030 137.465 ;
        RECT -71.090 137.265 -68.920 137.295 ;
        RECT -71.090 136.930 -69.590 137.265 ;
        RECT -71.090 136.900 -68.970 136.930 ;
        RECT -71.090 136.730 -68.030 136.900 ;
        RECT -71.090 136.700 -68.970 136.730 ;
        RECT -71.090 135.950 -69.590 136.700 ;
        RECT -71.090 135.920 -68.945 135.950 ;
        RECT -71.090 135.750 -68.030 135.920 ;
        RECT -71.090 135.720 -68.945 135.750 ;
        RECT -71.090 135.385 -69.590 135.720 ;
        RECT -71.090 135.350 -68.965 135.385 ;
        RECT -71.090 135.180 -68.030 135.350 ;
        RECT -71.090 135.155 -68.965 135.180 ;
        RECT -71.090 134.395 -69.590 135.155 ;
        RECT -58.665 134.515 -58.350 139.140 ;
        RECT -49.840 138.895 -49.525 141.350 ;
        RECT -44.885 141.350 -44.545 141.860 ;
        RECT -36.085 141.575 -35.745 144.230 ;
        RECT -37.540 141.405 -35.745 141.575 ;
        RECT -44.885 138.895 -44.570 141.350 ;
        RECT -36.085 140.595 -35.745 141.405 ;
        RECT -37.540 140.425 -35.745 140.595 ;
        RECT -32.985 140.425 -32.305 140.440 ;
        RECT -36.085 139.850 -32.305 140.425 ;
        RECT -36.085 139.615 -35.745 139.850 ;
        RECT -32.985 139.825 -32.305 139.850 ;
        RECT -29.150 140.430 -28.470 140.445 ;
        RECT -24.285 140.430 -23.320 147.290 ;
        RECT -29.150 139.855 -23.320 140.430 ;
        RECT -29.150 139.830 -28.470 139.855 ;
        RECT -37.540 139.445 -35.745 139.615 ;
        RECT -36.085 139.140 -35.745 139.445 ;
        RECT -49.840 137.550 -44.570 138.895 ;
        RECT -49.840 136.860 -49.525 137.550 ;
        RECT -49.865 136.555 -49.525 136.860 ;
        RECT -51.320 136.385 -49.525 136.555 ;
        RECT -49.865 135.575 -49.525 136.385 ;
        RECT -51.320 135.405 -49.525 135.575 ;
        RECT -49.865 134.595 -49.525 135.405 ;
        RECT -71.090 134.370 -68.945 134.395 ;
        RECT -71.090 134.200 -68.030 134.370 ;
        RECT -71.090 134.165 -68.945 134.200 ;
        RECT -71.090 133.420 -69.590 134.165 ;
        RECT -71.090 133.390 -68.945 133.420 ;
        RECT -71.090 133.220 -68.030 133.390 ;
        RECT -71.090 128.895 -70.125 133.220 ;
        RECT -58.680 132.905 -58.340 134.515 ;
        RECT -51.320 134.510 -49.525 134.595 ;
        RECT -44.885 136.860 -44.570 137.550 ;
        RECT -44.885 136.555 -44.545 136.860 ;
        RECT -44.885 136.385 -43.090 136.555 ;
        RECT -44.885 135.575 -44.545 136.385 ;
        RECT -44.885 135.405 -43.090 135.575 ;
        RECT -44.885 134.595 -44.545 135.405 ;
        RECT -44.885 134.510 -43.090 134.595 ;
        RECT -36.060 134.515 -35.745 139.140 ;
        RECT -24.285 138.480 -23.320 139.855 ;
        RECT -25.430 138.445 -23.320 138.480 ;
        RECT -26.380 138.275 -23.320 138.445 ;
        RECT -25.430 138.250 -23.320 138.275 ;
        RECT -24.820 137.495 -23.320 138.250 ;
        RECT -25.490 137.465 -23.320 137.495 ;
        RECT -26.380 137.295 -23.320 137.465 ;
        RECT -25.490 137.265 -23.320 137.295 ;
        RECT -24.820 136.930 -23.320 137.265 ;
        RECT -25.440 136.900 -23.320 136.930 ;
        RECT -26.380 136.730 -23.320 136.900 ;
        RECT -25.440 136.700 -23.320 136.730 ;
        RECT -24.820 135.950 -23.320 136.700 ;
        RECT -25.465 135.920 -23.320 135.950 ;
        RECT -26.380 135.750 -23.320 135.920 ;
        RECT -25.465 135.720 -23.320 135.750 ;
        RECT -24.820 135.385 -23.320 135.720 ;
        RECT -25.445 135.350 -23.320 135.385 ;
        RECT -26.380 135.180 -23.320 135.350 ;
        RECT -25.445 135.155 -23.320 135.180 ;
        RECT -51.320 134.425 -43.090 134.510 ;
        RECT -49.865 133.165 -44.545 134.425 ;
        RECT -58.680 132.860 -58.325 132.905 ;
        RECT -58.680 132.690 -56.870 132.860 ;
        RECT -58.680 131.880 -58.325 132.690 ;
        RECT -49.865 132.370 -49.525 133.165 ;
        RECT -51.320 132.200 -49.525 132.370 ;
        RECT -58.680 131.710 -56.870 131.880 ;
        RECT -49.865 131.780 -49.525 132.200 ;
        RECT -44.885 132.370 -44.545 133.165 ;
        RECT -36.070 133.825 -35.730 134.515 ;
        RECT -24.820 134.395 -23.320 135.155 ;
        RECT -25.465 134.370 -23.320 134.395 ;
        RECT -26.380 134.200 -23.320 134.370 ;
        RECT -25.465 134.165 -23.320 134.200 ;
        RECT -33.780 133.825 -33.440 133.955 ;
        RECT -36.070 133.655 -33.440 133.825 ;
        RECT -36.070 133.485 -31.985 133.655 ;
        RECT -36.070 133.385 -33.440 133.485 ;
        RECT -24.820 133.420 -23.320 134.165 ;
        RECT -25.465 133.390 -23.320 133.420 ;
        RECT -36.070 132.915 -35.730 133.385 ;
        RECT -33.780 132.915 -33.440 133.385 ;
        RECT -26.380 133.220 -23.320 133.390 ;
        RECT -36.070 132.905 -33.440 132.915 ;
        RECT -36.085 132.860 -33.440 132.905 ;
        RECT -37.540 132.690 -33.440 132.860 ;
        RECT -36.085 132.675 -33.440 132.690 ;
        RECT -36.085 132.505 -31.985 132.675 ;
        RECT -36.085 132.475 -33.440 132.505 ;
        RECT -44.885 132.200 -43.090 132.370 ;
        RECT -44.885 131.780 -44.545 132.200 ;
        RECT -36.085 132.000 -35.730 132.475 ;
        RECT -33.780 132.000 -33.440 132.475 ;
        RECT -36.085 131.880 -33.440 132.000 ;
        RECT -58.680 130.900 -58.325 131.710 ;
        RECT -49.865 131.390 -44.545 131.780 ;
        RECT -37.540 131.710 -33.440 131.880 ;
        RECT -36.085 131.695 -33.440 131.710 ;
        RECT -36.085 131.560 -31.985 131.695 ;
        RECT -51.320 131.220 -43.090 131.390 ;
        RECT -58.680 130.730 -56.870 130.900 ;
        RECT -58.680 130.430 -58.325 130.730 ;
        RECT -49.865 130.435 -44.545 131.220 ;
        RECT -36.085 130.900 -35.730 131.560 ;
        RECT -33.780 131.525 -31.985 131.560 ;
        RECT -33.780 131.480 -33.440 131.525 ;
        RECT -37.540 130.730 -35.730 130.900 ;
        RECT -58.680 129.440 -58.340 130.430 ;
        RECT -49.865 130.410 -49.525 130.435 ;
        RECT -51.320 130.240 -49.525 130.410 ;
        RECT -49.865 129.445 -49.525 130.240 ;
        RECT -44.885 130.410 -44.545 130.435 ;
        RECT -36.085 130.430 -35.730 130.730 ;
        RECT -44.885 130.240 -43.090 130.410 ;
        RECT -49.865 129.440 -49.080 129.445 ;
        RECT -44.885 129.440 -44.545 130.240 ;
        RECT -36.070 129.440 -35.730 130.430 ;
        RECT -58.680 128.995 -35.730 129.440 ;
        RECT -48.505 126.105 -48.080 128.995 ;
        RECT -24.285 126.405 -23.320 133.220 ;
        RECT -24.285 126.395 -23.375 126.405 ;
        RECT -49.120 126.080 -48.080 126.105 ;
        RECT -52.070 125.910 -48.080 126.080 ;
        RECT -23.820 125.970 -23.375 126.395 ;
        RECT -24.450 125.945 -23.375 125.970 ;
        RECT -49.120 125.880 -48.080 125.910 ;
        RECT -48.505 125.130 -48.080 125.880 ;
        RECT -27.400 125.775 -23.375 125.945 ;
        RECT -24.450 125.745 -23.375 125.775 ;
        RECT -49.105 125.100 -48.080 125.130 ;
        RECT -52.070 124.930 -48.080 125.100 ;
        RECT -23.820 124.995 -23.375 125.745 ;
        RECT -24.435 124.965 -23.375 124.995 ;
        RECT -49.105 124.905 -48.080 124.930 ;
        RECT -48.505 123.020 -48.080 124.905 ;
        RECT -27.400 124.795 -23.375 124.965 ;
        RECT -24.435 124.770 -23.375 124.795 ;
        RECT -49.110 122.985 -48.080 123.020 ;
        RECT -52.070 122.815 -48.080 122.985 ;
        RECT -23.820 122.885 -23.375 124.770 ;
        RECT -24.440 122.850 -23.375 122.885 ;
        RECT -49.110 122.795 -48.080 122.815 ;
        RECT -57.330 120.115 -56.990 120.160 ;
        RECT -57.330 119.945 -55.535 120.115 ;
        RECT -57.330 119.135 -56.990 119.945 ;
        RECT -57.330 118.965 -55.535 119.135 ;
        RECT -57.330 118.155 -56.990 118.965 ;
        RECT -57.330 117.985 -55.535 118.155 ;
        RECT -57.330 115.705 -56.990 117.985 ;
        RECT -57.330 115.535 -55.535 115.705 ;
        RECT -57.330 114.725 -56.990 115.535 ;
        RECT -57.330 114.555 -55.535 114.725 ;
        RECT -57.330 113.745 -56.990 114.555 ;
        RECT -57.330 113.575 -55.535 113.745 ;
        RECT -57.330 113.270 -56.990 113.575 ;
        RECT -57.330 108.600 -57.015 113.270 ;
        RECT -48.505 110.990 -48.080 122.795 ;
        RECT -27.400 122.680 -23.375 122.850 ;
        RECT -24.440 122.660 -23.375 122.680 ;
        RECT -48.530 110.685 -48.080 110.990 ;
        RECT -49.985 110.515 -48.080 110.685 ;
        RECT -48.530 110.015 -48.080 110.515 ;
        RECT -32.695 120.115 -32.355 120.160 ;
        RECT -32.695 119.945 -30.900 120.115 ;
        RECT -32.695 119.135 -32.355 119.945 ;
        RECT -32.695 118.965 -30.900 119.135 ;
        RECT -32.695 118.155 -32.355 118.965 ;
        RECT -32.695 117.985 -30.900 118.155 ;
        RECT -32.695 115.705 -32.355 117.985 ;
        RECT -23.820 115.750 -23.375 122.660 ;
        RECT -32.695 115.535 -30.900 115.705 ;
        RECT -32.695 114.725 -32.355 115.535 ;
        RECT -23.870 114.750 -23.375 115.750 ;
        RECT -32.695 114.555 -30.900 114.725 ;
        RECT -32.695 113.745 -32.355 114.555 ;
        RECT -32.695 113.575 -30.900 113.745 ;
        RECT -32.695 113.270 -32.355 113.575 ;
        RECT -48.530 109.705 -48.190 110.015 ;
        RECT -49.985 109.535 -48.190 109.705 ;
        RECT -48.530 108.725 -48.190 109.535 ;
        RECT -57.335 107.035 -56.995 108.600 ;
        RECT -49.985 108.555 -48.190 108.725 ;
        RECT -32.695 108.600 -32.380 113.270 ;
        RECT -23.870 110.990 -23.555 114.750 ;
        RECT -23.895 110.685 -23.555 110.990 ;
        RECT -25.350 110.515 -23.555 110.685 ;
        RECT -23.895 109.705 -23.555 110.515 ;
        RECT -25.350 109.535 -23.555 109.705 ;
        RECT -23.895 108.725 -23.555 109.535 ;
        RECT -57.335 106.990 -56.990 107.035 ;
        RECT -57.335 106.820 -55.535 106.990 ;
        RECT -57.335 106.235 -56.990 106.820 ;
        RECT -48.530 106.500 -48.190 108.555 ;
        RECT -42.750 107.145 -42.255 107.385 ;
        RECT -43.580 106.975 -42.255 107.145 ;
        RECT -32.700 107.035 -32.360 108.600 ;
        RECT -25.350 108.555 -23.555 108.725 ;
        RECT -49.985 106.330 -48.190 106.500 ;
        RECT -57.330 106.010 -56.990 106.235 ;
        RECT -57.330 105.840 -55.535 106.010 ;
        RECT -57.330 105.030 -56.990 105.840 ;
        RECT -48.530 105.520 -48.190 106.330 ;
        RECT -42.750 106.165 -42.255 106.975 ;
        RECT -41.400 106.515 -41.070 107.020 ;
        RECT -32.700 106.990 -32.355 107.035 ;
        RECT -32.700 106.820 -30.900 106.990 ;
        RECT -41.400 106.500 -40.450 106.515 ;
        RECT -43.580 105.995 -42.255 106.165 ;
        RECT -49.985 105.350 -48.190 105.520 ;
        RECT -57.330 104.860 -55.535 105.030 ;
        RECT -57.330 102.205 -56.990 104.860 ;
        RECT -48.530 104.540 -48.190 105.350 ;
        RECT -42.750 105.185 -42.255 105.995 ;
        RECT -43.580 105.015 -42.255 105.185 ;
        RECT -49.985 104.370 -48.190 104.540 ;
        RECT -57.330 102.035 -55.535 102.205 ;
        RECT -57.330 101.225 -56.990 102.035 ;
        RECT -48.530 101.980 -48.190 104.370 ;
        RECT -42.750 104.205 -42.255 105.015 ;
        RECT -43.580 104.035 -42.255 104.205 ;
        RECT -42.750 103.150 -42.255 104.035 ;
        RECT -41.955 106.495 -40.450 106.500 ;
        RECT -41.955 106.325 -37.490 106.495 ;
        RECT -41.955 106.290 -40.450 106.325 ;
        RECT -41.955 104.405 -41.070 106.290 ;
        RECT -32.700 106.235 -32.355 106.820 ;
        RECT -23.895 106.500 -23.555 108.555 ;
        RECT -25.350 106.330 -23.555 106.500 ;
        RECT -32.695 106.010 -32.355 106.235 ;
        RECT -32.695 105.840 -30.900 106.010 ;
        RECT -32.695 105.030 -32.355 105.840 ;
        RECT -23.895 105.520 -23.555 106.330 ;
        RECT -25.350 105.350 -23.555 105.520 ;
        RECT -32.695 104.860 -30.900 105.030 ;
        RECT -41.955 104.380 -40.455 104.405 ;
        RECT -41.955 104.210 -37.490 104.380 ;
        RECT -41.955 104.180 -40.455 104.210 ;
        RECT -41.955 104.025 -41.070 104.180 ;
        RECT -42.040 103.430 -41.070 104.025 ;
        RECT -42.040 103.400 -40.440 103.430 ;
        RECT -42.040 103.230 -37.490 103.400 ;
        RECT -42.040 103.205 -40.440 103.230 ;
        RECT -42.040 103.175 -41.070 103.205 ;
        RECT -42.040 103.150 -41.190 103.175 ;
        RECT -42.750 103.120 -41.190 103.150 ;
        RECT -44.585 102.950 -41.190 103.120 ;
        RECT -42.500 102.140 -41.190 102.950 ;
        RECT -57.330 101.055 -55.535 101.225 ;
        RECT -57.330 100.245 -56.990 101.055 ;
        RECT -57.330 100.075 -55.535 100.245 ;
        RECT -57.330 99.770 -56.990 100.075 ;
        RECT -57.330 95.145 -57.015 99.770 ;
        RECT -48.505 97.490 -48.190 101.980 ;
        RECT -44.585 101.970 -41.190 102.140 ;
        RECT -42.500 101.160 -41.190 101.970 ;
        RECT -44.585 100.990 -41.190 101.160 ;
        RECT -42.500 100.940 -41.190 100.990 ;
        RECT -42.185 100.935 -41.190 100.940 ;
        RECT -43.400 99.235 -42.905 99.475 ;
        RECT -44.730 99.065 -42.905 99.235 ;
        RECT -43.400 98.255 -42.905 99.065 ;
        RECT -44.730 98.085 -42.905 98.255 ;
        RECT -48.530 97.185 -48.190 97.490 ;
        RECT -43.400 97.655 -42.905 98.085 ;
        RECT -41.955 99.085 -41.190 100.935 ;
        RECT -40.875 102.150 -40.380 102.390 ;
        RECT -32.695 102.205 -32.355 104.860 ;
        RECT -23.895 104.540 -23.555 105.350 ;
        RECT -25.350 104.370 -23.555 104.540 ;
        RECT -40.875 101.980 -39.550 102.150 ;
        RECT -32.695 102.035 -30.900 102.205 ;
        RECT -40.875 101.170 -40.380 101.980 ;
        RECT -32.695 101.225 -32.355 102.035 ;
        RECT -23.895 101.980 -23.555 104.370 ;
        RECT -40.875 101.000 -39.550 101.170 ;
        RECT -32.695 101.055 -30.900 101.225 ;
        RECT -40.875 100.190 -40.380 101.000 ;
        RECT -32.695 100.245 -32.355 101.055 ;
        RECT -40.875 100.020 -39.550 100.190 ;
        RECT -32.695 100.075 -30.900 100.245 ;
        RECT -40.875 99.210 -40.380 100.020 ;
        RECT -32.695 99.770 -32.355 100.075 ;
        RECT -41.955 98.140 -41.120 99.085 ;
        RECT -40.875 99.040 -39.550 99.210 ;
        RECT -40.875 98.155 -40.380 99.040 ;
        RECT -41.955 97.955 -41.155 98.140 ;
        RECT -40.950 98.125 -40.380 98.155 ;
        RECT -40.950 97.955 -38.545 98.125 ;
        RECT -41.955 97.655 -41.190 97.955 ;
        RECT -43.400 97.275 -41.190 97.655 ;
        RECT -49.985 97.015 -48.190 97.185 ;
        RECT -44.730 97.105 -41.190 97.275 ;
        RECT -48.530 96.205 -48.190 97.015 ;
        RECT -43.400 96.795 -41.190 97.105 ;
        RECT -43.400 96.295 -42.905 96.795 ;
        RECT -49.985 96.035 -48.190 96.205 ;
        RECT -44.730 96.125 -42.905 96.295 ;
        RECT -48.530 95.225 -48.190 96.035 ;
        RECT -43.400 95.885 -42.905 96.125 ;
        RECT -57.345 93.535 -57.005 95.145 ;
        RECT -49.985 95.055 -48.190 95.225 ;
        RECT -57.345 93.490 -56.990 93.535 ;
        RECT -57.345 93.320 -55.535 93.490 ;
        RECT -57.345 92.510 -56.990 93.320 ;
        RECT -48.530 93.000 -48.190 95.055 ;
        RECT -49.985 92.830 -48.190 93.000 ;
        RECT -48.530 92.700 -48.190 92.830 ;
        RECT -41.955 92.700 -41.190 96.795 ;
        RECT -40.950 97.145 -40.630 97.955 ;
        RECT -40.950 96.975 -38.545 97.145 ;
        RECT -40.950 96.165 -40.630 96.975 ;
        RECT -40.950 95.995 -38.545 96.165 ;
        RECT -40.950 95.945 -40.630 95.995 ;
        RECT -32.695 95.145 -32.380 99.770 ;
        RECT -23.870 97.490 -23.555 101.980 ;
        RECT -23.895 97.185 -23.555 97.490 ;
        RECT -25.350 97.015 -23.555 97.185 ;
        RECT -23.895 96.205 -23.555 97.015 ;
        RECT -25.350 96.035 -23.555 96.205 ;
        RECT -23.895 95.225 -23.555 96.035 ;
        RECT -32.710 93.535 -32.370 95.145 ;
        RECT -25.350 95.055 -23.555 95.225 ;
        RECT -32.710 93.490 -32.355 93.535 ;
        RECT -32.710 93.320 -30.900 93.490 ;
        RECT -32.710 92.700 -32.355 93.320 ;
        RECT -23.895 93.000 -23.555 95.055 ;
        RECT -25.350 92.830 -23.555 93.000 ;
        RECT -48.530 92.510 -32.355 92.700 ;
        RECT -57.345 92.340 -55.535 92.510 ;
        RECT -48.530 92.340 -30.900 92.510 ;
        RECT -57.345 91.530 -56.990 92.340 ;
        RECT -48.530 92.020 -32.355 92.340 ;
        RECT -23.895 92.020 -23.555 92.830 ;
        RECT -49.985 91.935 -32.355 92.020 ;
        RECT -49.985 91.850 -48.190 91.935 ;
        RECT -57.345 91.360 -55.535 91.530 ;
        RECT -57.345 91.060 -56.990 91.360 ;
        RECT -57.345 90.070 -57.005 91.060 ;
        RECT -48.530 91.040 -48.190 91.850 ;
        RECT -49.985 90.870 -48.190 91.040 ;
        RECT -52.490 90.070 -51.655 90.075 ;
        RECT -48.530 90.070 -48.190 90.870 ;
        RECT -57.345 89.625 -48.190 90.070 ;
        RECT -32.710 91.530 -32.355 91.935 ;
        RECT -25.350 91.850 -23.555 92.020 ;
        RECT -32.710 91.360 -30.900 91.530 ;
        RECT -32.710 91.060 -32.355 91.360 ;
        RECT -32.710 90.070 -32.370 91.060 ;
        RECT -23.895 91.040 -23.555 91.850 ;
        RECT -25.350 90.870 -23.555 91.040 ;
        RECT -23.895 90.070 -23.555 90.870 ;
        RECT -32.710 89.625 -23.555 90.070 ;
        RECT -62.870 82.200 -62.375 82.440 ;
        RECT -63.700 82.030 -62.375 82.200 ;
        RECT -62.870 81.220 -62.375 82.030 ;
        RECT -61.520 81.570 -61.190 82.075 ;
        RECT -61.520 81.555 -60.570 81.570 ;
        RECT -63.700 81.050 -62.375 81.220 ;
        RECT -62.870 80.240 -62.375 81.050 ;
        RECT -63.700 80.070 -62.375 80.240 ;
        RECT -62.870 79.260 -62.375 80.070 ;
        RECT -63.700 79.090 -62.375 79.260 ;
        RECT -62.870 78.205 -62.375 79.090 ;
        RECT -62.075 81.550 -60.570 81.555 ;
        RECT -62.075 81.380 -57.610 81.550 ;
        RECT -62.075 81.345 -60.570 81.380 ;
        RECT -62.075 79.460 -61.190 81.345 ;
        RECT -62.075 79.435 -60.575 79.460 ;
        RECT -62.075 79.265 -57.610 79.435 ;
        RECT -62.075 79.235 -60.575 79.265 ;
        RECT -62.075 79.080 -61.190 79.235 ;
        RECT -62.160 78.485 -61.190 79.080 ;
        RECT -62.160 78.455 -60.560 78.485 ;
        RECT -62.160 78.285 -57.610 78.455 ;
        RECT -62.160 78.260 -60.560 78.285 ;
        RECT -62.160 78.230 -61.190 78.260 ;
        RECT -62.160 78.205 -61.310 78.230 ;
        RECT -62.870 78.175 -61.310 78.205 ;
        RECT -64.705 78.005 -61.310 78.175 ;
        RECT -62.620 77.195 -61.310 78.005 ;
        RECT -64.705 77.025 -61.310 77.195 ;
        RECT -62.620 76.215 -61.310 77.025 ;
        RECT -64.705 76.045 -61.310 76.215 ;
        RECT -62.620 75.995 -61.310 76.045 ;
        RECT -62.305 75.990 -61.310 75.995 ;
        RECT -63.520 74.290 -63.025 74.530 ;
        RECT -64.850 74.120 -63.025 74.290 ;
        RECT -63.520 73.310 -63.025 74.120 ;
        RECT -64.850 73.140 -63.025 73.310 ;
        RECT -63.520 72.710 -63.025 73.140 ;
        RECT -62.075 74.140 -61.310 75.990 ;
        RECT -60.995 77.205 -60.500 77.445 ;
        RECT -60.995 77.035 -59.670 77.205 ;
        RECT -60.995 76.225 -60.500 77.035 ;
        RECT -60.995 76.055 -59.670 76.225 ;
        RECT -60.995 75.245 -60.500 76.055 ;
        RECT -60.995 75.075 -59.670 75.245 ;
        RECT -60.995 74.265 -60.500 75.075 ;
        RECT -62.075 73.195 -61.240 74.140 ;
        RECT -60.995 74.095 -59.670 74.265 ;
        RECT -60.995 73.210 -60.500 74.095 ;
        RECT -62.075 73.010 -61.275 73.195 ;
        RECT -61.070 73.180 -60.500 73.210 ;
        RECT -61.070 73.010 -58.665 73.180 ;
        RECT -62.075 72.710 -61.310 73.010 ;
        RECT -63.520 72.330 -61.310 72.710 ;
        RECT -64.850 72.160 -61.310 72.330 ;
        RECT -63.520 71.850 -61.310 72.160 ;
        RECT -63.520 71.350 -63.025 71.850 ;
        RECT -64.850 71.180 -63.025 71.350 ;
        RECT -63.520 70.940 -63.025 71.180 ;
        RECT -70.300 58.600 -69.840 65.700 ;
        RECT -67.580 65.690 -67.145 65.700 ;
        RECT -62.170 65.690 -61.310 71.850 ;
        RECT -61.070 72.200 -60.750 73.010 ;
        RECT -61.070 72.030 -58.665 72.200 ;
        RECT -61.070 71.220 -60.750 72.030 ;
        RECT -61.070 71.050 -58.665 71.220 ;
        RECT -61.070 71.000 -60.750 71.050 ;
        RECT -67.580 64.830 -61.310 65.690 ;
        RECT -53.470 66.740 -53.125 66.750 ;
        RECT -52.490 66.740 -51.655 89.625 ;
        RECT -37.870 82.200 -37.375 82.440 ;
        RECT -38.700 82.030 -37.375 82.200 ;
        RECT -37.870 81.220 -37.375 82.030 ;
        RECT -36.520 81.570 -36.190 82.075 ;
        RECT -36.520 81.555 -35.570 81.570 ;
        RECT -38.700 81.050 -37.375 81.220 ;
        RECT -37.870 80.240 -37.375 81.050 ;
        RECT -38.700 80.070 -37.375 80.240 ;
        RECT -37.870 79.260 -37.375 80.070 ;
        RECT -38.700 79.090 -37.375 79.260 ;
        RECT -37.870 78.205 -37.375 79.090 ;
        RECT -37.075 81.550 -35.570 81.555 ;
        RECT -37.075 81.380 -32.610 81.550 ;
        RECT -37.075 81.345 -35.570 81.380 ;
        RECT -37.075 79.460 -36.190 81.345 ;
        RECT -37.075 79.435 -35.575 79.460 ;
        RECT -37.075 79.265 -32.610 79.435 ;
        RECT -37.075 79.235 -35.575 79.265 ;
        RECT -37.075 79.080 -36.190 79.235 ;
        RECT -37.160 78.485 -36.190 79.080 ;
        RECT -37.160 78.455 -35.560 78.485 ;
        RECT -37.160 78.285 -32.610 78.455 ;
        RECT -37.160 78.260 -35.560 78.285 ;
        RECT -37.160 78.230 -36.190 78.260 ;
        RECT -37.160 78.205 -36.310 78.230 ;
        RECT -37.870 78.175 -36.310 78.205 ;
        RECT -39.705 78.005 -36.310 78.175 ;
        RECT -37.620 77.195 -36.310 78.005 ;
        RECT -39.705 77.025 -36.310 77.195 ;
        RECT -37.620 76.215 -36.310 77.025 ;
        RECT -39.705 76.045 -36.310 76.215 ;
        RECT -37.620 75.995 -36.310 76.045 ;
        RECT -37.305 75.990 -36.310 75.995 ;
        RECT -38.520 74.290 -38.025 74.530 ;
        RECT -39.850 74.120 -38.025 74.290 ;
        RECT -38.520 73.310 -38.025 74.120 ;
        RECT -39.850 73.140 -38.025 73.310 ;
        RECT -38.520 72.710 -38.025 73.140 ;
        RECT -37.075 74.140 -36.310 75.990 ;
        RECT -35.995 77.205 -35.500 77.445 ;
        RECT -35.995 77.035 -34.670 77.205 ;
        RECT -35.995 76.225 -35.500 77.035 ;
        RECT -35.995 76.055 -34.670 76.225 ;
        RECT -35.995 75.245 -35.500 76.055 ;
        RECT -35.995 75.075 -34.670 75.245 ;
        RECT -35.995 74.265 -35.500 75.075 ;
        RECT -37.075 73.195 -36.240 74.140 ;
        RECT -35.995 74.095 -34.670 74.265 ;
        RECT -35.995 73.210 -35.500 74.095 ;
        RECT -37.075 73.010 -36.275 73.195 ;
        RECT -36.070 73.180 -35.500 73.210 ;
        RECT -36.070 73.010 -33.665 73.180 ;
        RECT -37.075 72.710 -36.310 73.010 ;
        RECT -38.520 72.330 -36.310 72.710 ;
        RECT -39.850 72.160 -36.310 72.330 ;
        RECT -38.520 71.850 -36.310 72.160 ;
        RECT -38.520 71.350 -38.025 71.850 ;
        RECT -39.850 71.180 -38.025 71.350 ;
        RECT -38.520 70.940 -38.025 71.180 ;
        RECT -37.075 71.000 -36.310 71.850 ;
        RECT -36.070 72.200 -35.750 73.010 ;
        RECT -36.070 72.030 -33.665 72.200 ;
        RECT -36.070 71.220 -35.750 72.030 ;
        RECT -36.070 71.050 -33.665 71.220 ;
        RECT -36.070 71.000 -35.750 71.050 ;
        RECT -37.075 68.875 -36.510 71.000 ;
        RECT -28.560 69.245 -28.065 69.265 ;
        RECT -27.755 69.245 -26.690 89.625 ;
        RECT -28.560 69.025 -26.690 69.245 ;
        RECT -37.505 68.825 -36.510 68.875 ;
        RECT -29.390 68.855 -26.690 69.025 ;
        RECT -38.965 68.655 -36.510 68.825 ;
        RECT -37.670 67.845 -36.510 68.655 ;
        RECT -28.560 68.045 -26.690 68.855 ;
        RECT -29.390 67.875 -26.690 68.045 ;
        RECT -38.965 67.675 -36.510 67.845 ;
        RECT -53.470 65.230 -51.655 66.740 ;
        RECT -54.135 65.190 -51.655 65.230 ;
        RECT -56.060 65.020 -51.655 65.190 ;
        RECT -37.670 65.135 -36.510 67.675 ;
        RECT -28.560 67.065 -26.690 67.875 ;
        RECT -29.390 66.895 -26.690 67.065 ;
        RECT -28.560 66.085 -26.690 66.895 ;
        RECT -29.390 65.915 -26.690 66.085 ;
        RECT -54.135 64.990 -51.655 65.020 ;
        RECT -67.580 64.820 -67.145 64.830 ;
        RECT -53.470 64.245 -51.655 64.990 ;
        RECT -38.965 64.965 -36.510 65.135 ;
        RECT -28.560 65.000 -26.690 65.915 ;
        RECT -54.105 64.210 -51.655 64.245 ;
        RECT -56.060 64.040 -51.655 64.210 ;
        RECT -37.670 64.155 -36.510 64.965 ;
        RECT -30.395 64.830 -26.690 65.000 ;
        RECT -54.105 64.005 -51.655 64.040 ;
        RECT -53.470 63.980 -51.655 64.005 ;
        RECT -38.965 63.985 -36.510 64.155 ;
        RECT -28.340 64.020 -26.690 64.830 ;
        RECT -53.330 63.975 -51.655 63.980 ;
        RECT -53.465 62.120 -53.120 62.225 ;
        RECT -52.490 62.120 -51.655 63.975 ;
        RECT -37.670 63.175 -36.510 63.985 ;
        RECT -30.395 63.850 -26.690 64.020 ;
        RECT -38.965 63.005 -36.510 63.175 ;
        RECT -28.340 63.040 -26.690 63.850 ;
        RECT -37.670 62.195 -36.510 63.005 ;
        RECT -30.395 62.870 -26.690 63.040 ;
        RECT -28.340 62.610 -26.690 62.870 ;
        RECT -53.465 60.705 -51.655 62.120 ;
        RECT -38.965 62.025 -36.510 62.195 ;
        RECT -54.130 60.665 -51.655 60.705 ;
        RECT -56.055 60.495 -51.655 60.665 ;
        RECT -54.130 60.465 -51.655 60.495 ;
        RECT -53.465 59.720 -51.655 60.465 ;
        RECT -54.100 59.685 -51.655 59.720 ;
        RECT -56.055 59.530 -51.655 59.685 ;
        RECT -37.670 59.555 -36.510 62.025 ;
        RECT -27.755 59.725 -26.690 62.610 ;
        RECT -27.825 59.675 -26.690 59.725 ;
        RECT -56.055 59.515 -53.120 59.530 ;
        RECT -54.100 59.480 -53.120 59.515 ;
        RECT -53.465 59.455 -53.120 59.480 ;
        RECT -70.300 58.430 -68.460 58.600 ;
        RECT -70.300 57.620 -69.840 58.430 ;
        RECT -53.850 57.650 -53.185 57.780 ;
        RECT -52.490 57.650 -51.655 59.530 ;
        RECT -38.105 59.315 -36.510 59.555 ;
        RECT -29.285 59.505 -26.690 59.675 ;
        RECT -38.935 59.145 -36.510 59.315 ;
        RECT -38.105 58.335 -36.510 59.145 ;
        RECT -27.825 58.695 -26.690 59.505 ;
        RECT -29.285 58.525 -26.690 58.695 ;
        RECT -27.825 58.500 -26.690 58.525 ;
        RECT -38.935 58.165 -36.510 58.335 ;
        RECT -70.300 57.450 -68.460 57.620 ;
        RECT -70.300 56.640 -69.840 57.450 ;
        RECT -70.300 56.470 -68.460 56.640 ;
        RECT -70.300 55.660 -69.840 56.470 ;
        RECT -70.300 55.490 -68.460 55.660 ;
        RECT -70.300 52.950 -69.840 55.490 ;
        RECT -53.850 54.685 -51.655 57.650 ;
        RECT -38.105 57.355 -36.510 58.165 ;
        RECT -38.935 57.185 -36.510 57.355 ;
        RECT -38.105 56.375 -36.510 57.185 ;
        RECT -38.935 56.205 -36.510 56.375 ;
        RECT -38.105 55.290 -36.510 56.205 ;
        RECT -27.755 55.985 -26.690 58.500 ;
        RECT -29.285 55.815 -26.690 55.985 ;
        RECT -39.940 55.120 -36.510 55.290 ;
        RECT -54.490 54.635 -51.655 54.685 ;
        RECT -57.410 54.465 -51.655 54.635 ;
        RECT -54.490 54.420 -51.655 54.465 ;
        RECT -53.850 53.740 -51.655 54.420 ;
        RECT -37.855 54.310 -36.510 55.120 ;
        RECT -27.805 55.005 -26.690 55.815 ;
        RECT -29.285 54.835 -26.690 55.005 ;
        RECT -39.940 54.140 -36.510 54.310 ;
        RECT -53.850 53.705 -53.185 53.740 ;
        RECT -54.410 53.655 -53.185 53.705 ;
        RECT -57.410 53.485 -53.185 53.655 ;
        RECT -54.410 53.440 -53.185 53.485 ;
        RECT -70.300 52.780 -68.460 52.950 ;
        RECT -70.300 52.690 -69.840 52.780 ;
        RECT -70.255 51.970 -69.920 52.690 ;
        RECT -70.255 51.800 -68.460 51.970 ;
        RECT -52.490 51.890 -51.655 53.740 ;
        RECT -37.855 53.330 -36.510 54.140 ;
        RECT -27.805 54.025 -26.690 54.835 ;
        RECT -29.285 53.855 -26.690 54.025 ;
        RECT -39.940 53.160 -36.510 53.330 ;
        RECT -37.855 53.110 -36.510 53.160 ;
        RECT -70.255 51.750 -69.920 51.800 ;
        RECT -37.670 46.170 -36.510 53.110 ;
        RECT -27.805 53.045 -26.690 53.855 ;
        RECT -29.285 52.875 -26.690 53.045 ;
        RECT -27.805 46.170 -26.690 52.875 ;
        RECT 72.985 51.285 79.335 51.455 ;
        RECT 72.985 51.075 73.155 51.285 ;
        RECT 72.345 49.545 73.310 51.075 ;
        RECT 79.165 50.835 79.335 51.285 ;
        RECT 77.920 50.665 79.335 50.835 ;
        RECT 72.345 49.375 74.945 49.545 ;
        RECT 72.345 49.035 73.310 49.375 ;
        RECT -37.670 44.810 -26.690 46.170 ;
        RECT 17.140 46.965 73.310 49.035 ;
        RECT 79.165 48.255 79.335 50.665 ;
        RECT 77.920 48.085 79.335 48.255 ;
        RECT 17.140 46.795 74.945 46.965 ;
        RECT 17.140 45.860 73.310 46.795 ;
        RECT 17.140 41.000 20.315 45.860 ;
        RECT 72.345 45.265 73.310 45.860 ;
        RECT 79.165 45.675 79.335 48.085 ;
        RECT 77.920 45.505 79.335 45.675 ;
        RECT 79.165 45.030 79.335 45.505 ;
        RECT 78.610 44.860 79.450 45.030 ;
        RECT 16.875 39.590 20.515 41.000 ;
        RECT 16.875 39.200 44.270 39.590 ;
        RECT 16.875 38.295 63.570 39.200 ;
        RECT 16.875 37.825 20.515 38.295 ;
        RECT 40.720 38.290 63.570 38.295 ;
        RECT -64.875 34.015 -57.020 34.715 ;
        RECT -64.875 27.790 -11.940 34.015 ;
        RECT 40.720 33.460 40.890 38.290 ;
        RECT 49.300 33.460 49.470 38.290 ;
        RECT 57.880 33.460 58.700 38.290 ;
        RECT 63.110 33.460 63.280 38.290 ;
        RECT -64.875 26.860 -57.020 27.790 ;
        RECT 119.645 21.835 305.605 23.705 ;
        RECT 119.645 21.450 493.990 21.835 ;
        RECT 79.085 20.840 81.655 20.855 ;
        RECT 119.645 20.840 121.900 21.450 ;
        RECT 74.095 18.585 121.900 20.840 ;
        RECT 74.095 18.460 76.350 18.585 ;
        RECT -66.035 16.205 76.350 18.460 ;
        RECT 106.940 17.955 108.060 18.585 ;
        RECT 105.015 17.695 111.120 17.955 ;
        RECT 101.340 17.665 103.285 17.670 ;
        RECT 105.015 17.665 105.650 17.695 ;
        RECT 98.925 17.325 105.650 17.665 ;
        RECT 107.835 17.635 110.510 17.695 ;
        RECT -66.630 11.020 -46.610 11.525 ;
        RECT -10.990 11.250 -8.735 16.205 ;
        RECT 30.055 12.130 31.770 16.205 ;
        RECT 58.740 12.430 62.750 16.205 ;
        RECT 98.970 15.870 99.140 17.325 ;
        RECT 99.950 15.870 100.120 17.325 ;
        RECT 100.930 15.870 101.100 17.325 ;
        RECT 103.220 15.870 103.390 17.325 ;
        RECT 104.200 15.870 104.370 17.325 ;
        RECT 105.180 15.870 105.350 17.325 ;
        RECT 28.620 11.870 34.725 12.130 ;
        RECT 38.110 12.100 75.300 12.430 ;
        RECT 24.945 11.840 26.890 11.845 ;
        RECT 28.620 11.840 29.255 11.870 ;
        RECT 22.530 11.500 29.255 11.840 ;
        RECT 31.440 11.810 34.115 11.870 ;
        RECT -66.735 10.690 -29.545 11.020 ;
        RECT -11.875 10.990 -5.770 11.250 ;
        RECT -15.550 10.960 -13.605 10.965 ;
        RECT -11.875 10.960 -11.240 10.990 ;
        RECT -61.795 10.330 -61.500 10.690 ;
        RECT -59.410 10.330 -59.115 10.690 ;
        RECT -58.255 10.330 -57.960 10.690 ;
        RECT -57.075 10.330 -56.780 10.690 ;
        RECT -55.885 10.330 -55.590 10.690 ;
        RECT -54.685 10.330 -54.390 10.690 ;
        RECT -53.535 10.330 -53.240 10.690 ;
        RECT -52.350 10.330 -52.055 10.690 ;
        RECT -51.180 10.330 -50.885 10.690 ;
        RECT -50.010 10.330 -49.715 10.690 ;
        RECT -46.385 10.330 -46.090 10.690 ;
        RECT -45.230 10.330 -44.935 10.690 ;
        RECT -44.050 10.330 -43.755 10.690 ;
        RECT -42.875 10.330 -42.580 10.690 ;
        RECT -41.680 10.330 -41.385 10.690 ;
        RECT -40.535 10.330 -40.240 10.690 ;
        RECT -37.505 10.330 -37.210 10.690 ;
        RECT -36.345 10.330 -36.050 10.690 ;
        RECT -35.140 10.330 -34.845 10.690 ;
        RECT -33.785 10.330 -33.490 10.690 ;
        RECT -30.845 10.330 -30.550 10.690 ;
        RECT -17.965 10.620 -11.240 10.960 ;
        RECT -9.055 10.930 -6.380 10.990 ;
        RECT -67.285 10.090 -29.525 10.330 ;
        RECT -66.455 7.855 -66.285 10.090 ;
        RECT -65.275 7.855 -65.105 10.090 ;
        RECT -64.095 7.855 -63.925 10.090 ;
        RECT -62.915 7.855 -62.745 10.090 ;
        RECT -61.735 7.855 -61.565 10.090 ;
        RECT -60.555 7.855 -60.385 10.090 ;
        RECT -59.375 7.855 -59.205 10.090 ;
        RECT -58.195 7.855 -58.025 10.090 ;
        RECT -57.015 7.855 -56.845 10.090 ;
        RECT -55.835 7.855 -55.665 10.090 ;
        RECT -54.655 7.855 -54.485 10.090 ;
        RECT -53.475 7.855 -53.305 10.090 ;
        RECT -52.295 7.855 -52.125 10.090 ;
        RECT -51.115 7.855 -50.945 10.090 ;
        RECT -49.935 7.855 -49.765 10.090 ;
        RECT -48.755 7.855 -48.585 10.090 ;
        RECT -47.515 7.855 -47.345 10.090 ;
        RECT -46.335 7.855 -46.165 10.090 ;
        RECT -45.155 7.855 -44.985 10.090 ;
        RECT -43.975 7.855 -43.805 10.090 ;
        RECT -42.795 7.855 -42.625 10.090 ;
        RECT -41.615 7.855 -41.445 10.090 ;
        RECT -40.435 7.855 -40.265 10.090 ;
        RECT -39.255 7.855 -39.085 10.090 ;
        RECT -38.075 7.855 -37.905 10.090 ;
        RECT -37.425 7.855 -37.255 10.090 ;
        RECT -36.245 7.855 -36.075 10.090 ;
        RECT -35.065 7.855 -34.895 10.090 ;
        RECT -33.885 7.855 -33.715 10.090 ;
        RECT -32.705 7.855 -32.535 10.090 ;
        RECT -32.055 7.855 -31.885 10.090 ;
        RECT -30.875 7.855 -30.705 10.090 ;
        RECT -29.695 7.855 -29.525 10.090 ;
        RECT -17.920 9.165 -17.750 10.620 ;
        RECT -16.940 9.165 -16.770 10.620 ;
        RECT -15.960 9.165 -15.790 10.620 ;
        RECT -13.670 9.165 -13.500 10.620 ;
        RECT -12.690 9.165 -12.520 10.620 ;
        RECT -11.710 9.165 -11.540 10.620 ;
        RECT -13.670 3.375 -13.500 4.830 ;
        RECT -12.690 3.375 -12.520 4.830 ;
        RECT -11.710 3.375 -11.540 4.830 ;
        RECT -13.715 3.035 -11.240 3.375 ;
        RECT -12.020 3.005 -11.240 3.035 ;
        RECT -9.055 3.005 -6.380 3.065 ;
        RECT -6.030 3.005 -5.770 10.990 ;
        RECT 22.575 10.045 22.745 11.500 ;
        RECT 23.555 10.045 23.725 11.500 ;
        RECT 24.535 10.045 24.705 11.500 ;
        RECT 26.825 10.045 26.995 11.500 ;
        RECT 27.805 10.045 27.975 11.500 ;
        RECT 28.785 10.045 28.955 11.500 ;
        RECT 3.565 7.955 3.735 9.125 ;
        RECT 2.885 7.880 3.975 7.955 ;
        RECT 5.245 7.880 5.415 9.115 ;
        RECT 2.885 7.695 5.415 7.880 ;
        RECT 6.125 7.695 6.295 9.115 ;
        RECT 7.005 7.880 7.175 9.115 ;
        RECT 8.450 7.880 8.620 9.115 ;
        RECT 9.180 7.880 9.350 9.115 ;
        RECT 12.500 7.955 12.670 9.125 ;
        RECT 14.045 7.955 14.215 9.125 ;
        RECT 12.260 7.880 14.895 7.955 ;
        RECT 7.005 7.870 14.895 7.880 ;
        RECT 17.500 7.870 19.375 8.270 ;
        RECT 7.005 7.695 19.375 7.870 ;
        RECT 2.885 6.615 19.375 7.695 ;
        RECT 2.885 6.430 5.415 6.615 ;
        RECT 2.885 6.355 3.975 6.430 ;
        RECT 3.565 5.185 3.735 6.355 ;
        RECT 5.245 5.195 5.415 6.430 ;
        RECT 6.125 5.195 6.295 6.615 ;
        RECT 7.005 6.595 19.375 6.615 ;
        RECT 7.005 6.430 14.895 6.595 ;
        RECT 7.005 5.195 7.175 6.430 ;
        RECT 8.450 5.195 8.620 6.430 ;
        RECT 9.180 5.195 9.350 6.430 ;
        RECT 12.260 6.355 14.895 6.430 ;
        RECT 17.500 6.395 19.375 6.595 ;
        RECT 12.500 5.185 12.670 6.355 ;
        RECT 14.045 5.185 14.215 6.355 ;
        RECT 26.825 4.255 26.995 5.710 ;
        RECT 27.805 4.255 27.975 5.710 ;
        RECT 28.785 4.255 28.955 5.710 ;
        RECT 26.780 3.915 29.255 4.255 ;
        RECT 28.620 3.885 29.255 3.915 ;
        RECT 31.440 3.885 34.115 3.945 ;
        RECT 34.465 3.885 34.725 11.870 ;
        RECT 39.115 11.740 39.410 12.100 ;
        RECT 42.055 11.740 42.350 12.100 ;
        RECT 43.410 11.740 43.705 12.100 ;
        RECT 44.615 11.740 44.910 12.100 ;
        RECT 45.775 11.740 46.070 12.100 ;
        RECT 48.805 11.740 49.100 12.100 ;
        RECT 49.950 11.740 50.245 12.100 ;
        RECT 51.145 11.740 51.440 12.100 ;
        RECT 52.320 11.740 52.615 12.100 ;
        RECT 53.500 11.740 53.795 12.100 ;
        RECT 54.655 11.740 54.950 12.100 ;
        RECT 58.280 11.740 58.575 12.100 ;
        RECT 59.450 11.740 59.745 12.100 ;
        RECT 60.620 11.740 60.915 12.100 ;
        RECT 61.805 11.740 62.100 12.100 ;
        RECT 62.955 11.740 63.250 12.100 ;
        RECT 64.155 11.740 64.450 12.100 ;
        RECT 65.345 11.740 65.640 12.100 ;
        RECT 66.525 11.740 66.820 12.100 ;
        RECT 67.680 11.740 67.975 12.100 ;
        RECT 70.065 11.740 70.360 12.100 ;
        RECT 38.090 11.500 75.850 11.740 ;
        RECT 38.090 9.265 38.260 11.500 ;
        RECT 39.270 9.265 39.440 11.500 ;
        RECT 40.450 9.265 40.620 11.500 ;
        RECT 41.100 9.265 41.270 11.500 ;
        RECT 42.280 9.265 42.450 11.500 ;
        RECT 43.460 9.265 43.630 11.500 ;
        RECT 44.640 9.265 44.810 11.500 ;
        RECT 45.820 9.265 45.990 11.500 ;
        RECT 46.470 9.265 46.640 11.500 ;
        RECT 47.650 9.265 47.820 11.500 ;
        RECT 48.830 9.265 49.000 11.500 ;
        RECT 50.010 9.265 50.180 11.500 ;
        RECT 51.190 9.265 51.360 11.500 ;
        RECT 52.370 9.265 52.540 11.500 ;
        RECT 53.550 9.265 53.720 11.500 ;
        RECT 54.730 9.265 54.900 11.500 ;
        RECT 55.910 9.265 56.080 11.500 ;
        RECT 57.150 9.265 57.320 11.500 ;
        RECT 58.330 9.265 58.500 11.500 ;
        RECT 59.510 9.265 59.680 11.500 ;
        RECT 60.690 9.265 60.860 11.500 ;
        RECT 61.870 9.265 62.040 11.500 ;
        RECT 63.050 9.265 63.220 11.500 ;
        RECT 64.230 9.265 64.400 11.500 ;
        RECT 65.410 9.265 65.580 11.500 ;
        RECT 66.590 9.265 66.760 11.500 ;
        RECT 67.770 9.265 67.940 11.500 ;
        RECT 68.950 9.265 69.120 11.500 ;
        RECT 70.130 9.265 70.300 11.500 ;
        RECT 71.310 9.265 71.480 11.500 ;
        RECT 72.490 9.265 72.660 11.500 ;
        RECT 73.670 9.265 73.840 11.500 ;
        RECT 74.850 9.265 75.020 11.500 ;
        RECT 103.220 10.080 103.390 11.535 ;
        RECT 104.200 10.080 104.370 11.535 ;
        RECT 105.180 10.080 105.350 11.535 ;
        RECT 103.175 9.740 105.650 10.080 ;
        RECT 105.015 9.710 105.650 9.740 ;
        RECT 107.835 9.710 110.510 9.770 ;
        RECT 110.860 9.710 111.120 17.695 ;
        RECT 255.675 16.315 258.650 21.450 ;
        RECT 266.560 16.315 269.535 21.450 ;
        RECT 276.305 16.315 279.280 21.450 ;
        RECT 288.090 16.315 291.065 21.450 ;
        RECT 209.075 15.465 221.025 16.190 ;
        RECT 254.500 15.985 291.690 16.315 ;
        RECT 255.505 15.625 255.800 15.985 ;
        RECT 258.445 15.625 258.740 15.985 ;
        RECT 259.800 15.625 260.095 15.985 ;
        RECT 261.005 15.625 261.300 15.985 ;
        RECT 262.165 15.625 262.460 15.985 ;
        RECT 265.195 15.625 265.490 15.985 ;
        RECT 266.340 15.625 266.635 15.985 ;
        RECT 267.535 15.625 267.830 15.985 ;
        RECT 268.710 15.625 269.005 15.985 ;
        RECT 269.890 15.625 270.185 15.985 ;
        RECT 271.045 15.625 271.340 15.985 ;
        RECT 274.670 15.625 274.965 15.985 ;
        RECT 275.840 15.625 276.135 15.985 ;
        RECT 277.010 15.625 277.305 15.985 ;
        RECT 278.195 15.625 278.490 15.985 ;
        RECT 279.345 15.625 279.640 15.985 ;
        RECT 280.545 15.625 280.840 15.985 ;
        RECT 281.735 15.625 282.030 15.985 ;
        RECT 282.915 15.625 283.210 15.985 ;
        RECT 284.070 15.625 284.365 15.985 ;
        RECT 286.455 15.625 286.750 15.985 ;
        RECT 209.075 15.455 226.420 15.465 ;
        RECT 207.445 15.450 226.420 15.455 ;
        RECT 195.885 15.135 226.420 15.450 ;
        RECT 195.885 15.110 202.775 15.135 ;
        RECT 207.445 15.115 216.275 15.135 ;
        RECT 220.900 15.125 226.420 15.135 ;
        RECT 209.010 15.110 216.275 15.115 ;
        RECT 222.510 15.110 224.985 15.125 ;
        RECT 133.440 14.290 134.815 14.380 ;
        RECT 133.440 13.345 140.070 14.290 ;
        RECT 195.930 13.655 196.100 15.110 ;
        RECT 196.910 13.655 197.080 15.110 ;
        RECT 197.890 13.655 198.060 15.110 ;
        RECT 200.340 13.655 200.510 15.110 ;
        RECT 201.320 13.655 201.490 15.110 ;
        RECT 202.300 13.655 202.470 15.110 ;
        RECT 209.055 13.655 209.225 15.110 ;
        RECT 210.035 13.655 210.205 15.110 ;
        RECT 211.015 13.655 211.185 15.110 ;
        RECT 213.840 13.655 214.010 15.110 ;
        RECT 214.820 13.655 214.990 15.110 ;
        RECT 215.800 13.655 215.970 15.110 ;
        RECT 222.555 13.655 222.725 15.110 ;
        RECT 223.535 13.655 223.705 15.110 ;
        RECT 224.515 13.655 224.685 15.110 ;
        RECT 133.440 13.265 134.815 13.345 ;
        RECT 139.125 11.570 140.070 13.345 ;
        RECT 140.660 11.570 145.665 11.635 ;
        RECT 105.015 9.450 111.120 9.710 ;
        RECT 138.605 11.545 145.665 11.570 ;
        RECT 138.605 11.400 147.525 11.545 ;
        RECT 164.935 11.535 169.940 11.600 ;
        RECT 138.605 10.530 138.775 11.400 ;
        RECT 140.660 11.375 147.525 11.400 ;
        RECT 140.660 11.310 145.665 11.375 ;
        RECT 141.680 10.915 141.885 11.310 ;
        RECT 143.660 10.915 143.865 11.310 ;
        RECT 147.355 10.980 147.525 11.375 ;
        RECT 141.335 10.745 145.315 10.915 ;
        RECT 138.605 10.185 139.570 10.530 ;
        RECT 28.620 3.625 34.725 3.885 ;
        RECT 28.650 3.430 31.040 3.625 ;
        RECT -12.020 2.745 -5.770 3.005 ;
        RECT -12.020 1.820 -10.375 2.745 ;
        RECT -15.960 0.175 -10.375 1.820 ;
        RECT 79.090 1.375 81.340 1.725 ;
        RECT -15.960 -0.610 -14.315 0.175 ;
        RECT -19.215 -0.870 -13.110 -0.610 ;
        RECT -22.890 -0.900 -20.945 -0.895 ;
        RECT -19.215 -0.900 -18.580 -0.870 ;
        RECT -25.305 -1.240 -18.580 -0.900 ;
        RECT -16.395 -0.930 -13.720 -0.870 ;
        RECT -25.260 -2.695 -25.090 -1.240 ;
        RECT -24.280 -2.695 -24.110 -1.240 ;
        RECT -23.300 -2.695 -23.130 -1.240 ;
        RECT -21.010 -2.695 -20.840 -1.240 ;
        RECT -20.030 -2.695 -19.860 -1.240 ;
        RECT -19.050 -2.695 -18.880 -1.240 ;
        RECT -21.010 -8.485 -20.840 -7.030 ;
        RECT -20.030 -8.485 -19.860 -7.030 ;
        RECT -19.050 -8.485 -18.880 -7.030 ;
        RECT -21.055 -8.825 -18.580 -8.485 ;
        RECT -19.215 -8.855 -18.580 -8.825 ;
        RECT -16.395 -8.855 -13.720 -8.795 ;
        RECT -13.370 -8.855 -13.110 -0.870 ;
        RECT 29.285 -0.880 81.340 1.375 ;
        RECT 106.440 1.205 107.705 9.450 ;
        RECT 109.575 1.205 110.335 9.450 ;
        RECT 138.605 7.320 138.775 10.185 ;
        RECT 139.395 7.320 139.565 10.185 ;
        RECT 141.335 9.265 141.505 10.745 ;
        RECT 142.915 9.265 143.085 10.745 ;
        RECT 145.145 9.290 145.315 10.745 ;
        RECT 146.795 10.615 147.525 10.980 ;
        RECT 146.565 9.290 146.735 10.330 ;
        RECT 147.355 9.290 147.525 10.615 ;
        RECT 162.880 11.510 169.940 11.535 ;
        RECT 162.880 11.365 171.800 11.510 ;
        RECT 162.880 10.495 163.050 11.365 ;
        RECT 164.935 11.340 171.800 11.365 ;
        RECT 164.935 11.275 169.940 11.340 ;
        RECT 165.955 10.880 166.160 11.275 ;
        RECT 167.935 10.880 168.140 11.275 ;
        RECT 171.630 10.945 171.800 11.340 ;
        RECT 165.610 10.710 169.590 10.880 ;
        RECT 162.880 10.150 163.845 10.495 ;
        RECT 141.335 7.320 141.505 8.360 ;
        RECT 142.915 7.320 143.085 8.360 ;
        RECT 145.145 7.320 145.315 8.360 ;
        RECT 146.585 7.315 146.755 8.355 ;
        RECT 147.375 7.315 147.545 8.355 ;
        RECT 151.650 6.430 151.820 9.220 ;
        RECT 153.230 6.430 153.400 9.220 ;
        RECT 154.810 6.430 154.980 9.220 ;
        RECT 156.390 6.430 156.560 9.220 ;
        RECT 157.970 6.430 158.140 9.220 ;
        RECT 162.880 7.285 163.050 10.150 ;
        RECT 163.670 7.285 163.840 10.150 ;
        RECT 165.610 9.230 165.780 10.710 ;
        RECT 167.190 9.230 167.360 10.710 ;
        RECT 169.420 9.255 169.590 10.710 ;
        RECT 171.070 10.580 171.800 10.945 ;
        RECT 170.840 9.255 171.010 10.295 ;
        RECT 171.630 9.255 171.800 10.580 ;
        RECT 165.610 7.285 165.780 8.325 ;
        RECT 167.190 7.285 167.360 8.325 ;
        RECT 169.420 7.285 169.590 8.325 ;
        RECT 170.860 7.280 171.030 8.320 ;
        RECT 171.650 7.280 171.820 8.320 ;
        RECT 175.325 6.540 175.495 9.330 ;
        RECT 176.905 6.540 177.075 9.330 ;
        RECT 178.485 6.540 178.655 9.330 ;
        RECT 180.065 6.540 180.235 9.330 ;
        RECT 181.645 6.815 181.815 9.330 ;
        RECT 183.930 6.815 184.100 9.115 ;
        RECT 181.645 6.540 184.100 6.815 ;
        RECT 151.605 5.895 158.140 6.430 ;
        RECT 175.280 6.495 184.100 6.540 ;
        RECT 175.280 6.005 181.815 6.495 ;
        RECT 183.930 6.325 184.100 6.495 ;
        RECT 185.510 6.325 185.680 9.115 ;
        RECT 187.090 6.325 187.260 9.115 ;
        RECT 188.670 6.325 188.840 9.115 ;
        RECT 190.250 6.630 190.420 9.115 ;
        RECT 205.360 6.650 205.530 8.105 ;
        RECT 206.340 6.650 206.510 8.105 ;
        RECT 207.320 6.650 207.490 8.105 ;
        RECT 209.545 6.650 209.715 8.105 ;
        RECT 210.525 6.650 210.695 8.105 ;
        RECT 211.505 6.650 211.675 8.105 ;
        RECT 218.860 6.650 219.030 8.105 ;
        RECT 219.840 6.650 220.010 8.105 ;
        RECT 220.820 6.650 220.990 8.105 ;
        RECT 223.045 6.650 223.215 8.105 ;
        RECT 224.025 6.650 224.195 8.105 ;
        RECT 225.005 6.650 225.175 8.105 ;
        RECT 225.975 7.360 226.420 15.125 ;
        RECT 254.480 15.385 292.240 15.625 ;
        RECT 254.480 13.150 254.650 15.385 ;
        RECT 255.660 13.150 255.830 15.385 ;
        RECT 256.840 13.150 257.010 15.385 ;
        RECT 257.490 13.150 257.660 15.385 ;
        RECT 258.670 13.150 258.840 15.385 ;
        RECT 259.850 13.150 260.020 15.385 ;
        RECT 261.030 13.150 261.200 15.385 ;
        RECT 262.210 13.150 262.380 15.385 ;
        RECT 262.860 13.150 263.030 15.385 ;
        RECT 264.040 13.150 264.210 15.385 ;
        RECT 265.220 13.150 265.390 15.385 ;
        RECT 266.400 13.150 266.570 15.385 ;
        RECT 267.580 13.150 267.750 15.385 ;
        RECT 268.760 13.150 268.930 15.385 ;
        RECT 269.940 13.150 270.110 15.385 ;
        RECT 271.120 13.150 271.290 15.385 ;
        RECT 272.300 13.150 272.470 15.385 ;
        RECT 273.540 13.150 273.710 15.385 ;
        RECT 274.720 13.150 274.890 15.385 ;
        RECT 275.900 13.150 276.070 15.385 ;
        RECT 277.080 13.150 277.250 15.385 ;
        RECT 278.260 13.150 278.430 15.385 ;
        RECT 279.440 13.150 279.610 15.385 ;
        RECT 280.620 13.150 280.790 15.385 ;
        RECT 281.800 13.150 281.970 15.385 ;
        RECT 282.980 13.150 283.150 15.385 ;
        RECT 284.160 13.150 284.330 15.385 ;
        RECT 285.340 13.150 285.510 15.385 ;
        RECT 286.520 13.150 286.690 15.385 ;
        RECT 287.700 13.150 287.870 15.385 ;
        RECT 288.880 13.150 289.050 15.385 ;
        RECT 290.060 13.150 290.230 15.385 ;
        RECT 291.240 13.150 291.410 15.385 ;
        RECT 227.895 7.360 228.065 8.555 ;
        RECT 225.975 7.100 228.065 7.360 ;
        RECT 228.875 7.100 229.045 8.555 ;
        RECT 229.855 7.100 230.025 8.555 ;
        RECT 225.975 7.075 230.325 7.100 ;
        RECT 225.975 6.650 226.420 7.075 ;
        RECT 227.850 6.760 230.325 7.075 ;
        RECT 303.350 6.990 493.990 21.450 ;
        RECT 190.245 6.625 200.490 6.630 ;
        RECT 205.055 6.625 214.065 6.650 ;
        RECT 218.555 6.625 226.420 6.650 ;
        RECT 190.245 6.325 226.420 6.625 ;
        RECT 303.350 6.550 305.605 6.990 ;
        RECT 175.325 5.620 175.495 6.005 ;
        RECT 176.905 5.620 177.075 6.005 ;
        RECT 178.485 5.620 178.655 6.005 ;
        RECT 180.065 5.620 180.235 6.005 ;
        RECT 181.645 5.620 181.815 6.005 ;
        RECT 151.605 4.970 158.140 5.505 ;
        RECT 175.280 5.085 181.815 5.620 ;
        RECT 183.885 6.310 226.420 6.325 ;
        RECT 183.885 6.210 200.490 6.310 ;
        RECT 183.885 5.300 190.420 6.210 ;
        RECT 151.650 2.180 151.820 4.970 ;
        RECT 153.230 2.180 153.400 4.970 ;
        RECT 154.810 2.180 154.980 4.970 ;
        RECT 156.390 2.180 156.560 4.970 ;
        RECT 157.970 2.180 158.140 4.970 ;
        RECT 175.325 2.295 175.495 5.085 ;
        RECT 176.905 2.295 177.075 5.085 ;
        RECT 178.485 2.295 178.655 5.085 ;
        RECT 180.065 2.295 180.235 5.085 ;
        RECT 181.645 5.055 181.815 5.085 ;
        RECT 183.930 5.055 184.100 5.300 ;
        RECT 181.645 4.735 184.100 5.055 ;
        RECT 181.645 2.295 181.815 4.735 ;
        RECT 183.930 2.510 184.100 4.735 ;
        RECT 185.510 2.510 185.680 5.300 ;
        RECT 187.090 2.510 187.260 5.300 ;
        RECT 188.670 2.510 188.840 5.300 ;
        RECT 190.250 2.510 190.420 5.300 ;
        RECT 266.810 4.295 322.665 6.550 ;
        RECT 266.810 1.760 270.000 4.295 ;
        RECT 273.795 1.760 276.985 4.295 ;
        RECT 280.865 1.760 284.055 4.295 ;
        RECT 286.295 1.760 289.485 4.295 ;
        RECT 253.485 1.430 290.675 1.760 ;
        RECT 105.875 0.945 111.980 1.205 ;
        RECT 254.490 1.070 254.785 1.430 ;
        RECT 257.430 1.070 257.725 1.430 ;
        RECT 258.785 1.070 259.080 1.430 ;
        RECT 259.990 1.070 260.285 1.430 ;
        RECT 261.150 1.070 261.445 1.430 ;
        RECT 264.180 1.070 264.475 1.430 ;
        RECT 265.325 1.070 265.620 1.430 ;
        RECT 266.520 1.070 266.815 1.430 ;
        RECT 267.695 1.070 267.990 1.430 ;
        RECT 268.875 1.070 269.170 1.430 ;
        RECT 270.030 1.070 270.325 1.430 ;
        RECT 273.655 1.070 273.950 1.430 ;
        RECT 274.825 1.070 275.120 1.430 ;
        RECT 275.995 1.070 276.290 1.430 ;
        RECT 277.180 1.070 277.475 1.430 ;
        RECT 278.330 1.070 278.625 1.430 ;
        RECT 279.530 1.070 279.825 1.430 ;
        RECT 280.720 1.070 281.015 1.430 ;
        RECT 281.900 1.070 282.195 1.430 ;
        RECT 283.055 1.070 283.350 1.430 ;
        RECT 285.440 1.070 285.735 1.430 ;
        RECT 102.200 0.915 104.145 0.920 ;
        RECT 105.875 0.915 106.510 0.945 ;
        RECT 99.785 0.575 106.510 0.915 ;
        RECT 108.695 0.885 111.370 0.945 ;
        RECT 99.830 -0.880 100.000 0.575 ;
        RECT 100.810 -0.880 100.980 0.575 ;
        RECT 101.790 -0.880 101.960 0.575 ;
        RECT 104.080 -0.880 104.250 0.575 ;
        RECT 105.060 -0.880 105.230 0.575 ;
        RECT 106.040 -0.880 106.210 0.575 ;
        RECT 29.385 -1.320 31.055 -0.880 ;
        RECT 28.695 -1.580 34.800 -1.320 ;
        RECT 41.515 -1.350 43.770 -0.880 ;
        RECT 49.455 -1.350 51.710 -0.880 ;
        RECT 57.160 -1.350 59.415 -0.880 ;
        RECT 63.250 -1.350 65.505 -0.880 ;
        RECT 69.240 -1.350 71.495 -0.880 ;
        RECT 79.090 -1.045 81.340 -0.880 ;
        RECT 25.020 -1.610 26.965 -1.605 ;
        RECT 28.695 -1.610 29.330 -1.580 ;
        RECT 22.605 -1.950 29.330 -1.610 ;
        RECT 31.515 -1.640 34.190 -1.580 ;
        RECT 22.650 -3.405 22.820 -1.950 ;
        RECT 23.630 -3.405 23.800 -1.950 ;
        RECT 24.610 -3.405 24.780 -1.950 ;
        RECT 26.900 -3.405 27.070 -1.950 ;
        RECT 27.880 -3.405 28.050 -1.950 ;
        RECT 28.860 -3.405 29.030 -1.950 ;
        RECT -19.215 -9.115 -13.110 -8.855 ;
        RECT 26.900 -9.195 27.070 -7.740 ;
        RECT 27.880 -9.195 28.050 -7.740 ;
        RECT 28.860 -9.195 29.030 -7.740 ;
        RECT 26.855 -9.535 29.330 -9.195 ;
        RECT 28.695 -9.565 29.330 -9.535 ;
        RECT 31.515 -9.565 34.190 -9.505 ;
        RECT 34.540 -9.565 34.800 -1.580 ;
        RECT 37.905 -1.680 75.095 -1.350 ;
        RECT 38.910 -2.040 39.205 -1.680 ;
        RECT 41.850 -2.040 42.145 -1.680 ;
        RECT 43.205 -2.040 43.500 -1.680 ;
        RECT 44.410 -2.040 44.705 -1.680 ;
        RECT 45.570 -2.040 45.865 -1.680 ;
        RECT 48.600 -2.040 48.895 -1.680 ;
        RECT 49.745 -2.040 50.040 -1.680 ;
        RECT 50.940 -2.040 51.235 -1.680 ;
        RECT 52.115 -2.040 52.410 -1.680 ;
        RECT 53.295 -2.040 53.590 -1.680 ;
        RECT 54.450 -2.040 54.745 -1.680 ;
        RECT 58.075 -2.040 58.370 -1.680 ;
        RECT 59.245 -2.040 59.540 -1.680 ;
        RECT 60.415 -2.040 60.710 -1.680 ;
        RECT 61.600 -2.040 61.895 -1.680 ;
        RECT 62.750 -2.040 63.045 -1.680 ;
        RECT 63.950 -2.040 64.245 -1.680 ;
        RECT 65.140 -2.040 65.435 -1.680 ;
        RECT 66.320 -2.040 66.615 -1.680 ;
        RECT 67.475 -2.040 67.770 -1.680 ;
        RECT 69.860 -2.040 70.155 -1.680 ;
        RECT 37.885 -2.280 75.645 -2.040 ;
        RECT 37.885 -4.515 38.055 -2.280 ;
        RECT 39.065 -4.515 39.235 -2.280 ;
        RECT 40.245 -4.515 40.415 -2.280 ;
        RECT 40.895 -4.515 41.065 -2.280 ;
        RECT 42.075 -4.515 42.245 -2.280 ;
        RECT 43.255 -4.515 43.425 -2.280 ;
        RECT 44.435 -4.515 44.605 -2.280 ;
        RECT 45.615 -4.515 45.785 -2.280 ;
        RECT 46.265 -4.515 46.435 -2.280 ;
        RECT 47.445 -4.515 47.615 -2.280 ;
        RECT 48.625 -4.515 48.795 -2.280 ;
        RECT 49.805 -4.515 49.975 -2.280 ;
        RECT 50.985 -4.515 51.155 -2.280 ;
        RECT 52.165 -4.515 52.335 -2.280 ;
        RECT 53.345 -4.515 53.515 -2.280 ;
        RECT 54.525 -4.515 54.695 -2.280 ;
        RECT 55.705 -4.515 55.875 -2.280 ;
        RECT 56.945 -4.515 57.115 -2.280 ;
        RECT 58.125 -4.515 58.295 -2.280 ;
        RECT 59.305 -4.515 59.475 -2.280 ;
        RECT 60.485 -4.515 60.655 -2.280 ;
        RECT 61.665 -4.515 61.835 -2.280 ;
        RECT 62.845 -4.515 63.015 -2.280 ;
        RECT 64.025 -4.515 64.195 -2.280 ;
        RECT 65.205 -4.515 65.375 -2.280 ;
        RECT 66.385 -4.515 66.555 -2.280 ;
        RECT 67.565 -4.515 67.735 -2.280 ;
        RECT 68.745 -4.515 68.915 -2.280 ;
        RECT 69.925 -4.515 70.095 -2.280 ;
        RECT 71.105 -4.515 71.275 -2.280 ;
        RECT 72.285 -4.515 72.455 -2.280 ;
        RECT 73.465 -4.515 73.635 -2.280 ;
        RECT 74.645 -4.515 74.815 -2.280 ;
        RECT 104.080 -6.670 104.250 -5.215 ;
        RECT 105.060 -6.670 105.230 -5.215 ;
        RECT 106.040 -6.670 106.210 -5.215 ;
        RECT 104.035 -7.010 106.510 -6.670 ;
        RECT 105.875 -7.040 106.510 -7.010 ;
        RECT 108.695 -7.040 111.370 -6.980 ;
        RECT 111.720 -7.040 111.980 0.945 ;
        RECT 253.465 0.830 291.225 1.070 ;
        RECT 134.940 -0.345 136.520 -0.190 ;
        RECT 138.835 -0.345 139.600 -0.295 ;
        RECT 134.425 -0.745 136.520 -0.345 ;
        RECT 138.025 -0.665 139.600 -0.345 ;
        RECT 163.110 -0.360 163.875 -0.330 ;
        RECT 138.025 -0.745 138.835 -0.665 ;
        RECT 162.305 -0.700 163.875 -0.360 ;
        RECT 134.940 -0.830 136.520 -0.745 ;
        RECT 162.305 -0.760 163.115 -0.700 ;
        RECT 253.465 -1.405 253.635 0.830 ;
        RECT 254.645 -1.405 254.815 0.830 ;
        RECT 255.825 -1.405 255.995 0.830 ;
        RECT 256.475 -1.405 256.645 0.830 ;
        RECT 257.655 -1.405 257.825 0.830 ;
        RECT 258.835 -1.405 259.005 0.830 ;
        RECT 260.015 -1.405 260.185 0.830 ;
        RECT 261.195 -1.405 261.365 0.830 ;
        RECT 261.845 -1.405 262.015 0.830 ;
        RECT 263.025 -1.405 263.195 0.830 ;
        RECT 264.205 -1.405 264.375 0.830 ;
        RECT 265.385 -1.405 265.555 0.830 ;
        RECT 266.565 -1.405 266.735 0.830 ;
        RECT 267.745 -1.405 267.915 0.830 ;
        RECT 268.925 -1.405 269.095 0.830 ;
        RECT 270.105 -1.405 270.275 0.830 ;
        RECT 271.285 -1.405 271.455 0.830 ;
        RECT 272.525 -1.405 272.695 0.830 ;
        RECT 273.705 -1.405 273.875 0.830 ;
        RECT 274.885 -1.405 275.055 0.830 ;
        RECT 276.065 -1.405 276.235 0.830 ;
        RECT 277.245 -1.405 277.415 0.830 ;
        RECT 278.425 -1.405 278.595 0.830 ;
        RECT 279.605 -1.405 279.775 0.830 ;
        RECT 280.785 -1.405 280.955 0.830 ;
        RECT 281.965 -1.405 282.135 0.830 ;
        RECT 283.145 -1.405 283.315 0.830 ;
        RECT 284.325 -1.405 284.495 0.830 ;
        RECT 285.505 -1.405 285.675 0.830 ;
        RECT 286.685 -1.405 286.855 0.830 ;
        RECT 287.865 -1.405 288.035 0.830 ;
        RECT 289.045 -1.405 289.215 0.830 ;
        RECT 290.225 -1.405 290.395 0.830 ;
        RECT 105.875 -7.300 111.980 -7.040 ;
        RECT 276.660 -7.585 278.915 -7.580 ;
        RECT 283.345 -7.585 285.600 -7.580 ;
        RECT 289.280 -7.585 291.535 -7.580 ;
        RECT 320.410 -7.585 322.665 4.295 ;
        RECT 28.695 -9.825 34.800 -9.565 ;
        RECT 269.460 -9.840 322.665 -7.585 ;
        RECT 269.460 -13.475 271.715 -9.840 ;
        RECT 276.660 -13.475 278.915 -9.840 ;
        RECT 283.345 -13.475 285.600 -9.840 ;
        RECT 289.280 -13.475 291.535 -9.840 ;
        RECT 320.410 -13.125 322.665 -9.840 ;
        RECT 318.010 -13.385 324.115 -13.125 ;
        RECT 314.335 -13.415 316.280 -13.410 ;
        RECT 318.010 -13.415 318.645 -13.385 ;
        RECT 253.485 -13.655 291.535 -13.475 ;
        RECT 253.485 -13.805 290.675 -13.655 ;
        RECT 311.920 -13.755 318.645 -13.415 ;
        RECT 320.830 -13.445 323.505 -13.385 ;
        RECT 254.490 -14.165 254.785 -13.805 ;
        RECT 257.430 -14.165 257.725 -13.805 ;
        RECT 258.785 -14.165 259.080 -13.805 ;
        RECT 259.990 -14.165 260.285 -13.805 ;
        RECT 261.150 -14.165 261.445 -13.805 ;
        RECT 264.180 -14.165 264.475 -13.805 ;
        RECT 265.325 -14.165 265.620 -13.805 ;
        RECT 266.520 -14.165 266.815 -13.805 ;
        RECT 267.695 -14.165 267.990 -13.805 ;
        RECT 268.875 -14.165 269.170 -13.805 ;
        RECT 270.030 -14.165 270.325 -13.805 ;
        RECT 273.655 -14.165 273.950 -13.805 ;
        RECT 274.825 -14.165 275.120 -13.805 ;
        RECT 275.995 -14.165 276.290 -13.805 ;
        RECT 277.180 -14.165 277.475 -13.805 ;
        RECT 278.330 -14.165 278.625 -13.805 ;
        RECT 279.530 -14.165 279.825 -13.805 ;
        RECT 280.720 -14.165 281.015 -13.805 ;
        RECT 281.900 -14.165 282.195 -13.805 ;
        RECT 283.055 -14.165 283.350 -13.805 ;
        RECT 285.440 -14.165 285.735 -13.805 ;
        RECT 253.465 -14.405 291.225 -14.165 ;
        RECT 253.465 -16.640 253.635 -14.405 ;
        RECT 254.645 -16.640 254.815 -14.405 ;
        RECT 255.825 -16.640 255.995 -14.405 ;
        RECT 256.475 -16.640 256.645 -14.405 ;
        RECT 257.655 -16.640 257.825 -14.405 ;
        RECT 258.835 -16.640 259.005 -14.405 ;
        RECT 260.015 -16.640 260.185 -14.405 ;
        RECT 261.195 -16.640 261.365 -14.405 ;
        RECT 261.845 -16.640 262.015 -14.405 ;
        RECT 263.025 -16.640 263.195 -14.405 ;
        RECT 264.205 -16.640 264.375 -14.405 ;
        RECT 265.385 -16.640 265.555 -14.405 ;
        RECT 266.565 -16.640 266.735 -14.405 ;
        RECT 267.745 -16.640 267.915 -14.405 ;
        RECT 268.925 -16.640 269.095 -14.405 ;
        RECT 270.105 -16.640 270.275 -14.405 ;
        RECT 271.285 -16.640 271.455 -14.405 ;
        RECT 272.525 -16.640 272.695 -14.405 ;
        RECT 273.705 -16.640 273.875 -14.405 ;
        RECT 274.885 -16.640 275.055 -14.405 ;
        RECT 276.065 -16.640 276.235 -14.405 ;
        RECT 277.245 -16.640 277.415 -14.405 ;
        RECT 278.425 -16.640 278.595 -14.405 ;
        RECT 279.605 -16.640 279.775 -14.405 ;
        RECT 280.785 -16.640 280.955 -14.405 ;
        RECT 281.965 -16.640 282.135 -14.405 ;
        RECT 283.145 -16.640 283.315 -14.405 ;
        RECT 284.325 -16.640 284.495 -14.405 ;
        RECT 285.505 -16.640 285.675 -14.405 ;
        RECT 286.685 -16.640 286.855 -14.405 ;
        RECT 287.865 -16.640 288.035 -14.405 ;
        RECT 289.045 -16.640 289.215 -14.405 ;
        RECT 290.225 -16.640 290.395 -14.405 ;
        RECT 311.965 -15.210 312.135 -13.755 ;
        RECT 312.945 -15.210 313.115 -13.755 ;
        RECT 313.925 -15.210 314.095 -13.755 ;
        RECT 316.215 -15.210 316.385 -13.755 ;
        RECT 317.195 -15.210 317.365 -13.755 ;
        RECT 318.175 -15.210 318.345 -13.755 ;
        RECT 316.215 -21.000 316.385 -19.545 ;
        RECT 317.195 -21.000 317.365 -19.545 ;
        RECT 318.175 -21.000 318.345 -19.545 ;
        RECT 316.170 -21.340 318.645 -21.000 ;
        RECT 318.010 -21.370 318.645 -21.340 ;
        RECT 320.830 -21.370 323.505 -21.310 ;
        RECT 323.855 -21.370 324.115 -13.385 ;
        RECT 318.010 -21.630 324.115 -21.370 ;
        RECT 479.145 -23.490 493.990 6.990 ;
        RECT 478.715 -38.335 493.990 -23.490 ;
        RECT 479.145 -63.340 493.990 -38.335 ;
        RECT 406.890 -79.080 493.990 -63.340 ;
        RECT 406.890 -80.290 422.630 -79.080 ;
        RECT -74.655 -82.895 -74.485 -80.660 ;
        RECT -73.475 -82.895 -73.305 -80.660 ;
        RECT -72.295 -82.895 -72.125 -80.660 ;
        RECT -71.115 -82.895 -70.945 -80.660 ;
        RECT -69.935 -82.895 -69.765 -80.660 ;
        RECT -68.755 -82.895 -68.585 -80.660 ;
        RECT -67.575 -82.895 -67.405 -80.660 ;
        RECT -66.395 -82.895 -66.225 -80.660 ;
        RECT -65.215 -82.895 -65.045 -80.660 ;
        RECT -64.035 -82.895 -63.865 -80.660 ;
        RECT -62.855 -82.895 -62.685 -80.660 ;
        RECT -61.675 -82.895 -61.505 -80.660 ;
        RECT -60.495 -82.895 -60.325 -80.660 ;
        RECT -59.315 -82.895 -59.145 -80.660 ;
        RECT -58.135 -82.895 -57.965 -80.660 ;
        RECT -56.955 -82.895 -56.785 -80.660 ;
        RECT -55.715 -82.895 -55.545 -80.660 ;
        RECT -54.535 -82.895 -54.365 -80.660 ;
        RECT -53.355 -82.895 -53.185 -80.660 ;
        RECT -52.175 -82.895 -52.005 -80.660 ;
        RECT -50.995 -82.895 -50.825 -80.660 ;
        RECT -49.815 -82.895 -49.645 -80.660 ;
        RECT -48.635 -82.895 -48.465 -80.660 ;
        RECT -47.455 -82.895 -47.285 -80.660 ;
        RECT -46.275 -82.895 -46.105 -80.660 ;
        RECT -45.625 -82.895 -45.455 -80.660 ;
        RECT -44.445 -82.895 -44.275 -80.660 ;
        RECT -43.265 -82.895 -43.095 -80.660 ;
        RECT -42.085 -82.895 -41.915 -80.660 ;
        RECT -40.905 -82.895 -40.735 -80.660 ;
        RECT -40.255 -82.895 -40.085 -80.660 ;
        RECT -39.075 -82.895 -38.905 -80.660 ;
        RECT -37.895 -82.895 -37.725 -80.660 ;
        RECT 126.125 -81.395 431.865 -80.290 ;
        RECT -75.485 -83.135 -37.725 -82.895 ;
        RECT -69.995 -83.495 -69.700 -83.135 ;
        RECT -67.610 -83.495 -67.315 -83.135 ;
        RECT -66.455 -83.495 -66.160 -83.135 ;
        RECT -65.275 -83.495 -64.980 -83.135 ;
        RECT -64.085 -83.495 -63.790 -83.135 ;
        RECT -62.885 -83.495 -62.590 -83.135 ;
        RECT -61.735 -83.495 -61.440 -83.135 ;
        RECT -60.550 -83.495 -60.255 -83.135 ;
        RECT -59.380 -83.495 -59.085 -83.135 ;
        RECT -58.210 -83.495 -57.915 -83.135 ;
        RECT -54.585 -83.495 -54.290 -83.135 ;
        RECT -53.430 -83.495 -53.135 -83.135 ;
        RECT -52.250 -83.495 -51.955 -83.135 ;
        RECT -51.075 -83.495 -50.780 -83.135 ;
        RECT -49.880 -83.495 -49.585 -83.135 ;
        RECT -48.735 -83.495 -48.440 -83.135 ;
        RECT -45.705 -83.495 -45.410 -83.135 ;
        RECT -44.545 -83.495 -44.250 -83.135 ;
        RECT -43.340 -83.495 -43.045 -83.135 ;
        RECT -41.985 -83.495 -41.690 -83.135 ;
        RECT -39.045 -83.495 -38.750 -83.135 ;
        RECT -74.935 -83.825 -37.745 -83.495 ;
        RECT -70.530 -91.210 -68.780 -83.825 ;
        RECT -59.415 -91.210 -57.665 -83.825 ;
        RECT -49.050 -91.030 -47.050 -83.825 ;
        RECT 30.985 -85.205 431.865 -81.395 ;
        RECT 30.985 -90.975 34.795 -85.205 ;
        RECT 126.125 -85.805 431.865 -85.205 ;
        RECT -40.160 -91.030 37.140 -90.975 ;
        RECT -51.815 -91.210 37.140 -91.030 ;
        RECT -76.940 -91.475 37.140 -91.210 ;
        RECT -76.940 -91.525 -50.815 -91.475 ;
        RECT -76.940 -91.550 -69.075 -91.525 ;
        RECT -64.585 -91.550 -55.575 -91.525 ;
        RECT -76.940 -94.345 -76.495 -91.550 ;
        RECT -75.695 -93.005 -75.525 -91.550 ;
        RECT -74.715 -93.005 -74.545 -91.550 ;
        RECT -73.735 -93.005 -73.565 -91.550 ;
        RECT -71.510 -93.005 -71.340 -91.550 ;
        RECT -70.530 -93.005 -70.360 -91.550 ;
        RECT -69.550 -93.005 -69.380 -91.550 ;
        RECT -62.195 -93.005 -62.025 -91.550 ;
        RECT -61.215 -93.005 -61.045 -91.550 ;
        RECT -60.235 -93.005 -60.065 -91.550 ;
        RECT -58.010 -93.005 -57.840 -91.550 ;
        RECT -57.030 -93.005 -56.860 -91.550 ;
        RECT -56.050 -93.005 -55.880 -91.550 ;
        RECT -43.905 -92.095 -43.680 -91.475 ;
        RECT -41.795 -92.090 -41.570 -91.475 ;
        RECT -121.755 -95.410 -76.495 -94.345 ;
        RECT -43.885 -95.055 -43.715 -92.095 ;
        RECT -41.770 -95.055 -41.600 -92.090 ;
        RECT -40.820 -92.105 -40.595 -91.475 ;
        RECT -40.170 -91.940 37.140 -91.475 ;
        RECT -40.790 -95.055 -40.620 -92.105 ;
        RECT -33.345 -92.475 -28.085 -91.940 ;
        RECT -33.345 -93.120 -33.145 -92.475 ;
        RECT -32.400 -93.120 -32.170 -92.475 ;
        RECT -31.410 -93.100 -31.180 -92.475 ;
        RECT -33.345 -94.035 -33.175 -93.120 ;
        RECT -32.365 -94.035 -32.195 -93.120 ;
        RECT -31.385 -94.035 -31.215 -93.100 ;
        RECT -30.845 -93.120 -30.615 -92.475 ;
        RECT -29.865 -93.095 -29.635 -92.475 ;
        RECT -30.815 -94.035 -30.645 -93.120 ;
        RECT -29.835 -94.035 -29.665 -93.095 ;
        RECT -29.300 -93.145 -29.070 -92.475 ;
        RECT -28.315 -93.085 -28.085 -92.475 ;
        RECT -29.270 -94.035 -29.100 -93.145 ;
        RECT -28.290 -94.035 -28.120 -93.085 ;
        RECT -121.755 -95.460 -110.580 -95.410 ;
        RECT -121.755 -104.165 -120.395 -95.460 ;
        RECT -113.690 -96.940 -113.520 -95.460 ;
        RECT -112.710 -96.940 -112.540 -95.460 ;
        RECT -111.730 -96.940 -111.560 -95.460 ;
        RECT -110.750 -96.940 -110.580 -95.460 ;
        RECT -108.065 -95.480 -106.840 -95.410 ;
        RECT -108.040 -96.940 -107.870 -95.480 ;
        RECT -107.060 -96.940 -106.890 -95.480 ;
        RECT -103.955 -95.720 -97.320 -95.410 ;
        RECT -103.955 -95.995 -97.300 -95.720 ;
        RECT -103.695 -98.050 -103.525 -95.995 ;
        RECT -102.715 -98.050 -102.545 -95.995 ;
        RECT -101.735 -96.215 -97.300 -95.995 ;
        RECT -101.735 -98.050 -101.565 -96.215 ;
        RECT -100.650 -97.045 -100.480 -96.215 ;
        RECT -99.670 -97.045 -99.500 -96.215 ;
        RECT -98.690 -97.045 -98.520 -96.215 ;
        RECT -97.710 -97.045 -97.540 -96.215 ;
        RECT -76.940 -100.025 -76.495 -95.410 ;
        RECT -26.710 -96.125 -26.135 -91.940 ;
        RECT -19.275 -92.130 -16.310 -91.940 ;
        RECT -20.845 -92.475 -15.585 -92.130 ;
        RECT -20.845 -93.120 -20.645 -92.475 ;
        RECT -19.900 -93.120 -19.670 -92.475 ;
        RECT -18.910 -93.100 -18.680 -92.475 ;
        RECT -20.845 -94.035 -20.675 -93.120 ;
        RECT -19.865 -94.035 -19.695 -93.120 ;
        RECT -18.885 -94.035 -18.715 -93.100 ;
        RECT -18.345 -93.120 -18.115 -92.475 ;
        RECT -17.365 -93.095 -17.135 -92.475 ;
        RECT -18.315 -94.035 -18.145 -93.120 ;
        RECT -17.335 -94.035 -17.165 -93.095 ;
        RECT -16.800 -93.145 -16.570 -92.475 ;
        RECT -15.815 -93.085 -15.585 -92.475 ;
        RECT -16.770 -94.035 -16.600 -93.145 ;
        RECT -15.790 -94.035 -15.620 -93.085 ;
        RECT -26.735 -96.805 -26.120 -96.125 ;
        RECT -13.870 -96.300 -13.300 -91.940 ;
        RECT -6.695 -92.130 -3.730 -91.940 ;
        RECT -8.345 -92.475 -3.085 -92.130 ;
        RECT -8.345 -93.120 -8.145 -92.475 ;
        RECT -7.400 -93.120 -7.170 -92.475 ;
        RECT -6.410 -93.100 -6.180 -92.475 ;
        RECT -8.345 -94.035 -8.175 -93.120 ;
        RECT -7.365 -94.035 -7.195 -93.120 ;
        RECT -6.385 -94.035 -6.215 -93.100 ;
        RECT -5.845 -93.120 -5.615 -92.475 ;
        RECT -4.865 -93.095 -4.635 -92.475 ;
        RECT -5.815 -94.035 -5.645 -93.120 ;
        RECT -4.835 -94.035 -4.665 -93.095 ;
        RECT -4.300 -93.145 -4.070 -92.475 ;
        RECT -3.315 -93.085 -3.085 -92.475 ;
        RECT -4.270 -94.035 -4.100 -93.145 ;
        RECT -3.290 -94.035 -3.120 -93.085 ;
        RECT -1.460 -96.300 -0.885 -91.940 ;
        RECT 5.975 -92.130 8.940 -91.940 ;
        RECT 18.040 -92.130 21.005 -91.940 ;
        RECT 4.155 -92.475 9.415 -92.130 ;
        RECT 4.155 -93.120 4.355 -92.475 ;
        RECT 5.100 -93.120 5.330 -92.475 ;
        RECT 6.090 -93.100 6.320 -92.475 ;
        RECT 4.155 -94.035 4.325 -93.120 ;
        RECT 5.135 -94.035 5.305 -93.120 ;
        RECT 6.115 -94.035 6.285 -93.100 ;
        RECT 6.655 -93.120 6.885 -92.475 ;
        RECT 7.635 -93.095 7.865 -92.475 ;
        RECT 6.685 -94.035 6.855 -93.120 ;
        RECT 7.665 -94.035 7.835 -93.095 ;
        RECT 8.200 -93.145 8.430 -92.475 ;
        RECT 9.185 -93.085 9.415 -92.475 ;
        RECT 16.655 -92.475 21.915 -92.130 ;
        RECT 8.230 -94.035 8.400 -93.145 ;
        RECT 9.210 -94.035 9.380 -93.085 ;
        RECT 16.655 -93.120 16.855 -92.475 ;
        RECT 17.600 -93.120 17.830 -92.475 ;
        RECT 18.590 -93.100 18.820 -92.475 ;
        RECT 16.655 -94.035 16.825 -93.120 ;
        RECT 17.635 -94.035 17.805 -93.120 ;
        RECT 18.615 -94.035 18.785 -93.100 ;
        RECT 19.155 -93.120 19.385 -92.475 ;
        RECT 20.135 -93.095 20.365 -92.475 ;
        RECT 19.185 -94.035 19.355 -93.120 ;
        RECT 20.165 -94.035 20.335 -93.095 ;
        RECT 20.700 -93.145 20.930 -92.475 ;
        RECT 21.685 -93.085 21.915 -92.475 ;
        RECT 31.655 -92.475 36.915 -91.940 ;
        RECT 20.730 -94.035 20.900 -93.145 ;
        RECT 21.710 -94.035 21.880 -93.085 ;
        RECT 31.655 -93.120 31.855 -92.475 ;
        RECT 32.600 -93.120 32.830 -92.475 ;
        RECT 33.590 -93.100 33.820 -92.475 ;
        RECT 31.655 -94.035 31.825 -93.120 ;
        RECT 32.635 -94.035 32.805 -93.120 ;
        RECT 33.615 -94.035 33.785 -93.100 ;
        RECT 34.155 -93.120 34.385 -92.475 ;
        RECT 35.135 -93.095 35.365 -92.475 ;
        RECT 34.185 -94.035 34.355 -93.120 ;
        RECT 35.165 -94.035 35.335 -93.095 ;
        RECT 35.700 -93.145 35.930 -92.475 ;
        RECT 36.685 -93.085 36.915 -92.475 ;
        RECT 126.125 -92.750 131.640 -85.805 ;
        RECT 35.730 -94.035 35.900 -93.145 ;
        RECT 36.710 -94.035 36.880 -93.085 ;
        RECT -13.900 -96.980 -13.285 -96.300 ;
        RECT -1.485 -96.980 -0.870 -96.300 ;
        RECT -75.205 -100.010 -75.035 -98.555 ;
        RECT -74.225 -100.010 -74.055 -98.555 ;
        RECT -73.245 -100.010 -73.075 -98.555 ;
        RECT -66.490 -100.010 -66.320 -98.555 ;
        RECT -65.510 -100.010 -65.340 -98.555 ;
        RECT -64.530 -100.010 -64.360 -98.555 ;
        RECT -61.705 -100.010 -61.535 -98.555 ;
        RECT -60.725 -100.010 -60.555 -98.555 ;
        RECT -59.745 -100.010 -59.575 -98.555 ;
        RECT -52.990 -100.010 -52.820 -98.555 ;
        RECT -52.010 -100.010 -51.840 -98.555 ;
        RECT -51.030 -100.010 -50.860 -98.555 ;
        RECT -48.580 -100.010 -48.410 -98.555 ;
        RECT -47.600 -100.010 -47.430 -98.555 ;
        RECT -46.620 -100.010 -46.450 -98.555 ;
        RECT -1.490 -99.070 -0.875 -99.065 ;
        RECT -75.505 -100.025 -73.030 -100.010 ;
        RECT -66.795 -100.015 -59.530 -100.010 ;
        RECT -76.940 -100.035 -71.420 -100.025 ;
        RECT -66.795 -100.035 -57.965 -100.015 ;
        RECT -53.295 -100.035 -46.405 -100.010 ;
        RECT -95.515 -103.405 -95.345 -101.320 ;
        RECT -94.535 -103.405 -94.365 -101.320 ;
        RECT -93.555 -103.155 -93.385 -101.320 ;
        RECT -92.470 -103.155 -92.300 -102.325 ;
        RECT -91.490 -103.155 -91.320 -102.325 ;
        RECT -90.510 -103.155 -90.340 -102.325 ;
        RECT -89.530 -103.155 -89.360 -102.325 ;
        RECT -93.555 -103.405 -89.120 -103.155 ;
        RECT -88.280 -103.215 -88.110 -100.265 ;
        RECT -95.565 -103.650 -89.120 -103.405 ;
        RECT -95.565 -103.725 -93.355 -103.650 ;
        RECT -88.305 -103.845 -88.080 -103.215 ;
        RECT -87.300 -103.230 -87.130 -100.265 ;
        RECT -85.185 -103.225 -85.015 -100.265 ;
        RECT -76.940 -100.350 -46.405 -100.035 ;
        RECT -76.940 -100.365 -71.420 -100.350 ;
        RECT -60.330 -100.355 -57.965 -100.350 ;
        RECT -87.330 -103.845 -87.105 -103.230 ;
        RECT -85.220 -103.845 -84.995 -103.225 ;
        RECT -93.370 -103.930 -92.425 -103.895 ;
        RECT -93.555 -103.965 -92.425 -103.930 ;
        RECT -88.335 -103.965 -84.490 -103.845 ;
        RECT -95.565 -104.165 -84.490 -103.965 ;
        RECT -121.755 -104.175 -84.490 -104.165 ;
        RECT -121.755 -104.730 -85.010 -104.175 ;
        RECT -121.755 -105.160 -97.690 -104.730 ;
        RECT -121.755 -105.325 -97.740 -105.160 ;
        RECT -113.455 -105.510 -107.010 -105.325 ;
        RECT -113.405 -107.595 -113.235 -105.510 ;
        RECT -112.425 -107.595 -112.255 -105.510 ;
        RECT -111.445 -105.760 -107.010 -105.510 ;
        RECT -111.445 -107.595 -111.275 -105.760 ;
        RECT -110.360 -106.590 -110.190 -105.760 ;
        RECT -109.380 -106.590 -109.210 -105.760 ;
        RECT -108.400 -106.590 -108.230 -105.760 ;
        RECT -107.420 -106.590 -107.250 -105.760 ;
        RECT -104.540 -106.620 -104.370 -105.325 ;
        RECT -103.560 -106.620 -103.390 -105.325 ;
        RECT -102.580 -106.620 -102.410 -105.325 ;
        RECT -101.600 -106.620 -101.430 -105.325 ;
        RECT -98.890 -106.620 -98.720 -105.325 ;
        RECT -97.910 -106.620 -97.740 -105.325 ;
        RECT -94.715 -105.680 -93.855 -104.730 ;
        RECT -90.575 -104.815 -87.485 -104.730 ;
        RECT -90.575 -104.960 -88.360 -104.815 ;
        RECT -90.570 -105.030 -88.360 -104.960 ;
        RECT -90.570 -105.275 -84.125 -105.030 ;
        RECT -95.625 -106.175 -92.035 -105.680 ;
        RECT -95.385 -107.505 -95.215 -106.175 ;
        RECT -94.405 -107.505 -94.235 -106.175 ;
        RECT -93.425 -107.505 -93.255 -106.175 ;
        RECT -92.445 -107.505 -92.275 -106.175 ;
        RECT -90.520 -107.360 -90.350 -105.275 ;
        RECT -89.540 -107.360 -89.370 -105.275 ;
        RECT -88.560 -105.525 -84.125 -105.275 ;
        RECT -88.560 -107.360 -88.390 -105.525 ;
        RECT -87.475 -106.355 -87.305 -105.525 ;
        RECT -86.495 -106.355 -86.325 -105.525 ;
        RECT -85.515 -106.355 -85.345 -105.525 ;
        RECT -84.535 -106.355 -84.365 -105.525 ;
        RECT -74.630 -108.845 -73.865 -100.365 ;
        RECT -35.040 -101.095 -34.870 -99.640 ;
        RECT -34.060 -101.095 -33.890 -99.640 ;
        RECT -33.080 -101.095 -32.910 -99.640 ;
        RECT -13.905 -99.920 -13.290 -99.240 ;
        RECT -1.490 -99.380 0.040 -99.070 ;
        RECT -26.740 -100.640 -26.125 -99.960 ;
        RECT -35.085 -101.435 -32.610 -101.095 ;
        RECT -35.005 -103.385 -34.565 -101.435 ;
        RECT -34.090 -103.385 -33.650 -101.435 ;
        RECT -33.180 -103.385 -32.740 -101.435 ;
        RECT -37.570 -103.400 -32.050 -103.385 ;
        RECT -26.715 -103.400 -26.140 -100.640 ;
        RECT -20.960 -103.400 -18.595 -103.395 ;
        RECT -13.885 -103.400 -13.310 -99.920 ;
        RECT -7.610 -103.400 -6.995 -103.290 ;
        RECT -37.570 -103.715 -6.995 -103.400 ;
        RECT -37.570 -103.725 -32.050 -103.715 ;
        RECT -70.570 -108.285 -70.400 -106.200 ;
        RECT -69.590 -108.285 -69.420 -106.200 ;
        RECT -68.610 -108.035 -68.440 -106.200 ;
        RECT -67.525 -108.035 -67.355 -107.205 ;
        RECT -66.545 -108.035 -66.375 -107.205 ;
        RECT -65.565 -108.035 -65.395 -107.205 ;
        RECT -64.585 -108.035 -64.415 -107.205 ;
        RECT -68.610 -108.285 -64.175 -108.035 ;
        RECT -63.335 -108.095 -63.165 -105.145 ;
        RECT -70.620 -108.530 -64.175 -108.285 ;
        RECT -70.620 -108.605 -68.410 -108.530 ;
        RECT -63.360 -108.725 -63.135 -108.095 ;
        RECT -62.355 -108.110 -62.185 -105.145 ;
        RECT -60.240 -108.105 -60.070 -105.145 ;
        RECT -62.385 -108.725 -62.160 -108.110 ;
        RECT -60.275 -108.725 -60.050 -108.105 ;
        RECT -68.425 -108.810 -67.480 -108.775 ;
        RECT -68.610 -108.845 -67.480 -108.810 ;
        RECT -63.390 -108.845 -59.545 -108.725 ;
        RECT -74.630 -109.055 -59.545 -108.845 ;
        RECT -74.630 -109.610 -60.065 -109.055 ;
        RECT -74.630 -115.845 -73.865 -109.610 ;
        RECT -69.770 -110.560 -68.910 -109.610 ;
        RECT -65.630 -109.695 -62.540 -109.610 ;
        RECT -65.630 -109.840 -63.415 -109.695 ;
        RECT -65.625 -109.910 -63.415 -109.840 ;
        RECT -65.625 -110.155 -59.180 -109.910 ;
        RECT -70.680 -111.055 -67.090 -110.560 ;
        RECT -70.440 -112.385 -70.270 -111.055 ;
        RECT -69.460 -112.385 -69.290 -111.055 ;
        RECT -68.480 -112.385 -68.310 -111.055 ;
        RECT -67.500 -112.385 -67.330 -111.055 ;
        RECT -65.575 -112.240 -65.405 -110.155 ;
        RECT -64.595 -112.240 -64.425 -110.155 ;
        RECT -63.615 -110.405 -59.180 -110.155 ;
        RECT -63.615 -112.240 -63.445 -110.405 ;
        RECT -62.530 -111.235 -62.360 -110.405 ;
        RECT -61.550 -111.235 -61.380 -110.405 ;
        RECT -60.570 -111.235 -60.400 -110.405 ;
        RECT -59.590 -111.235 -59.420 -110.405 ;
        RECT -37.570 -112.200 -37.125 -103.725 ;
        RECT -36.135 -103.740 -33.660 -103.725 ;
        RECT -27.425 -103.735 -18.595 -103.715 ;
        RECT -27.425 -103.740 -20.160 -103.735 ;
        RECT -13.925 -103.740 -6.995 -103.715 ;
        RECT -35.835 -105.195 -35.665 -103.740 ;
        RECT -34.855 -105.195 -34.685 -103.740 ;
        RECT -33.875 -105.195 -33.705 -103.740 ;
        RECT -27.120 -105.195 -26.950 -103.740 ;
        RECT -26.140 -105.195 -25.970 -103.740 ;
        RECT -25.160 -105.195 -24.990 -103.740 ;
        RECT -22.335 -105.195 -22.165 -103.740 ;
        RECT -21.355 -105.195 -21.185 -103.740 ;
        RECT -20.375 -105.195 -20.205 -103.740 ;
        RECT -13.620 -105.195 -13.450 -103.740 ;
        RECT -12.640 -105.195 -12.470 -103.740 ;
        RECT -11.660 -105.195 -11.490 -103.740 ;
        RECT -9.210 -105.195 -9.040 -103.740 ;
        RECT -8.230 -105.195 -8.060 -103.740 ;
        RECT -7.610 -103.970 -6.995 -103.740 ;
        RECT -6.140 -103.420 -5.525 -103.285 ;
        RECT -1.465 -103.420 -0.890 -99.380 ;
        RECT 8.750 -103.420 9.365 -103.350 ;
        RECT -6.140 -103.815 9.365 -103.420 ;
        RECT -6.140 -103.820 -4.365 -103.815 ;
        RECT -6.140 -103.965 -5.370 -103.820 ;
        RECT -7.250 -105.195 -7.080 -103.970 ;
        RECT -5.540 -105.280 -5.370 -103.965 ;
        RECT -4.560 -105.280 -4.390 -103.820 ;
        RECT -1.850 -105.280 -1.680 -103.815 ;
        RECT -0.870 -105.280 -0.700 -103.815 ;
        RECT 0.110 -105.280 0.280 -103.815 ;
        RECT 1.090 -105.280 1.260 -103.815 ;
        RECT 2.885 -104.015 7.320 -103.815 ;
        RECT 3.125 -104.845 3.295 -104.015 ;
        RECT 4.105 -104.845 4.275 -104.015 ;
        RECT 5.085 -104.845 5.255 -104.015 ;
        RECT 6.065 -104.845 6.235 -104.015 ;
        RECT 7.150 -105.850 7.320 -104.015 ;
        RECT 8.130 -105.850 8.300 -103.815 ;
        RECT 8.750 -104.030 9.365 -103.815 ;
        RECT 10.695 -103.530 11.310 -103.345 ;
        RECT 16.835 -103.455 17.450 -103.230 ;
        RECT 15.145 -103.530 17.450 -103.455 ;
        RECT 10.695 -103.775 17.450 -103.530 ;
        RECT 10.695 -104.025 15.345 -103.775 ;
        RECT 9.110 -105.850 9.280 -104.030 ;
        RECT 11.150 -104.855 11.320 -104.025 ;
        RECT 12.130 -104.855 12.300 -104.025 ;
        RECT 13.110 -104.855 13.280 -104.025 ;
        RECT 14.090 -104.855 14.260 -104.025 ;
        RECT 15.175 -105.860 15.345 -104.025 ;
        RECT 16.155 -105.860 16.325 -103.775 ;
        RECT 16.835 -103.910 17.450 -103.775 ;
        RECT 18.840 -103.385 19.455 -103.220 ;
        RECT 18.840 -103.410 23.320 -103.385 ;
        RECT 25.620 -103.410 26.235 -103.245 ;
        RECT 18.840 -103.750 26.235 -103.410 ;
        RECT 18.840 -103.775 20.445 -103.750 ;
        RECT 22.960 -103.755 26.235 -103.750 ;
        RECT 18.840 -103.900 19.455 -103.775 ;
        RECT 17.135 -105.860 17.305 -103.910 ;
        RECT 19.270 -105.235 19.440 -103.900 ;
        RECT 20.250 -105.235 20.420 -103.775 ;
        RECT 22.960 -105.235 23.130 -103.755 ;
        RECT 23.940 -105.235 24.110 -103.755 ;
        RECT 24.920 -105.235 25.090 -103.755 ;
        RECT 25.620 -103.925 26.235 -103.755 ;
        RECT 31.700 -103.385 32.315 -103.250 ;
        RECT 31.700 -103.730 36.965 -103.385 ;
        RECT 25.900 -105.235 26.070 -103.925 ;
        RECT 31.700 -103.930 32.315 -103.730 ;
        RECT 31.705 -104.375 31.905 -103.930 ;
        RECT 32.650 -104.375 32.880 -103.730 ;
        RECT 33.640 -104.355 33.870 -103.730 ;
        RECT 31.705 -105.290 31.875 -104.375 ;
        RECT 32.685 -105.290 32.855 -104.375 ;
        RECT 33.665 -105.290 33.835 -104.355 ;
        RECT 34.205 -104.375 34.435 -103.730 ;
        RECT 35.185 -104.350 35.415 -103.730 ;
        RECT 34.235 -105.290 34.405 -104.375 ;
        RECT 35.215 -105.290 35.385 -104.350 ;
        RECT 35.750 -104.400 35.980 -103.730 ;
        RECT 36.735 -104.340 36.965 -103.730 ;
        RECT 35.780 -105.290 35.950 -104.400 ;
        RECT 36.760 -105.290 36.930 -104.340 ;
        RECT 97.865 -105.060 123.990 -104.745 ;
        RECT 102.625 -105.085 111.635 -105.060 ;
        RECT 116.125 -105.085 123.990 -105.060 ;
        RECT 134.790 -105.065 134.960 -103.735 ;
        RECT 135.770 -105.065 135.940 -103.735 ;
        RECT 136.750 -105.065 136.920 -103.735 ;
        RECT 137.730 -105.065 137.900 -103.735 ;
        RECT 102.930 -106.540 103.100 -105.085 ;
        RECT 103.910 -106.540 104.080 -105.085 ;
        RECT 104.890 -106.540 105.060 -105.085 ;
        RECT 107.115 -106.540 107.285 -105.085 ;
        RECT 108.095 -106.540 108.265 -105.085 ;
        RECT 109.075 -106.540 109.245 -105.085 ;
        RECT 116.430 -106.540 116.600 -105.085 ;
        RECT 117.410 -106.540 117.580 -105.085 ;
        RECT 118.390 -106.540 118.560 -105.085 ;
        RECT 120.615 -106.540 120.785 -105.085 ;
        RECT 121.595 -106.540 121.765 -105.085 ;
        RECT 122.575 -106.540 122.745 -105.085 ;
        RECT 123.545 -105.385 123.990 -105.085 ;
        RECT 134.550 -105.385 138.140 -105.065 ;
        RECT 123.545 -105.560 138.140 -105.385 ;
        RECT 123.545 -106.510 136.320 -105.560 ;
        RECT 139.655 -105.965 139.825 -103.880 ;
        RECT 140.635 -105.965 140.805 -103.880 ;
        RECT 141.615 -105.715 141.785 -103.880 ;
        RECT 142.700 -105.715 142.870 -104.885 ;
        RECT 143.680 -105.715 143.850 -104.885 ;
        RECT 144.660 -105.715 144.830 -104.885 ;
        RECT 145.640 -105.715 145.810 -104.885 ;
        RECT 176.990 -105.120 177.160 -103.790 ;
        RECT 177.970 -105.120 178.140 -103.790 ;
        RECT 178.950 -105.120 179.120 -103.790 ;
        RECT 179.930 -105.120 180.100 -103.790 ;
        RECT 176.750 -105.615 180.340 -105.120 ;
        RECT 141.615 -105.965 146.050 -105.715 ;
        RECT 139.605 -106.210 146.050 -105.965 ;
        RECT 139.605 -106.280 141.815 -106.210 ;
        RECT 151.840 -106.240 164.000 -105.890 ;
        RECT 139.600 -106.425 141.815 -106.280 ;
        RECT 139.600 -106.510 142.690 -106.425 ;
        RECT 150.005 -106.500 164.000 -106.240 ;
        RECT 150.005 -106.505 158.770 -106.500 ;
        RECT 123.545 -106.855 145.165 -106.510 ;
        RECT -36.325 -112.200 -36.155 -110.745 ;
        RECT -35.345 -112.200 -35.175 -110.745 ;
        RECT -34.365 -112.200 -34.195 -110.745 ;
        RECT -32.140 -112.200 -31.970 -110.745 ;
        RECT -31.160 -112.200 -30.990 -110.745 ;
        RECT -30.180 -112.200 -30.010 -110.745 ;
        RECT -22.825 -112.200 -22.655 -110.745 ;
        RECT -21.845 -112.200 -21.675 -110.745 ;
        RECT -20.865 -112.200 -20.695 -110.745 ;
        RECT -18.640 -112.200 -18.470 -110.745 ;
        RECT -17.660 -112.200 -17.490 -110.745 ;
        RECT -16.680 -112.200 -16.510 -110.745 ;
        RECT -37.570 -112.225 -29.705 -112.200 ;
        RECT -25.215 -112.225 -16.205 -112.200 ;
        RECT -37.570 -112.540 -11.445 -112.225 ;
        RECT 86.895 -112.490 87.065 -109.490 ;
        RECT 87.875 -112.410 88.045 -109.490 ;
        RECT -37.570 -115.735 -37.125 -112.540 ;
        RECT -56.550 -115.845 -37.125 -115.735 ;
        RECT -76.940 -116.160 -37.125 -115.845 ;
        RECT -76.940 -116.185 -69.075 -116.160 ;
        RECT -64.585 -116.185 -55.575 -116.160 ;
        RECT -76.940 -119.310 -76.495 -116.185 ;
        RECT -75.695 -117.640 -75.525 -116.185 ;
        RECT -74.715 -117.640 -74.545 -116.185 ;
        RECT -73.735 -117.640 -73.565 -116.185 ;
        RECT -71.510 -117.640 -71.340 -116.185 ;
        RECT -70.530 -117.640 -70.360 -116.185 ;
        RECT -69.550 -117.640 -69.380 -116.185 ;
        RECT -62.195 -117.640 -62.025 -116.185 ;
        RECT -61.215 -117.640 -61.045 -116.185 ;
        RECT -60.235 -117.640 -60.065 -116.185 ;
        RECT -58.010 -117.640 -57.840 -116.185 ;
        RECT -57.030 -117.640 -56.860 -116.185 ;
        RECT -56.050 -117.640 -55.880 -116.185 ;
        RECT -43.770 -116.765 -43.545 -116.160 ;
        RECT -41.660 -116.760 -41.435 -116.160 ;
        RECT -114.675 -120.145 -76.490 -119.310 ;
        RECT -43.750 -119.725 -43.580 -116.765 ;
        RECT -41.635 -119.725 -41.465 -116.760 ;
        RECT -40.685 -116.775 -40.460 -116.160 ;
        RECT -37.570 -116.735 -37.125 -116.160 ;
        RECT -40.655 -119.725 -40.485 -116.775 ;
        RECT -37.570 -117.180 -37.120 -116.735 ;
        RECT -36.130 -117.180 -34.785 -112.540 ;
        RECT -33.400 -117.180 -32.055 -112.540 ;
        RECT -29.015 -117.180 -27.670 -112.540 ;
        RECT -24.705 -117.180 -23.360 -112.540 ;
        RECT -20.190 -117.180 -18.845 -112.540 ;
        RECT -15.035 -117.180 -13.690 -112.540 ;
        RECT 86.850 -113.050 87.115 -112.490 ;
        RECT 87.830 -113.050 88.095 -112.410 ;
        RECT 86.850 -113.715 91.190 -113.050 ;
        RECT 93.500 -113.545 93.670 -112.090 ;
        RECT 94.480 -113.545 94.650 -112.090 ;
        RECT 95.460 -113.545 95.630 -112.090 ;
        RECT 97.910 -113.545 98.080 -112.090 ;
        RECT 98.890 -113.545 99.060 -112.090 ;
        RECT 99.870 -113.545 100.040 -112.090 ;
        RECT 106.625 -113.545 106.795 -112.090 ;
        RECT 107.605 -113.545 107.775 -112.090 ;
        RECT 108.585 -113.545 108.755 -112.090 ;
        RECT 111.410 -113.545 111.580 -112.090 ;
        RECT 112.390 -113.545 112.560 -112.090 ;
        RECT 113.370 -113.545 113.540 -112.090 ;
        RECT 120.125 -113.545 120.295 -112.090 ;
        RECT 121.105 -113.545 121.275 -112.090 ;
        RECT 122.085 -113.545 122.255 -112.090 ;
        RECT 93.455 -113.570 100.345 -113.545 ;
        RECT 106.580 -113.550 113.845 -113.545 ;
        RECT 105.015 -113.570 113.845 -113.550 ;
        RECT 120.080 -113.560 122.555 -113.545 ;
        RECT 123.545 -113.560 123.990 -106.855 ;
        RECT 134.610 -107.065 145.165 -106.855 ;
        RECT 150.005 -106.825 152.030 -106.505 ;
        RECT 147.190 -106.875 147.680 -106.860 ;
        RECT 150.005 -106.875 150.590 -106.825 ;
        RECT 134.610 -107.100 145.685 -107.065 ;
        RECT 146.050 -107.100 146.360 -106.960 ;
        RECT 134.610 -107.275 146.360 -107.100 ;
        RECT 136.620 -107.310 137.750 -107.275 ;
        RECT 136.805 -107.345 137.750 -107.310 ;
        RECT 141.840 -107.360 146.360 -107.275 ;
        RECT 141.840 -107.395 145.685 -107.360 ;
        RECT 134.610 -107.590 136.820 -107.515 ;
        RECT 134.610 -107.835 141.055 -107.590 ;
        RECT 134.660 -109.920 134.830 -107.835 ;
        RECT 135.640 -109.920 135.810 -107.835 ;
        RECT 136.620 -108.085 141.055 -107.835 ;
        RECT 141.870 -108.025 142.095 -107.395 ;
        RECT 142.845 -108.010 143.070 -107.395 ;
        RECT 136.620 -109.920 136.790 -108.085 ;
        RECT 137.705 -108.915 137.875 -108.085 ;
        RECT 138.685 -108.915 138.855 -108.085 ;
        RECT 139.665 -108.915 139.835 -108.085 ;
        RECT 140.645 -108.915 140.815 -108.085 ;
        RECT 141.895 -110.975 142.065 -108.025 ;
        RECT 142.875 -110.975 143.045 -108.010 ;
        RECT 144.955 -108.015 145.180 -107.395 ;
        RECT 146.050 -107.430 146.360 -107.360 ;
        RECT 147.190 -107.460 150.590 -106.875 ;
        RECT 151.840 -107.300 152.030 -106.825 ;
        RECT 152.825 -107.290 153.015 -106.505 ;
        RECT 147.190 -107.490 147.680 -107.460 ;
        RECT 144.990 -110.975 145.160 -108.015 ;
        RECT 151.855 -109.765 152.025 -107.300 ;
        RECT 152.835 -109.765 153.005 -107.290 ;
        RECT 155.785 -107.405 156.035 -106.505 ;
        RECT 156.415 -107.390 156.665 -106.505 ;
        RECT 157.570 -107.315 157.785 -106.505 ;
        RECT 158.555 -107.305 158.770 -106.505 ;
        RECT 163.390 -106.565 164.000 -106.500 ;
        RECT 177.660 -106.565 178.520 -105.615 ;
        RECT 181.855 -106.020 182.025 -103.935 ;
        RECT 182.835 -106.020 183.005 -103.935 ;
        RECT 183.815 -105.770 183.985 -103.935 ;
        RECT 184.900 -105.770 185.070 -104.940 ;
        RECT 185.880 -105.770 186.050 -104.940 ;
        RECT 186.860 -105.770 187.030 -104.940 ;
        RECT 187.840 -105.770 188.010 -104.940 ;
        RECT 221.305 -105.315 221.475 -103.985 ;
        RECT 222.285 -105.315 222.455 -103.985 ;
        RECT 223.265 -105.315 223.435 -103.985 ;
        RECT 224.245 -105.315 224.415 -103.985 ;
        RECT 221.065 -105.735 224.655 -105.315 ;
        RECT 183.815 -106.020 188.250 -105.770 ;
        RECT 200.900 -105.810 224.655 -105.735 ;
        RECT 200.900 -105.945 222.835 -105.810 ;
        RECT 181.805 -106.265 188.250 -106.020 ;
        RECT 181.805 -106.335 184.015 -106.265 ;
        RECT 194.040 -106.295 222.835 -105.945 ;
        RECT 226.170 -106.215 226.340 -104.130 ;
        RECT 227.150 -106.215 227.320 -104.130 ;
        RECT 228.130 -105.965 228.300 -104.130 ;
        RECT 229.215 -105.965 229.385 -105.135 ;
        RECT 230.195 -105.965 230.365 -105.135 ;
        RECT 231.175 -105.965 231.345 -105.135 ;
        RECT 232.155 -105.965 232.325 -105.135 ;
        RECT 267.295 -105.145 267.465 -103.815 ;
        RECT 268.275 -105.145 268.445 -103.815 ;
        RECT 269.255 -105.145 269.425 -103.815 ;
        RECT 270.235 -105.145 270.405 -103.815 ;
        RECT 267.055 -105.485 270.645 -105.145 ;
        RECT 245.155 -105.640 270.645 -105.485 ;
        RECT 228.130 -106.215 232.565 -105.965 ;
        RECT 245.155 -106.140 268.825 -105.640 ;
        RECT 272.160 -106.045 272.330 -103.960 ;
        RECT 273.140 -106.045 273.310 -103.960 ;
        RECT 274.120 -105.795 274.290 -103.960 ;
        RECT 311.065 -104.815 311.235 -103.485 ;
        RECT 312.045 -104.815 312.215 -103.485 ;
        RECT 313.025 -104.815 313.195 -103.485 ;
        RECT 314.005 -104.815 314.175 -103.485 ;
        RECT 275.205 -105.795 275.375 -104.965 ;
        RECT 276.185 -105.795 276.355 -104.965 ;
        RECT 277.165 -105.795 277.335 -104.965 ;
        RECT 278.145 -105.795 278.315 -104.965 ;
        RECT 310.825 -105.000 314.415 -104.815 ;
        RECT 291.070 -105.310 314.415 -105.000 ;
        RECT 274.120 -106.045 278.555 -105.795 ;
        RECT 291.070 -105.970 312.595 -105.310 ;
        RECT 315.930 -105.715 316.100 -103.630 ;
        RECT 316.910 -105.715 317.080 -103.630 ;
        RECT 317.890 -105.465 318.060 -103.630 ;
        RECT 318.975 -105.465 319.145 -104.635 ;
        RECT 319.955 -105.465 320.125 -104.635 ;
        RECT 320.935 -105.465 321.105 -104.635 ;
        RECT 321.915 -105.465 322.085 -104.635 ;
        RECT 356.830 -104.730 357.000 -103.400 ;
        RECT 357.810 -104.730 357.980 -103.400 ;
        RECT 358.790 -104.730 358.960 -103.400 ;
        RECT 359.770 -104.730 359.940 -103.400 ;
        RECT 356.590 -105.105 360.180 -104.730 ;
        RECT 334.805 -105.225 360.180 -105.105 ;
        RECT 317.890 -105.715 322.325 -105.465 ;
        RECT 334.805 -105.640 358.360 -105.225 ;
        RECT 361.695 -105.630 361.865 -103.545 ;
        RECT 362.675 -105.630 362.845 -103.545 ;
        RECT 363.655 -105.380 363.825 -103.545 ;
        RECT 403.650 -104.540 403.820 -103.210 ;
        RECT 404.630 -104.540 404.800 -103.210 ;
        RECT 405.610 -104.540 405.780 -103.210 ;
        RECT 406.590 -104.540 406.760 -103.210 ;
        RECT 364.740 -105.380 364.910 -104.550 ;
        RECT 365.720 -105.380 365.890 -104.550 ;
        RECT 366.700 -105.380 366.870 -104.550 ;
        RECT 367.680 -105.380 367.850 -104.550 ;
        RECT 403.410 -104.760 407.000 -104.540 ;
        RECT 380.615 -105.035 407.000 -104.760 ;
        RECT 363.655 -105.630 368.090 -105.380 ;
        RECT 380.615 -105.555 405.180 -105.035 ;
        RECT 408.515 -105.440 408.685 -103.355 ;
        RECT 409.495 -105.440 409.665 -103.355 ;
        RECT 410.475 -105.190 410.645 -103.355 ;
        RECT 411.560 -105.190 411.730 -104.360 ;
        RECT 412.540 -105.190 412.710 -104.360 ;
        RECT 413.520 -105.190 413.690 -104.360 ;
        RECT 414.500 -105.190 414.670 -104.360 ;
        RECT 410.475 -105.440 414.910 -105.190 ;
        RECT 429.490 -105.365 431.865 -85.805 ;
        RECT 181.800 -106.480 184.015 -106.335 ;
        RECT 181.800 -106.565 184.890 -106.480 ;
        RECT 192.205 -106.560 222.835 -106.295 ;
        RECT 226.120 -106.460 232.565 -106.215 ;
        RECT 226.120 -106.530 228.330 -106.460 ;
        RECT 238.355 -106.490 268.825 -106.140 ;
        RECT 272.110 -106.290 278.555 -106.045 ;
        RECT 284.345 -106.260 312.595 -105.970 ;
        RECT 315.880 -105.960 322.325 -105.715 ;
        RECT 315.880 -106.030 318.090 -105.960 ;
        RECT 328.115 -105.990 358.360 -105.640 ;
        RECT 361.645 -105.875 368.090 -105.630 ;
        RECT 361.645 -105.945 363.855 -105.875 ;
        RECT 373.880 -105.905 405.180 -105.555 ;
        RECT 408.465 -105.685 414.910 -105.440 ;
        RECT 408.465 -105.755 410.675 -105.685 ;
        RECT 420.700 -105.715 432.860 -105.365 ;
        RECT 315.875 -106.175 318.090 -106.030 ;
        RECT 326.280 -106.175 358.360 -105.990 ;
        RECT 361.640 -106.090 363.855 -105.945 ;
        RECT 372.045 -105.985 405.180 -105.905 ;
        RECT 408.460 -105.900 410.675 -105.755 ;
        RECT 408.460 -105.985 411.550 -105.900 ;
        RECT 418.865 -105.975 432.860 -105.715 ;
        RECT 418.865 -105.980 427.630 -105.975 ;
        RECT 361.640 -106.175 364.730 -106.090 ;
        RECT 372.045 -106.170 414.025 -105.985 ;
        RECT 315.875 -106.260 318.965 -106.175 ;
        RECT 326.280 -106.255 367.205 -106.175 ;
        RECT 272.110 -106.360 274.320 -106.290 ;
        RECT 284.345 -106.320 321.440 -106.260 ;
        RECT 163.390 -107.120 187.365 -106.565 ;
        RECT 192.205 -106.880 194.230 -106.560 ;
        RECT 189.390 -106.930 189.880 -106.915 ;
        RECT 192.205 -106.930 192.790 -106.880 ;
        RECT 163.390 -107.155 187.885 -107.120 ;
        RECT 188.250 -107.155 188.560 -107.015 ;
        RECT 155.810 -109.765 155.980 -107.405 ;
        RECT 156.460 -109.765 156.630 -107.390 ;
        RECT 157.600 -108.765 157.770 -107.315 ;
        RECT 158.580 -108.765 158.750 -107.305 ;
        RECT 163.390 -107.330 188.560 -107.155 ;
        RECT 118.470 -113.570 123.990 -113.560 ;
        RECT 93.455 -113.885 123.990 -113.570 ;
        RECT 105.015 -113.890 107.380 -113.885 ;
        RECT 105.965 -114.985 107.125 -113.890 ;
        RECT 118.470 -113.900 123.990 -113.885 ;
        RECT 105.675 -115.305 107.885 -114.985 ;
        RECT -37.570 -117.495 -11.445 -117.180 ;
        RECT -37.570 -117.520 -29.705 -117.495 ;
        RECT -25.215 -117.520 -16.205 -117.495 ;
        RECT -112.825 -120.840 -108.915 -120.145 ;
        RECT -107.035 -120.775 -104.445 -120.145 ;
        RECT -113.125 -121.505 -108.785 -120.840 ;
        RECT -107.110 -121.120 -104.340 -120.775 ;
        RECT -102.590 -120.780 -99.825 -120.145 ;
        RECT -102.590 -120.985 -99.815 -120.780 ;
        RECT -113.125 -122.065 -112.860 -121.505 ;
        RECT -113.080 -125.065 -112.910 -122.065 ;
        RECT -112.145 -122.145 -111.880 -121.505 ;
        RECT -107.085 -121.755 -106.845 -121.120 ;
        RECT -112.100 -125.065 -111.930 -122.145 ;
        RECT -107.050 -123.710 -106.880 -121.755 ;
        RECT -106.100 -121.785 -105.860 -121.120 ;
        RECT -102.585 -121.125 -99.815 -120.985 ;
        RECT -102.560 -121.760 -102.320 -121.125 ;
        RECT -106.070 -123.710 -105.900 -121.785 ;
        RECT -102.525 -123.715 -102.355 -121.760 ;
        RECT -101.575 -121.790 -101.335 -121.125 ;
        RECT -101.545 -123.715 -101.375 -121.790 ;
        RECT -76.940 -124.660 -76.495 -120.145 ;
        RECT -75.205 -124.645 -75.035 -123.190 ;
        RECT -74.225 -124.645 -74.055 -123.190 ;
        RECT -73.245 -124.645 -73.075 -123.190 ;
        RECT -66.490 -124.645 -66.320 -123.190 ;
        RECT -65.510 -124.645 -65.340 -123.190 ;
        RECT -64.530 -124.645 -64.360 -123.190 ;
        RECT -61.705 -124.645 -61.535 -123.190 ;
        RECT -60.725 -124.645 -60.555 -123.190 ;
        RECT -59.745 -124.645 -59.575 -123.190 ;
        RECT -52.990 -124.645 -52.820 -123.190 ;
        RECT -52.010 -124.645 -51.840 -123.190 ;
        RECT -51.030 -124.645 -50.860 -123.190 ;
        RECT -48.580 -124.645 -48.410 -123.190 ;
        RECT -47.600 -124.645 -47.430 -123.190 ;
        RECT -46.620 -124.645 -46.450 -123.190 ;
        RECT -75.505 -124.660 -73.030 -124.645 ;
        RECT -66.795 -124.650 -59.530 -124.645 ;
        RECT -76.940 -124.670 -71.420 -124.660 ;
        RECT -66.795 -124.670 -57.965 -124.650 ;
        RECT -53.295 -124.670 -46.405 -124.645 ;
        RECT -76.940 -124.985 -46.405 -124.670 ;
        RECT -76.940 -125.000 -71.420 -124.985 ;
        RECT -60.330 -124.990 -57.965 -124.985 ;
        RECT -95.515 -128.405 -95.345 -126.320 ;
        RECT -94.535 -128.405 -94.365 -126.320 ;
        RECT -93.555 -128.155 -93.385 -126.320 ;
        RECT -92.470 -128.155 -92.300 -127.325 ;
        RECT -91.490 -128.155 -91.320 -127.325 ;
        RECT -90.510 -128.155 -90.340 -127.325 ;
        RECT -89.530 -128.155 -89.360 -127.325 ;
        RECT -93.555 -128.405 -89.120 -128.155 ;
        RECT -88.280 -128.215 -88.110 -125.265 ;
        RECT -95.565 -128.650 -89.120 -128.405 ;
        RECT -95.565 -128.725 -93.355 -128.650 ;
        RECT -88.305 -128.845 -88.080 -128.215 ;
        RECT -87.300 -128.230 -87.130 -125.265 ;
        RECT -85.185 -128.225 -85.015 -125.265 ;
        RECT -37.570 -125.995 -37.125 -117.520 ;
        RECT -36.325 -118.975 -36.155 -117.520 ;
        RECT -35.345 -118.975 -35.175 -117.520 ;
        RECT -34.365 -118.975 -34.195 -117.520 ;
        RECT -32.140 -118.975 -31.970 -117.520 ;
        RECT -31.160 -118.975 -30.990 -117.520 ;
        RECT -30.180 -118.975 -30.010 -117.520 ;
        RECT -22.825 -118.975 -22.655 -117.520 ;
        RECT -21.845 -118.975 -21.675 -117.520 ;
        RECT -20.865 -118.975 -20.695 -117.520 ;
        RECT -18.640 -118.975 -18.470 -117.520 ;
        RECT -17.660 -118.975 -17.490 -117.520 ;
        RECT -16.680 -118.975 -16.510 -117.520 ;
        RECT 105.725 -117.890 105.895 -115.305 ;
        RECT 106.705 -117.890 106.875 -115.305 ;
        RECT 107.685 -117.890 107.855 -115.305 ;
        RECT -35.835 -125.980 -35.665 -124.525 ;
        RECT -34.855 -125.980 -34.685 -124.525 ;
        RECT -33.875 -125.980 -33.705 -124.525 ;
        RECT -27.120 -125.980 -26.950 -124.525 ;
        RECT -26.140 -125.980 -25.970 -124.525 ;
        RECT -25.160 -125.980 -24.990 -124.525 ;
        RECT -22.335 -125.980 -22.165 -124.525 ;
        RECT -21.355 -125.980 -21.185 -124.525 ;
        RECT -20.375 -125.980 -20.205 -124.525 ;
        RECT -13.620 -125.980 -13.450 -124.525 ;
        RECT -12.640 -125.980 -12.470 -124.525 ;
        RECT -11.660 -125.980 -11.490 -124.525 ;
        RECT -9.210 -125.980 -9.040 -124.525 ;
        RECT -8.230 -125.980 -8.060 -124.525 ;
        RECT -7.250 -125.750 -7.080 -124.525 ;
        RECT -7.610 -125.980 -6.995 -125.750 ;
        RECT -5.540 -125.755 -5.370 -124.440 ;
        RECT -36.135 -125.995 -33.660 -125.980 ;
        RECT -27.425 -125.985 -20.160 -125.980 ;
        RECT -37.570 -126.005 -32.050 -125.995 ;
        RECT -27.425 -126.005 -18.595 -125.985 ;
        RECT -13.925 -126.005 -6.995 -125.980 ;
        RECT -37.570 -126.320 -6.995 -126.005 ;
        RECT -37.570 -126.335 -32.050 -126.320 ;
        RECT -87.330 -128.845 -87.105 -128.230 ;
        RECT -85.220 -128.845 -84.995 -128.225 ;
        RECT -93.370 -128.930 -92.425 -128.895 ;
        RECT -93.555 -128.965 -92.425 -128.930 ;
        RECT -88.335 -128.965 -84.490 -128.845 ;
        RECT -101.735 -129.175 -84.490 -128.965 ;
        RECT -26.715 -129.080 -26.140 -126.320 ;
        RECT -20.960 -126.325 -18.595 -126.320 ;
        RECT -101.735 -129.730 -85.010 -129.175 ;
        RECT -101.735 -129.825 -93.855 -129.730 ;
        RECT -101.735 -134.800 -100.875 -129.825 ;
        RECT -94.715 -130.680 -93.855 -129.825 ;
        RECT -90.575 -129.815 -87.485 -129.730 ;
        RECT -26.740 -129.760 -26.125 -129.080 ;
        RECT -13.885 -129.800 -13.310 -126.320 ;
        RECT -7.610 -126.430 -6.995 -126.320 ;
        RECT -6.140 -125.900 -5.370 -125.755 ;
        RECT -4.560 -125.900 -4.390 -124.440 ;
        RECT -6.140 -125.905 -4.365 -125.900 ;
        RECT -1.850 -125.905 -1.680 -124.440 ;
        RECT -0.870 -125.905 -0.700 -124.440 ;
        RECT 0.110 -125.905 0.280 -124.440 ;
        RECT 1.090 -125.905 1.260 -124.440 ;
        RECT 3.125 -125.705 3.295 -124.875 ;
        RECT 4.105 -125.705 4.275 -124.875 ;
        RECT 5.085 -125.705 5.255 -124.875 ;
        RECT 6.065 -125.705 6.235 -124.875 ;
        RECT 7.150 -125.705 7.320 -123.870 ;
        RECT 2.885 -125.905 7.320 -125.705 ;
        RECT 8.130 -125.905 8.300 -123.870 ;
        RECT 9.110 -125.690 9.280 -123.870 ;
        RECT 8.750 -125.905 9.365 -125.690 ;
        RECT 11.150 -125.695 11.320 -124.865 ;
        RECT 12.130 -125.695 12.300 -124.865 ;
        RECT 13.110 -125.695 13.280 -124.865 ;
        RECT 14.090 -125.695 14.260 -124.865 ;
        RECT 15.175 -125.695 15.345 -123.860 ;
        RECT -6.140 -126.300 9.365 -125.905 ;
        RECT -6.140 -126.435 -5.525 -126.300 ;
        RECT -90.575 -129.960 -88.360 -129.815 ;
        RECT -90.570 -130.030 -88.360 -129.960 ;
        RECT -90.570 -130.275 -84.125 -130.030 ;
        RECT -95.625 -131.175 -92.035 -130.680 ;
        RECT -95.385 -132.505 -95.215 -131.175 ;
        RECT -94.405 -132.505 -94.235 -131.175 ;
        RECT -93.425 -132.505 -93.255 -131.175 ;
        RECT -92.445 -132.505 -92.275 -131.175 ;
        RECT -90.520 -132.360 -90.350 -130.275 ;
        RECT -89.540 -132.360 -89.370 -130.275 ;
        RECT -88.560 -130.525 -84.125 -130.275 ;
        RECT -13.905 -130.480 -13.290 -129.800 ;
        RECT -1.465 -130.340 -0.890 -126.300 ;
        RECT 8.750 -126.370 9.365 -126.300 ;
        RECT 10.695 -125.945 15.345 -125.695 ;
        RECT 16.155 -125.945 16.325 -123.860 ;
        RECT 17.135 -125.810 17.305 -123.860 ;
        RECT 86.870 -124.175 87.040 -122.220 ;
        RECT 87.850 -124.145 88.020 -122.220 ;
        RECT 16.835 -125.945 17.450 -125.810 ;
        RECT 19.270 -125.820 19.440 -124.485 ;
        RECT 10.695 -126.190 17.450 -125.945 ;
        RECT 10.695 -126.375 11.310 -126.190 ;
        RECT 15.145 -126.265 17.450 -126.190 ;
        RECT 16.835 -126.490 17.450 -126.265 ;
        RECT 18.840 -125.945 19.455 -125.820 ;
        RECT 20.250 -125.945 20.420 -124.485 ;
        RECT 18.840 -125.970 20.445 -125.945 ;
        RECT 22.960 -125.965 23.130 -124.485 ;
        RECT 23.940 -125.965 24.110 -124.485 ;
        RECT 24.920 -125.965 25.090 -124.485 ;
        RECT 25.900 -125.795 26.070 -124.485 ;
        RECT 31.705 -125.345 31.875 -124.430 ;
        RECT 32.685 -125.345 32.855 -124.430 ;
        RECT 31.705 -125.790 31.905 -125.345 ;
        RECT 25.620 -125.965 26.235 -125.795 ;
        RECT 22.960 -125.970 26.235 -125.965 ;
        RECT 18.840 -126.310 26.235 -125.970 ;
        RECT 18.840 -126.335 23.320 -126.310 ;
        RECT 18.840 -126.500 19.455 -126.335 ;
        RECT 25.620 -126.475 26.235 -126.310 ;
        RECT 31.700 -125.990 32.315 -125.790 ;
        RECT 32.650 -125.990 32.880 -125.345 ;
        RECT 33.665 -125.365 33.835 -124.430 ;
        RECT 34.235 -125.345 34.405 -124.430 ;
        RECT 33.640 -125.990 33.870 -125.365 ;
        RECT 34.205 -125.990 34.435 -125.345 ;
        RECT 35.215 -125.370 35.385 -124.430 ;
        RECT 35.780 -125.320 35.950 -124.430 ;
        RECT 35.185 -125.990 35.415 -125.370 ;
        RECT 35.750 -125.990 35.980 -125.320 ;
        RECT 36.760 -125.380 36.930 -124.430 ;
        RECT 86.835 -124.810 87.075 -124.175 ;
        RECT 87.820 -124.810 88.060 -124.145 ;
        RECT 91.600 -124.175 91.770 -122.220 ;
        RECT 92.580 -124.145 92.750 -122.220 ;
        RECT 91.565 -124.810 91.805 -124.175 ;
        RECT 92.550 -124.810 92.790 -124.145 ;
        RECT 94.955 -124.810 95.385 -124.770 ;
        RECT 82.720 -124.870 95.385 -124.810 ;
        RECT 96.180 -124.870 96.350 -123.390 ;
        RECT 97.160 -124.870 97.330 -123.390 ;
        RECT 98.140 -124.870 98.310 -123.390 ;
        RECT 99.120 -124.870 99.290 -123.390 ;
        RECT 100.555 -124.850 100.870 -124.780 ;
        RECT 101.830 -124.850 102.000 -123.390 ;
        RECT 102.810 -124.850 102.980 -123.390 ;
        RECT 103.960 -124.810 104.330 -124.780 ;
        RECT 105.475 -124.810 105.645 -123.355 ;
        RECT 106.455 -124.810 106.625 -123.355 ;
        RECT 107.435 -124.675 107.605 -123.355 ;
        RECT 109.875 -124.675 110.045 -120.500 ;
        RECT 110.855 -124.675 111.025 -120.500 ;
        RECT 111.875 -124.675 112.045 -120.500 ;
        RECT 112.855 -124.675 113.025 -120.500 ;
        RECT 114.875 -124.675 115.045 -120.500 ;
        RECT 115.855 -124.675 116.025 -120.500 ;
        RECT 116.875 -124.675 117.045 -120.500 ;
        RECT 117.855 -124.675 118.025 -120.500 ;
        RECT 119.875 -124.675 120.045 -120.500 ;
        RECT 120.855 -124.675 121.025 -120.500 ;
        RECT 121.875 -124.675 122.045 -120.500 ;
        RECT 122.855 -124.675 123.025 -120.500 ;
        RECT 123.545 -124.675 123.990 -113.900 ;
        RECT 147.225 -117.450 149.235 -117.120 ;
        RECT 134.750 -122.330 134.920 -121.000 ;
        RECT 135.730 -122.330 135.900 -121.000 ;
        RECT 136.710 -122.330 136.880 -121.000 ;
        RECT 137.690 -122.330 137.860 -121.000 ;
        RECT 134.510 -122.825 138.100 -122.330 ;
        RECT 135.420 -123.775 136.280 -122.825 ;
        RECT 139.615 -123.230 139.785 -121.145 ;
        RECT 140.595 -123.230 140.765 -121.145 ;
        RECT 141.575 -122.980 141.745 -121.145 ;
        RECT 142.660 -122.980 142.830 -122.150 ;
        RECT 143.640 -122.980 143.810 -122.150 ;
        RECT 144.620 -122.980 144.790 -122.150 ;
        RECT 145.600 -122.980 145.770 -122.150 ;
        RECT 141.575 -123.230 146.010 -122.980 ;
        RECT 139.565 -123.475 146.010 -123.230 ;
        RECT 139.565 -123.545 141.775 -123.475 ;
        RECT 139.560 -123.690 141.775 -123.545 ;
        RECT 139.560 -123.775 142.650 -123.690 ;
        RECT 134.570 -124.330 145.125 -123.775 ;
        RECT 147.225 -123.955 147.555 -117.450 ;
        RECT 134.570 -124.540 145.645 -124.330 ;
        RECT 147.140 -124.520 147.560 -123.955 ;
        RECT 148.905 -124.100 149.235 -117.450 ;
        RECT 163.390 -118.485 164.000 -107.330 ;
        RECT 178.820 -107.365 179.950 -107.330 ;
        RECT 179.005 -107.400 179.950 -107.365 ;
        RECT 184.040 -107.415 188.560 -107.330 ;
        RECT 184.040 -107.450 187.885 -107.415 ;
        RECT 176.810 -107.645 179.020 -107.570 ;
        RECT 176.810 -107.890 183.255 -107.645 ;
        RECT 176.860 -109.975 177.030 -107.890 ;
        RECT 177.840 -109.975 178.010 -107.890 ;
        RECT 178.820 -108.140 183.255 -107.890 ;
        RECT 184.070 -108.080 184.295 -107.450 ;
        RECT 185.045 -108.065 185.270 -107.450 ;
        RECT 178.820 -109.975 178.990 -108.140 ;
        RECT 179.905 -108.970 180.075 -108.140 ;
        RECT 180.885 -108.970 181.055 -108.140 ;
        RECT 181.865 -108.970 182.035 -108.140 ;
        RECT 182.845 -108.970 183.015 -108.140 ;
        RECT 184.095 -111.030 184.265 -108.080 ;
        RECT 185.075 -111.030 185.245 -108.065 ;
        RECT 187.155 -108.070 187.380 -107.450 ;
        RECT 188.250 -107.485 188.560 -107.415 ;
        RECT 189.390 -107.515 192.790 -106.930 ;
        RECT 194.040 -107.355 194.230 -106.880 ;
        RECT 195.025 -107.345 195.215 -106.560 ;
        RECT 189.390 -107.545 189.880 -107.515 ;
        RECT 187.190 -111.030 187.360 -108.070 ;
        RECT 194.055 -109.820 194.225 -107.355 ;
        RECT 195.035 -109.820 195.205 -107.345 ;
        RECT 197.985 -107.460 198.235 -106.560 ;
        RECT 198.615 -107.445 198.865 -106.560 ;
        RECT 199.770 -107.370 199.985 -106.560 ;
        RECT 200.755 -106.760 222.835 -106.560 ;
        RECT 226.115 -106.675 228.330 -106.530 ;
        RECT 236.520 -106.590 268.825 -106.490 ;
        RECT 272.105 -106.505 274.320 -106.360 ;
        RECT 272.105 -106.590 275.195 -106.505 ;
        RECT 282.510 -106.585 321.440 -106.320 ;
        RECT 226.115 -106.760 229.205 -106.675 ;
        RECT 236.520 -106.755 277.670 -106.590 ;
        RECT 200.755 -107.005 231.680 -106.760 ;
        RECT 200.755 -107.360 200.970 -107.005 ;
        RECT 198.010 -109.820 198.180 -107.460 ;
        RECT 198.660 -109.820 198.830 -107.445 ;
        RECT 199.800 -108.820 199.970 -107.370 ;
        RECT 200.780 -108.820 200.950 -107.360 ;
        RECT 189.425 -117.505 191.435 -117.175 ;
        RECT 163.390 -119.095 166.550 -118.485 ;
        RECT 153.090 -122.485 153.260 -121.155 ;
        RECT 154.070 -122.485 154.240 -121.155 ;
        RECT 155.050 -122.485 155.220 -121.155 ;
        RECT 156.030 -122.485 156.200 -121.155 ;
        RECT 152.850 -122.980 156.440 -122.485 ;
        RECT 153.760 -123.930 154.620 -122.980 ;
        RECT 157.955 -123.385 158.125 -121.300 ;
        RECT 158.935 -123.385 159.105 -121.300 ;
        RECT 159.915 -123.135 160.085 -121.300 ;
        RECT 161.000 -123.135 161.170 -122.305 ;
        RECT 161.980 -123.135 162.150 -122.305 ;
        RECT 162.960 -123.135 163.130 -122.305 ;
        RECT 163.940 -123.135 164.110 -122.305 ;
        RECT 159.915 -123.385 164.350 -123.135 ;
        RECT 157.905 -123.630 164.350 -123.385 ;
        RECT 157.905 -123.700 160.115 -123.630 ;
        RECT 157.900 -123.845 160.115 -123.700 ;
        RECT 157.900 -123.930 160.990 -123.845 ;
        RECT 152.910 -124.100 163.465 -123.930 ;
        RECT 165.940 -124.075 166.550 -119.095 ;
        RECT 176.950 -122.385 177.120 -121.055 ;
        RECT 177.930 -122.385 178.100 -121.055 ;
        RECT 178.910 -122.385 179.080 -121.055 ;
        RECT 179.890 -122.385 180.060 -121.055 ;
        RECT 176.710 -122.880 180.300 -122.385 ;
        RECT 177.620 -123.830 178.480 -122.880 ;
        RECT 181.815 -123.285 181.985 -121.200 ;
        RECT 182.795 -123.285 182.965 -121.200 ;
        RECT 183.775 -123.035 183.945 -121.200 ;
        RECT 184.860 -123.035 185.030 -122.205 ;
        RECT 185.840 -123.035 186.010 -122.205 ;
        RECT 186.820 -123.035 186.990 -122.205 ;
        RECT 187.800 -123.035 187.970 -122.205 ;
        RECT 183.775 -123.285 188.210 -123.035 ;
        RECT 181.765 -123.530 188.210 -123.285 ;
        RECT 181.765 -123.600 183.975 -123.530 ;
        RECT 181.760 -123.745 183.975 -123.600 ;
        RECT 181.760 -123.830 184.850 -123.745 ;
        RECT 148.905 -124.430 163.465 -124.100 ;
        RECT 164.240 -124.305 164.635 -124.150 ;
        RECT 152.910 -124.485 163.465 -124.430 ;
        RECT 163.740 -124.485 164.635 -124.305 ;
        RECT 136.580 -124.575 137.710 -124.540 ;
        RECT 136.765 -124.610 137.710 -124.575 ;
        RECT 141.800 -124.660 145.645 -124.540 ;
        RECT 107.435 -124.810 123.990 -124.675 ;
        RECT 103.960 -124.850 123.990 -124.810 ;
        RECT 100.555 -124.870 123.990 -124.850 ;
        RECT 82.720 -125.150 123.990 -124.870 ;
        RECT 134.570 -124.855 136.780 -124.780 ;
        RECT 134.570 -125.100 141.015 -124.855 ;
        RECT 82.720 -125.155 104.330 -125.150 ;
        RECT 36.735 -125.990 36.965 -125.380 ;
        RECT 31.700 -126.335 36.965 -125.990 ;
        RECT 31.700 -126.470 32.315 -126.335 ;
        RECT 82.720 -127.510 83.350 -125.155 ;
        RECT 94.955 -125.185 104.330 -125.155 ;
        RECT 94.955 -125.215 100.870 -125.185 ;
        RECT 103.960 -125.215 104.330 -125.185 ;
        RECT 107.545 -125.190 123.990 -125.150 ;
        RECT 94.955 -125.235 95.385 -125.215 ;
        RECT 100.555 -125.270 100.870 -125.215 ;
        RECT 134.620 -127.185 134.790 -125.100 ;
        RECT 135.600 -127.185 135.770 -125.100 ;
        RECT 136.580 -125.350 141.015 -125.100 ;
        RECT 141.830 -125.290 142.055 -124.660 ;
        RECT 142.805 -125.275 143.030 -124.660 ;
        RECT 136.580 -127.185 136.750 -125.350 ;
        RECT 137.665 -126.180 137.835 -125.350 ;
        RECT 138.645 -126.180 138.815 -125.350 ;
        RECT 139.625 -126.180 139.795 -125.350 ;
        RECT 140.605 -126.180 140.775 -125.350 ;
        RECT 64.375 -127.525 66.740 -127.520 ;
        RECT 77.830 -127.525 83.350 -127.510 ;
        RECT 52.815 -127.840 83.350 -127.525 ;
        RECT 52.815 -127.865 59.705 -127.840 ;
        RECT 64.375 -127.860 73.205 -127.840 ;
        RECT 77.830 -127.850 83.350 -127.840 ;
        RECT 65.940 -127.865 73.205 -127.860 ;
        RECT 79.440 -127.865 81.915 -127.850 ;
        RECT 52.860 -129.320 53.030 -127.865 ;
        RECT 53.840 -129.320 54.010 -127.865 ;
        RECT 54.820 -129.320 54.990 -127.865 ;
        RECT 57.270 -129.320 57.440 -127.865 ;
        RECT 58.250 -129.320 58.420 -127.865 ;
        RECT 59.230 -129.320 59.400 -127.865 ;
        RECT 65.985 -129.320 66.155 -127.865 ;
        RECT 66.965 -129.320 67.135 -127.865 ;
        RECT 67.945 -129.320 68.115 -127.865 ;
        RECT 70.770 -129.320 70.940 -127.865 ;
        RECT 71.750 -129.320 71.920 -127.865 ;
        RECT 72.730 -129.320 72.900 -127.865 ;
        RECT 79.485 -129.320 79.655 -127.865 ;
        RECT 80.465 -129.320 80.635 -127.865 ;
        RECT 81.445 -129.320 81.615 -127.865 ;
        RECT -88.560 -132.360 -88.390 -130.525 ;
        RECT -87.475 -131.355 -87.305 -130.525 ;
        RECT -86.495 -131.355 -86.325 -130.525 ;
        RECT -85.515 -131.355 -85.345 -130.525 ;
        RECT -84.535 -131.355 -84.365 -130.525 ;
        RECT -1.490 -130.650 0.040 -130.340 ;
        RECT -1.490 -130.655 -0.875 -130.650 ;
        RECT -26.735 -133.595 -26.120 -132.915 ;
        RECT -13.900 -133.420 -13.285 -132.740 ;
        RECT -1.485 -133.420 -0.870 -132.740 ;
        RECT -101.745 -135.235 -100.865 -134.800 ;
        RECT -114.765 -137.575 -114.595 -136.115 ;
        RECT -113.785 -137.495 -113.615 -136.115 ;
        RECT -111.075 -137.495 -110.905 -136.115 ;
        RECT -110.095 -137.495 -109.925 -136.115 ;
        RECT -109.115 -137.495 -108.945 -136.115 ;
        RECT -108.135 -137.495 -107.965 -136.115 ;
        RECT -33.345 -136.600 -33.175 -135.685 ;
        RECT -32.365 -136.600 -32.195 -135.685 ;
        RECT -33.345 -137.245 -33.145 -136.600 ;
        RECT -32.400 -137.245 -32.170 -136.600 ;
        RECT -31.385 -136.620 -31.215 -135.685 ;
        RECT -30.815 -136.600 -30.645 -135.685 ;
        RECT -31.410 -137.245 -31.180 -136.620 ;
        RECT -30.845 -137.245 -30.615 -136.600 ;
        RECT -29.835 -136.625 -29.665 -135.685 ;
        RECT -29.270 -136.575 -29.100 -135.685 ;
        RECT -29.865 -137.245 -29.635 -136.625 ;
        RECT -29.300 -137.245 -29.070 -136.575 ;
        RECT -28.290 -136.635 -28.120 -135.685 ;
        RECT -28.315 -137.245 -28.085 -136.635 ;
        RECT -113.875 -137.575 -100.865 -137.495 ;
        RECT -114.815 -137.910 -100.865 -137.575 ;
        RECT -33.345 -137.780 -28.085 -137.245 ;
        RECT -26.710 -137.780 -26.135 -133.595 ;
        RECT -20.845 -136.600 -20.675 -135.685 ;
        RECT -19.865 -136.600 -19.695 -135.685 ;
        RECT -20.845 -137.245 -20.645 -136.600 ;
        RECT -19.900 -137.245 -19.670 -136.600 ;
        RECT -18.885 -136.620 -18.715 -135.685 ;
        RECT -18.315 -136.600 -18.145 -135.685 ;
        RECT -18.910 -137.245 -18.680 -136.620 ;
        RECT -18.345 -137.245 -18.115 -136.600 ;
        RECT -17.335 -136.625 -17.165 -135.685 ;
        RECT -16.770 -136.575 -16.600 -135.685 ;
        RECT -17.365 -137.245 -17.135 -136.625 ;
        RECT -16.800 -137.245 -16.570 -136.575 ;
        RECT -15.790 -136.635 -15.620 -135.685 ;
        RECT -15.815 -137.245 -15.585 -136.635 ;
        RECT -20.845 -137.590 -15.585 -137.245 ;
        RECT -19.275 -137.780 -16.310 -137.590 ;
        RECT -13.870 -137.780 -13.300 -133.420 ;
        RECT -8.345 -136.600 -8.175 -135.685 ;
        RECT -7.365 -136.600 -7.195 -135.685 ;
        RECT -8.345 -137.245 -8.145 -136.600 ;
        RECT -7.400 -137.245 -7.170 -136.600 ;
        RECT -6.385 -136.620 -6.215 -135.685 ;
        RECT -5.815 -136.600 -5.645 -135.685 ;
        RECT -6.410 -137.245 -6.180 -136.620 ;
        RECT -5.845 -137.245 -5.615 -136.600 ;
        RECT -4.835 -136.625 -4.665 -135.685 ;
        RECT -4.270 -136.575 -4.100 -135.685 ;
        RECT -4.865 -137.245 -4.635 -136.625 ;
        RECT -4.300 -137.245 -4.070 -136.575 ;
        RECT -3.290 -136.635 -3.120 -135.685 ;
        RECT -3.315 -137.245 -3.085 -136.635 ;
        RECT -8.345 -137.590 -3.085 -137.245 ;
        RECT -6.695 -137.780 -3.730 -137.590 ;
        RECT -1.460 -137.780 -0.885 -133.420 ;
        RECT 4.155 -136.600 4.325 -135.685 ;
        RECT 5.135 -136.600 5.305 -135.685 ;
        RECT 4.155 -137.245 4.355 -136.600 ;
        RECT 5.100 -137.245 5.330 -136.600 ;
        RECT 6.115 -136.620 6.285 -135.685 ;
        RECT 6.685 -136.600 6.855 -135.685 ;
        RECT 6.090 -137.245 6.320 -136.620 ;
        RECT 6.655 -137.245 6.885 -136.600 ;
        RECT 7.665 -136.625 7.835 -135.685 ;
        RECT 8.230 -136.575 8.400 -135.685 ;
        RECT 7.635 -137.245 7.865 -136.625 ;
        RECT 8.200 -137.245 8.430 -136.575 ;
        RECT 9.210 -136.635 9.380 -135.685 ;
        RECT 16.655 -136.600 16.825 -135.685 ;
        RECT 17.635 -136.600 17.805 -135.685 ;
        RECT 9.185 -137.245 9.415 -136.635 ;
        RECT 4.155 -137.590 9.415 -137.245 ;
        RECT 16.655 -137.245 16.855 -136.600 ;
        RECT 17.600 -137.245 17.830 -136.600 ;
        RECT 18.615 -136.620 18.785 -135.685 ;
        RECT 19.185 -136.600 19.355 -135.685 ;
        RECT 18.590 -137.245 18.820 -136.620 ;
        RECT 19.155 -137.245 19.385 -136.600 ;
        RECT 20.165 -136.625 20.335 -135.685 ;
        RECT 20.730 -136.575 20.900 -135.685 ;
        RECT 20.135 -137.245 20.365 -136.625 ;
        RECT 20.700 -137.245 20.930 -136.575 ;
        RECT 21.710 -136.635 21.880 -135.685 ;
        RECT 31.655 -136.600 31.825 -135.685 ;
        RECT 32.635 -136.600 32.805 -135.685 ;
        RECT 21.685 -137.245 21.915 -136.635 ;
        RECT 16.655 -137.590 21.915 -137.245 ;
        RECT 31.655 -137.245 31.855 -136.600 ;
        RECT 32.600 -137.245 32.830 -136.600 ;
        RECT 33.615 -136.620 33.785 -135.685 ;
        RECT 34.185 -136.600 34.355 -135.685 ;
        RECT 33.590 -137.245 33.820 -136.620 ;
        RECT 34.155 -137.245 34.385 -136.600 ;
        RECT 35.165 -136.625 35.335 -135.685 ;
        RECT 35.730 -136.575 35.900 -135.685 ;
        RECT 35.135 -137.245 35.365 -136.625 ;
        RECT 35.700 -137.245 35.930 -136.575 ;
        RECT 36.710 -136.635 36.880 -135.685 ;
        RECT 62.290 -136.325 62.460 -134.870 ;
        RECT 63.270 -136.325 63.440 -134.870 ;
        RECT 64.250 -136.325 64.420 -134.870 ;
        RECT 66.475 -136.325 66.645 -134.870 ;
        RECT 67.455 -136.325 67.625 -134.870 ;
        RECT 68.435 -136.325 68.605 -134.870 ;
        RECT 75.790 -136.325 75.960 -134.870 ;
        RECT 76.770 -136.325 76.940 -134.870 ;
        RECT 77.750 -136.325 77.920 -134.870 ;
        RECT 79.975 -136.325 80.145 -134.870 ;
        RECT 80.955 -136.325 81.125 -134.870 ;
        RECT 81.935 -136.325 82.105 -134.870 ;
        RECT 82.905 -136.325 83.350 -127.850 ;
        RECT 141.855 -128.240 142.025 -125.290 ;
        RECT 142.835 -128.240 143.005 -125.275 ;
        RECT 144.915 -125.280 145.140 -124.660 ;
        RECT 152.910 -124.695 164.635 -124.485 ;
        RECT 154.920 -124.730 156.050 -124.695 ;
        RECT 155.105 -124.765 156.050 -124.730 ;
        RECT 160.140 -124.720 164.635 -124.695 ;
        RECT 160.140 -124.815 163.985 -124.720 ;
        RECT 152.910 -125.010 155.120 -124.935 ;
        RECT 152.910 -125.255 159.355 -125.010 ;
        RECT 144.950 -128.240 145.120 -125.280 ;
        RECT 152.960 -127.340 153.130 -125.255 ;
        RECT 153.940 -127.340 154.110 -125.255 ;
        RECT 154.920 -125.505 159.355 -125.255 ;
        RECT 160.170 -125.445 160.395 -124.815 ;
        RECT 161.145 -125.430 161.370 -124.815 ;
        RECT 154.920 -127.340 155.090 -125.505 ;
        RECT 156.005 -126.335 156.175 -125.505 ;
        RECT 156.985 -126.335 157.155 -125.505 ;
        RECT 157.965 -126.335 158.135 -125.505 ;
        RECT 158.945 -126.335 159.115 -125.505 ;
        RECT 160.195 -128.395 160.365 -125.445 ;
        RECT 161.175 -128.395 161.345 -125.430 ;
        RECT 163.255 -125.435 163.480 -124.815 ;
        RECT 164.240 -124.845 164.635 -124.720 ;
        RECT 165.490 -124.770 166.550 -124.075 ;
        RECT 176.770 -124.385 187.325 -123.830 ;
        RECT 189.425 -124.010 189.755 -117.505 ;
        RECT 176.770 -124.595 187.845 -124.385 ;
        RECT 189.340 -124.575 189.760 -124.010 ;
        RECT 191.105 -124.155 191.435 -117.505 ;
        RECT 205.590 -118.540 206.200 -107.005 ;
        RECT 221.125 -107.315 231.680 -107.005 ;
        RECT 236.520 -107.075 238.545 -106.755 ;
        RECT 233.705 -107.125 234.195 -107.110 ;
        RECT 236.520 -107.125 237.105 -107.075 ;
        RECT 221.125 -107.350 232.200 -107.315 ;
        RECT 232.565 -107.350 232.875 -107.210 ;
        RECT 221.125 -107.525 232.875 -107.350 ;
        RECT 223.135 -107.560 224.265 -107.525 ;
        RECT 223.320 -107.595 224.265 -107.560 ;
        RECT 228.355 -107.610 232.875 -107.525 ;
        RECT 228.355 -107.645 232.200 -107.610 ;
        RECT 221.125 -107.840 223.335 -107.765 ;
        RECT 221.125 -108.085 227.570 -107.840 ;
        RECT 221.175 -110.170 221.345 -108.085 ;
        RECT 222.155 -110.170 222.325 -108.085 ;
        RECT 223.135 -108.335 227.570 -108.085 ;
        RECT 228.385 -108.275 228.610 -107.645 ;
        RECT 229.360 -108.260 229.585 -107.645 ;
        RECT 223.135 -110.170 223.305 -108.335 ;
        RECT 224.220 -109.165 224.390 -108.335 ;
        RECT 225.200 -109.165 225.370 -108.335 ;
        RECT 226.180 -109.165 226.350 -108.335 ;
        RECT 227.160 -109.165 227.330 -108.335 ;
        RECT 228.410 -111.225 228.580 -108.275 ;
        RECT 229.390 -111.225 229.560 -108.260 ;
        RECT 231.470 -108.265 231.695 -107.645 ;
        RECT 232.565 -107.680 232.875 -107.610 ;
        RECT 233.705 -107.710 237.105 -107.125 ;
        RECT 238.355 -107.550 238.545 -107.075 ;
        RECT 239.340 -107.540 239.530 -106.755 ;
        RECT 233.705 -107.740 234.195 -107.710 ;
        RECT 231.505 -111.225 231.675 -108.265 ;
        RECT 238.370 -110.015 238.540 -107.550 ;
        RECT 239.350 -110.015 239.520 -107.540 ;
        RECT 242.300 -107.655 242.550 -106.755 ;
        RECT 242.930 -107.640 243.180 -106.755 ;
        RECT 244.085 -107.565 244.300 -106.755 ;
        RECT 245.070 -107.055 277.670 -106.755 ;
        RECT 282.510 -106.905 284.535 -106.585 ;
        RECT 279.695 -106.955 280.185 -106.940 ;
        RECT 282.510 -106.955 283.095 -106.905 ;
        RECT 245.070 -107.555 245.285 -107.055 ;
        RECT 242.325 -110.015 242.495 -107.655 ;
        RECT 242.975 -110.015 243.145 -107.640 ;
        RECT 244.115 -109.015 244.285 -107.565 ;
        RECT 245.095 -109.015 245.265 -107.555 ;
        RECT 233.740 -117.700 235.750 -117.370 ;
        RECT 205.590 -119.150 208.750 -118.540 ;
        RECT 195.290 -122.540 195.460 -121.210 ;
        RECT 196.270 -122.540 196.440 -121.210 ;
        RECT 197.250 -122.540 197.420 -121.210 ;
        RECT 198.230 -122.540 198.400 -121.210 ;
        RECT 195.050 -123.035 198.640 -122.540 ;
        RECT 195.960 -123.985 196.820 -123.035 ;
        RECT 200.155 -123.440 200.325 -121.355 ;
        RECT 201.135 -123.440 201.305 -121.355 ;
        RECT 202.115 -123.190 202.285 -121.355 ;
        RECT 203.200 -123.190 203.370 -122.360 ;
        RECT 204.180 -123.190 204.350 -122.360 ;
        RECT 205.160 -123.190 205.330 -122.360 ;
        RECT 206.140 -123.190 206.310 -122.360 ;
        RECT 202.115 -123.440 206.550 -123.190 ;
        RECT 200.105 -123.685 206.550 -123.440 ;
        RECT 200.105 -123.755 202.315 -123.685 ;
        RECT 200.100 -123.900 202.315 -123.755 ;
        RECT 200.100 -123.985 203.190 -123.900 ;
        RECT 195.110 -124.155 205.665 -123.985 ;
        RECT 208.140 -124.130 208.750 -119.150 ;
        RECT 221.265 -122.580 221.435 -121.250 ;
        RECT 222.245 -122.580 222.415 -121.250 ;
        RECT 223.225 -122.580 223.395 -121.250 ;
        RECT 224.205 -122.580 224.375 -121.250 ;
        RECT 221.025 -123.075 224.615 -122.580 ;
        RECT 221.935 -124.025 222.795 -123.075 ;
        RECT 226.130 -123.480 226.300 -121.395 ;
        RECT 227.110 -123.480 227.280 -121.395 ;
        RECT 228.090 -123.230 228.260 -121.395 ;
        RECT 229.175 -123.230 229.345 -122.400 ;
        RECT 230.155 -123.230 230.325 -122.400 ;
        RECT 231.135 -123.230 231.305 -122.400 ;
        RECT 232.115 -123.230 232.285 -122.400 ;
        RECT 228.090 -123.480 232.525 -123.230 ;
        RECT 226.080 -123.725 232.525 -123.480 ;
        RECT 226.080 -123.795 228.290 -123.725 ;
        RECT 226.075 -123.940 228.290 -123.795 ;
        RECT 226.075 -124.025 229.165 -123.940 ;
        RECT 191.105 -124.485 205.665 -124.155 ;
        RECT 206.440 -124.360 206.835 -124.205 ;
        RECT 195.110 -124.540 205.665 -124.485 ;
        RECT 205.940 -124.540 206.835 -124.360 ;
        RECT 178.780 -124.630 179.910 -124.595 ;
        RECT 178.965 -124.665 179.910 -124.630 ;
        RECT 184.000 -124.715 187.845 -124.595 ;
        RECT 165.490 -124.910 166.185 -124.770 ;
        RECT 176.770 -124.910 178.980 -124.835 ;
        RECT 176.770 -125.155 183.215 -124.910 ;
        RECT 163.290 -128.395 163.460 -125.435 ;
        RECT 176.820 -127.240 176.990 -125.155 ;
        RECT 177.800 -127.240 177.970 -125.155 ;
        RECT 178.780 -125.405 183.215 -125.155 ;
        RECT 184.030 -125.345 184.255 -124.715 ;
        RECT 185.005 -125.330 185.230 -124.715 ;
        RECT 178.780 -127.240 178.950 -125.405 ;
        RECT 179.865 -126.235 180.035 -125.405 ;
        RECT 180.845 -126.235 181.015 -125.405 ;
        RECT 181.825 -126.235 181.995 -125.405 ;
        RECT 182.805 -126.235 182.975 -125.405 ;
        RECT 184.055 -128.295 184.225 -125.345 ;
        RECT 185.035 -128.295 185.205 -125.330 ;
        RECT 187.115 -125.335 187.340 -124.715 ;
        RECT 195.110 -124.750 206.835 -124.540 ;
        RECT 197.120 -124.785 198.250 -124.750 ;
        RECT 197.305 -124.820 198.250 -124.785 ;
        RECT 202.340 -124.775 206.835 -124.750 ;
        RECT 202.340 -124.870 206.185 -124.775 ;
        RECT 195.110 -125.065 197.320 -124.990 ;
        RECT 195.110 -125.310 201.555 -125.065 ;
        RECT 187.150 -128.295 187.320 -125.335 ;
        RECT 195.160 -127.395 195.330 -125.310 ;
        RECT 196.140 -127.395 196.310 -125.310 ;
        RECT 197.120 -125.560 201.555 -125.310 ;
        RECT 202.370 -125.500 202.595 -124.870 ;
        RECT 203.345 -125.485 203.570 -124.870 ;
        RECT 197.120 -127.395 197.290 -125.560 ;
        RECT 198.205 -126.390 198.375 -125.560 ;
        RECT 199.185 -126.390 199.355 -125.560 ;
        RECT 200.165 -126.390 200.335 -125.560 ;
        RECT 201.145 -126.390 201.315 -125.560 ;
        RECT 202.395 -128.450 202.565 -125.500 ;
        RECT 203.375 -128.450 203.545 -125.485 ;
        RECT 205.455 -125.490 205.680 -124.870 ;
        RECT 206.440 -124.900 206.835 -124.775 ;
        RECT 207.690 -124.825 208.750 -124.130 ;
        RECT 221.085 -124.580 231.640 -124.025 ;
        RECT 233.740 -124.205 234.070 -117.700 ;
        RECT 221.085 -124.790 232.160 -124.580 ;
        RECT 233.655 -124.770 234.075 -124.205 ;
        RECT 235.420 -124.350 235.750 -117.700 ;
        RECT 249.905 -118.735 250.515 -107.055 ;
        RECT 267.115 -107.145 277.670 -107.055 ;
        RECT 267.115 -107.180 278.190 -107.145 ;
        RECT 278.555 -107.180 278.865 -107.040 ;
        RECT 267.115 -107.355 278.865 -107.180 ;
        RECT 269.125 -107.390 270.255 -107.355 ;
        RECT 269.310 -107.425 270.255 -107.390 ;
        RECT 274.345 -107.440 278.865 -107.355 ;
        RECT 274.345 -107.475 278.190 -107.440 ;
        RECT 267.115 -107.670 269.325 -107.595 ;
        RECT 267.115 -107.915 273.560 -107.670 ;
        RECT 267.165 -110.000 267.335 -107.915 ;
        RECT 268.145 -110.000 268.315 -107.915 ;
        RECT 269.125 -108.165 273.560 -107.915 ;
        RECT 274.375 -108.105 274.600 -107.475 ;
        RECT 275.350 -108.090 275.575 -107.475 ;
        RECT 269.125 -110.000 269.295 -108.165 ;
        RECT 270.210 -108.995 270.380 -108.165 ;
        RECT 271.190 -108.995 271.360 -108.165 ;
        RECT 272.170 -108.995 272.340 -108.165 ;
        RECT 273.150 -108.995 273.320 -108.165 ;
        RECT 274.400 -111.055 274.570 -108.105 ;
        RECT 275.380 -111.055 275.550 -108.090 ;
        RECT 277.460 -108.095 277.685 -107.475 ;
        RECT 278.555 -107.510 278.865 -107.440 ;
        RECT 279.695 -107.540 283.095 -106.955 ;
        RECT 284.345 -107.380 284.535 -106.905 ;
        RECT 285.330 -107.370 285.520 -106.585 ;
        RECT 279.695 -107.570 280.185 -107.540 ;
        RECT 277.495 -111.055 277.665 -108.095 ;
        RECT 284.360 -109.845 284.530 -107.380 ;
        RECT 285.340 -109.845 285.510 -107.370 ;
        RECT 288.290 -107.485 288.540 -106.585 ;
        RECT 288.920 -107.470 289.170 -106.585 ;
        RECT 290.075 -107.395 290.290 -106.585 ;
        RECT 291.060 -106.815 321.440 -106.585 ;
        RECT 326.280 -106.575 328.305 -106.255 ;
        RECT 323.465 -106.625 323.955 -106.610 ;
        RECT 326.280 -106.625 326.865 -106.575 ;
        RECT 291.060 -106.850 321.960 -106.815 ;
        RECT 322.325 -106.850 322.635 -106.710 ;
        RECT 291.060 -106.895 322.635 -106.850 ;
        RECT 291.060 -107.385 291.275 -106.895 ;
        RECT 288.315 -109.845 288.485 -107.485 ;
        RECT 288.965 -109.845 289.135 -107.470 ;
        RECT 290.105 -108.845 290.275 -107.395 ;
        RECT 291.085 -108.845 291.255 -107.385 ;
        RECT 279.730 -117.530 281.740 -117.200 ;
        RECT 249.905 -119.345 253.065 -118.735 ;
        RECT 239.605 -122.735 239.775 -121.405 ;
        RECT 240.585 -122.735 240.755 -121.405 ;
        RECT 241.565 -122.735 241.735 -121.405 ;
        RECT 242.545 -122.735 242.715 -121.405 ;
        RECT 239.365 -123.230 242.955 -122.735 ;
        RECT 240.275 -124.180 241.135 -123.230 ;
        RECT 244.470 -123.635 244.640 -121.550 ;
        RECT 245.450 -123.635 245.620 -121.550 ;
        RECT 246.430 -123.385 246.600 -121.550 ;
        RECT 247.515 -123.385 247.685 -122.555 ;
        RECT 248.495 -123.385 248.665 -122.555 ;
        RECT 249.475 -123.385 249.645 -122.555 ;
        RECT 250.455 -123.385 250.625 -122.555 ;
        RECT 246.430 -123.635 250.865 -123.385 ;
        RECT 244.420 -123.880 250.865 -123.635 ;
        RECT 244.420 -123.950 246.630 -123.880 ;
        RECT 244.415 -124.095 246.630 -123.950 ;
        RECT 244.415 -124.180 247.505 -124.095 ;
        RECT 239.425 -124.350 249.980 -124.180 ;
        RECT 252.455 -124.325 253.065 -119.345 ;
        RECT 267.255 -122.410 267.425 -121.080 ;
        RECT 268.235 -122.410 268.405 -121.080 ;
        RECT 269.215 -122.410 269.385 -121.080 ;
        RECT 270.195 -122.410 270.365 -121.080 ;
        RECT 267.015 -122.905 270.605 -122.410 ;
        RECT 267.925 -123.855 268.785 -122.905 ;
        RECT 272.120 -123.310 272.290 -121.225 ;
        RECT 273.100 -123.310 273.270 -121.225 ;
        RECT 274.080 -123.060 274.250 -121.225 ;
        RECT 275.165 -123.060 275.335 -122.230 ;
        RECT 276.145 -123.060 276.315 -122.230 ;
        RECT 277.125 -123.060 277.295 -122.230 ;
        RECT 278.105 -123.060 278.275 -122.230 ;
        RECT 274.080 -123.310 278.515 -123.060 ;
        RECT 272.070 -123.555 278.515 -123.310 ;
        RECT 272.070 -123.625 274.280 -123.555 ;
        RECT 272.065 -123.770 274.280 -123.625 ;
        RECT 272.065 -123.855 275.155 -123.770 ;
        RECT 235.420 -124.680 249.980 -124.350 ;
        RECT 250.755 -124.555 251.150 -124.400 ;
        RECT 239.425 -124.735 249.980 -124.680 ;
        RECT 250.255 -124.735 251.150 -124.555 ;
        RECT 223.095 -124.825 224.225 -124.790 ;
        RECT 207.690 -124.965 208.385 -124.825 ;
        RECT 223.280 -124.860 224.225 -124.825 ;
        RECT 228.315 -124.910 232.160 -124.790 ;
        RECT 221.085 -125.105 223.295 -125.030 ;
        RECT 221.085 -125.350 227.530 -125.105 ;
        RECT 205.490 -128.450 205.660 -125.490 ;
        RECT 221.135 -127.435 221.305 -125.350 ;
        RECT 222.115 -127.435 222.285 -125.350 ;
        RECT 223.095 -125.600 227.530 -125.350 ;
        RECT 228.345 -125.540 228.570 -124.910 ;
        RECT 229.320 -125.525 229.545 -124.910 ;
        RECT 223.095 -127.435 223.265 -125.600 ;
        RECT 224.180 -126.430 224.350 -125.600 ;
        RECT 225.160 -126.430 225.330 -125.600 ;
        RECT 226.140 -126.430 226.310 -125.600 ;
        RECT 227.120 -126.430 227.290 -125.600 ;
        RECT 228.370 -128.490 228.540 -125.540 ;
        RECT 229.350 -128.490 229.520 -125.525 ;
        RECT 231.430 -125.530 231.655 -124.910 ;
        RECT 239.425 -124.945 251.150 -124.735 ;
        RECT 241.435 -124.980 242.565 -124.945 ;
        RECT 241.620 -125.015 242.565 -124.980 ;
        RECT 246.655 -124.970 251.150 -124.945 ;
        RECT 246.655 -125.065 250.500 -124.970 ;
        RECT 239.425 -125.260 241.635 -125.185 ;
        RECT 239.425 -125.505 245.870 -125.260 ;
        RECT 231.465 -128.490 231.635 -125.530 ;
        RECT 239.475 -127.590 239.645 -125.505 ;
        RECT 240.455 -127.590 240.625 -125.505 ;
        RECT 241.435 -125.755 245.870 -125.505 ;
        RECT 246.685 -125.695 246.910 -125.065 ;
        RECT 247.660 -125.680 247.885 -125.065 ;
        RECT 241.435 -127.590 241.605 -125.755 ;
        RECT 242.520 -126.585 242.690 -125.755 ;
        RECT 243.500 -126.585 243.670 -125.755 ;
        RECT 244.480 -126.585 244.650 -125.755 ;
        RECT 245.460 -126.585 245.630 -125.755 ;
        RECT 246.710 -128.645 246.880 -125.695 ;
        RECT 247.690 -128.645 247.860 -125.680 ;
        RECT 249.770 -125.685 249.995 -125.065 ;
        RECT 250.755 -125.095 251.150 -124.970 ;
        RECT 252.005 -125.020 253.065 -124.325 ;
        RECT 267.075 -124.410 277.630 -123.855 ;
        RECT 279.730 -124.035 280.060 -117.530 ;
        RECT 267.075 -124.620 278.150 -124.410 ;
        RECT 279.645 -124.600 280.065 -124.035 ;
        RECT 281.410 -124.180 281.740 -117.530 ;
        RECT 295.895 -118.565 296.505 -106.895 ;
        RECT 310.885 -107.025 322.635 -106.895 ;
        RECT 312.895 -107.060 314.025 -107.025 ;
        RECT 313.080 -107.095 314.025 -107.060 ;
        RECT 318.115 -107.110 322.635 -107.025 ;
        RECT 318.115 -107.145 321.960 -107.110 ;
        RECT 310.885 -107.340 313.095 -107.265 ;
        RECT 310.885 -107.585 317.330 -107.340 ;
        RECT 310.935 -109.670 311.105 -107.585 ;
        RECT 311.915 -109.670 312.085 -107.585 ;
        RECT 312.895 -107.835 317.330 -107.585 ;
        RECT 318.145 -107.775 318.370 -107.145 ;
        RECT 319.120 -107.760 319.345 -107.145 ;
        RECT 312.895 -109.670 313.065 -107.835 ;
        RECT 313.980 -108.665 314.150 -107.835 ;
        RECT 314.960 -108.665 315.130 -107.835 ;
        RECT 315.940 -108.665 316.110 -107.835 ;
        RECT 316.920 -108.665 317.090 -107.835 ;
        RECT 318.170 -110.725 318.340 -107.775 ;
        RECT 319.150 -110.725 319.320 -107.760 ;
        RECT 321.230 -107.765 321.455 -107.145 ;
        RECT 322.325 -107.180 322.635 -107.110 ;
        RECT 323.465 -107.210 326.865 -106.625 ;
        RECT 328.115 -107.050 328.305 -106.575 ;
        RECT 329.100 -107.040 329.290 -106.255 ;
        RECT 323.465 -107.240 323.955 -107.210 ;
        RECT 321.265 -110.725 321.435 -107.765 ;
        RECT 328.130 -109.515 328.300 -107.050 ;
        RECT 329.110 -109.515 329.280 -107.040 ;
        RECT 332.060 -107.155 332.310 -106.255 ;
        RECT 332.690 -107.140 332.940 -106.255 ;
        RECT 333.845 -107.065 334.060 -106.255 ;
        RECT 334.805 -106.425 367.205 -106.255 ;
        RECT 334.830 -107.055 335.045 -106.425 ;
        RECT 332.085 -109.515 332.255 -107.155 ;
        RECT 332.735 -109.515 332.905 -107.140 ;
        RECT 333.875 -108.515 334.045 -107.065 ;
        RECT 334.855 -108.515 335.025 -107.055 ;
        RECT 323.500 -117.200 325.510 -116.870 ;
        RECT 295.895 -119.175 299.055 -118.565 ;
        RECT 285.595 -122.565 285.765 -121.235 ;
        RECT 286.575 -122.565 286.745 -121.235 ;
        RECT 287.555 -122.565 287.725 -121.235 ;
        RECT 288.535 -122.565 288.705 -121.235 ;
        RECT 285.355 -123.060 288.945 -122.565 ;
        RECT 286.265 -124.010 287.125 -123.060 ;
        RECT 290.460 -123.465 290.630 -121.380 ;
        RECT 291.440 -123.465 291.610 -121.380 ;
        RECT 292.420 -123.215 292.590 -121.380 ;
        RECT 293.505 -123.215 293.675 -122.385 ;
        RECT 294.485 -123.215 294.655 -122.385 ;
        RECT 295.465 -123.215 295.635 -122.385 ;
        RECT 296.445 -123.215 296.615 -122.385 ;
        RECT 292.420 -123.465 296.855 -123.215 ;
        RECT 290.410 -123.710 296.855 -123.465 ;
        RECT 290.410 -123.780 292.620 -123.710 ;
        RECT 290.405 -123.925 292.620 -123.780 ;
        RECT 290.405 -124.010 293.495 -123.925 ;
        RECT 285.415 -124.180 295.970 -124.010 ;
        RECT 298.445 -124.155 299.055 -119.175 ;
        RECT 311.025 -122.080 311.195 -120.750 ;
        RECT 312.005 -122.080 312.175 -120.750 ;
        RECT 312.985 -122.080 313.155 -120.750 ;
        RECT 313.965 -122.080 314.135 -120.750 ;
        RECT 310.785 -122.575 314.375 -122.080 ;
        RECT 311.695 -123.525 312.555 -122.575 ;
        RECT 315.890 -122.980 316.060 -120.895 ;
        RECT 316.870 -122.980 317.040 -120.895 ;
        RECT 317.850 -122.730 318.020 -120.895 ;
        RECT 318.935 -122.730 319.105 -121.900 ;
        RECT 319.915 -122.730 320.085 -121.900 ;
        RECT 320.895 -122.730 321.065 -121.900 ;
        RECT 321.875 -122.730 322.045 -121.900 ;
        RECT 317.850 -122.980 322.285 -122.730 ;
        RECT 315.840 -123.225 322.285 -122.980 ;
        RECT 315.840 -123.295 318.050 -123.225 ;
        RECT 315.835 -123.440 318.050 -123.295 ;
        RECT 315.835 -123.525 318.925 -123.440 ;
        RECT 281.410 -124.510 295.970 -124.180 ;
        RECT 296.745 -124.385 297.140 -124.230 ;
        RECT 285.415 -124.565 295.970 -124.510 ;
        RECT 296.245 -124.565 297.140 -124.385 ;
        RECT 269.085 -124.655 270.215 -124.620 ;
        RECT 269.270 -124.690 270.215 -124.655 ;
        RECT 274.305 -124.740 278.150 -124.620 ;
        RECT 267.075 -124.935 269.285 -124.860 ;
        RECT 252.005 -125.160 252.700 -125.020 ;
        RECT 267.075 -125.180 273.520 -124.935 ;
        RECT 249.805 -128.645 249.975 -125.685 ;
        RECT 267.125 -127.265 267.295 -125.180 ;
        RECT 268.105 -127.265 268.275 -125.180 ;
        RECT 269.085 -125.430 273.520 -125.180 ;
        RECT 274.335 -125.370 274.560 -124.740 ;
        RECT 275.310 -125.355 275.535 -124.740 ;
        RECT 269.085 -127.265 269.255 -125.430 ;
        RECT 270.170 -126.260 270.340 -125.430 ;
        RECT 271.150 -126.260 271.320 -125.430 ;
        RECT 272.130 -126.260 272.300 -125.430 ;
        RECT 273.110 -126.260 273.280 -125.430 ;
        RECT 274.360 -128.320 274.530 -125.370 ;
        RECT 275.340 -128.320 275.510 -125.355 ;
        RECT 277.420 -125.360 277.645 -124.740 ;
        RECT 285.415 -124.775 297.140 -124.565 ;
        RECT 287.425 -124.810 288.555 -124.775 ;
        RECT 287.610 -124.845 288.555 -124.810 ;
        RECT 292.645 -124.800 297.140 -124.775 ;
        RECT 292.645 -124.895 296.490 -124.800 ;
        RECT 285.415 -125.090 287.625 -125.015 ;
        RECT 285.415 -125.335 291.860 -125.090 ;
        RECT 277.455 -128.320 277.625 -125.360 ;
        RECT 285.465 -127.420 285.635 -125.335 ;
        RECT 286.445 -127.420 286.615 -125.335 ;
        RECT 287.425 -125.585 291.860 -125.335 ;
        RECT 292.675 -125.525 292.900 -124.895 ;
        RECT 293.650 -125.510 293.875 -124.895 ;
        RECT 287.425 -127.420 287.595 -125.585 ;
        RECT 288.510 -126.415 288.680 -125.585 ;
        RECT 289.490 -126.415 289.660 -125.585 ;
        RECT 290.470 -126.415 290.640 -125.585 ;
        RECT 291.450 -126.415 291.620 -125.585 ;
        RECT 292.700 -128.475 292.870 -125.525 ;
        RECT 293.680 -128.475 293.850 -125.510 ;
        RECT 295.760 -125.515 295.985 -124.895 ;
        RECT 296.745 -124.925 297.140 -124.800 ;
        RECT 297.995 -124.850 299.055 -124.155 ;
        RECT 310.845 -124.080 321.400 -123.525 ;
        RECT 323.500 -123.705 323.830 -117.200 ;
        RECT 310.845 -124.290 321.920 -124.080 ;
        RECT 323.415 -124.270 323.835 -123.705 ;
        RECT 325.180 -123.850 325.510 -117.200 ;
        RECT 339.665 -118.235 340.275 -106.425 ;
        RECT 356.650 -106.730 367.205 -106.425 ;
        RECT 372.045 -106.490 374.070 -106.170 ;
        RECT 369.230 -106.540 369.720 -106.525 ;
        RECT 372.045 -106.540 372.630 -106.490 ;
        RECT 356.650 -106.765 367.725 -106.730 ;
        RECT 368.090 -106.765 368.400 -106.625 ;
        RECT 356.650 -106.940 368.400 -106.765 ;
        RECT 358.660 -106.975 359.790 -106.940 ;
        RECT 358.845 -107.010 359.790 -106.975 ;
        RECT 363.880 -107.025 368.400 -106.940 ;
        RECT 363.880 -107.060 367.725 -107.025 ;
        RECT 356.650 -107.255 358.860 -107.180 ;
        RECT 356.650 -107.500 363.095 -107.255 ;
        RECT 356.700 -109.585 356.870 -107.500 ;
        RECT 357.680 -109.585 357.850 -107.500 ;
        RECT 358.660 -107.750 363.095 -107.500 ;
        RECT 363.910 -107.690 364.135 -107.060 ;
        RECT 364.885 -107.675 365.110 -107.060 ;
        RECT 358.660 -109.585 358.830 -107.750 ;
        RECT 359.745 -108.580 359.915 -107.750 ;
        RECT 360.725 -108.580 360.895 -107.750 ;
        RECT 361.705 -108.580 361.875 -107.750 ;
        RECT 362.685 -108.580 362.855 -107.750 ;
        RECT 363.935 -110.640 364.105 -107.690 ;
        RECT 364.915 -110.640 365.085 -107.675 ;
        RECT 366.995 -107.680 367.220 -107.060 ;
        RECT 368.090 -107.095 368.400 -107.025 ;
        RECT 369.230 -107.125 372.630 -106.540 ;
        RECT 373.880 -106.965 374.070 -106.490 ;
        RECT 374.865 -106.955 375.055 -106.170 ;
        RECT 369.230 -107.155 369.720 -107.125 ;
        RECT 367.030 -110.640 367.200 -107.680 ;
        RECT 373.895 -109.430 374.065 -106.965 ;
        RECT 374.875 -109.430 375.045 -106.955 ;
        RECT 377.825 -107.070 378.075 -106.170 ;
        RECT 378.455 -107.055 378.705 -106.170 ;
        RECT 379.610 -106.980 379.825 -106.170 ;
        RECT 380.595 -106.470 414.025 -106.170 ;
        RECT 418.865 -106.300 420.890 -105.980 ;
        RECT 416.050 -106.350 416.540 -106.335 ;
        RECT 418.865 -106.350 419.450 -106.300 ;
        RECT 380.595 -106.970 380.810 -106.470 ;
        RECT 377.850 -109.430 378.020 -107.070 ;
        RECT 378.500 -109.430 378.670 -107.055 ;
        RECT 379.640 -108.430 379.810 -106.980 ;
        RECT 380.620 -108.430 380.790 -106.970 ;
        RECT 369.265 -117.115 371.275 -116.785 ;
        RECT 339.665 -118.845 342.825 -118.235 ;
        RECT 329.365 -122.235 329.535 -120.905 ;
        RECT 330.345 -122.235 330.515 -120.905 ;
        RECT 331.325 -122.235 331.495 -120.905 ;
        RECT 332.305 -122.235 332.475 -120.905 ;
        RECT 329.125 -122.730 332.715 -122.235 ;
        RECT 330.035 -123.680 330.895 -122.730 ;
        RECT 334.230 -123.135 334.400 -121.050 ;
        RECT 335.210 -123.135 335.380 -121.050 ;
        RECT 336.190 -122.885 336.360 -121.050 ;
        RECT 337.275 -122.885 337.445 -122.055 ;
        RECT 338.255 -122.885 338.425 -122.055 ;
        RECT 339.235 -122.885 339.405 -122.055 ;
        RECT 340.215 -122.885 340.385 -122.055 ;
        RECT 336.190 -123.135 340.625 -122.885 ;
        RECT 334.180 -123.380 340.625 -123.135 ;
        RECT 334.180 -123.450 336.390 -123.380 ;
        RECT 334.175 -123.595 336.390 -123.450 ;
        RECT 334.175 -123.680 337.265 -123.595 ;
        RECT 329.185 -123.850 339.740 -123.680 ;
        RECT 342.215 -123.825 342.825 -118.845 ;
        RECT 356.790 -121.995 356.960 -120.665 ;
        RECT 357.770 -121.995 357.940 -120.665 ;
        RECT 358.750 -121.995 358.920 -120.665 ;
        RECT 359.730 -121.995 359.900 -120.665 ;
        RECT 356.550 -122.490 360.140 -121.995 ;
        RECT 357.460 -123.440 358.320 -122.490 ;
        RECT 361.655 -122.895 361.825 -120.810 ;
        RECT 362.635 -122.895 362.805 -120.810 ;
        RECT 363.615 -122.645 363.785 -120.810 ;
        RECT 364.700 -122.645 364.870 -121.815 ;
        RECT 365.680 -122.645 365.850 -121.815 ;
        RECT 366.660 -122.645 366.830 -121.815 ;
        RECT 367.640 -122.645 367.810 -121.815 ;
        RECT 363.615 -122.895 368.050 -122.645 ;
        RECT 361.605 -123.140 368.050 -122.895 ;
        RECT 361.605 -123.210 363.815 -123.140 ;
        RECT 361.600 -123.355 363.815 -123.210 ;
        RECT 361.600 -123.440 364.690 -123.355 ;
        RECT 325.180 -124.180 339.740 -123.850 ;
        RECT 340.515 -124.055 340.910 -123.900 ;
        RECT 329.185 -124.235 339.740 -124.180 ;
        RECT 340.015 -124.235 340.910 -124.055 ;
        RECT 312.855 -124.325 313.985 -124.290 ;
        RECT 313.040 -124.360 313.985 -124.325 ;
        RECT 318.075 -124.410 321.920 -124.290 ;
        RECT 310.845 -124.605 313.055 -124.530 ;
        RECT 310.845 -124.850 317.290 -124.605 ;
        RECT 297.995 -124.990 298.690 -124.850 ;
        RECT 295.795 -128.475 295.965 -125.515 ;
        RECT 310.895 -126.935 311.065 -124.850 ;
        RECT 311.875 -126.935 312.045 -124.850 ;
        RECT 312.855 -125.100 317.290 -124.850 ;
        RECT 318.105 -125.040 318.330 -124.410 ;
        RECT 319.080 -125.025 319.305 -124.410 ;
        RECT 312.855 -126.935 313.025 -125.100 ;
        RECT 313.940 -125.930 314.110 -125.100 ;
        RECT 314.920 -125.930 315.090 -125.100 ;
        RECT 315.900 -125.930 316.070 -125.100 ;
        RECT 316.880 -125.930 317.050 -125.100 ;
        RECT 318.130 -127.990 318.300 -125.040 ;
        RECT 319.110 -127.990 319.280 -125.025 ;
        RECT 321.190 -125.030 321.415 -124.410 ;
        RECT 329.185 -124.445 340.910 -124.235 ;
        RECT 331.195 -124.480 332.325 -124.445 ;
        RECT 331.380 -124.515 332.325 -124.480 ;
        RECT 336.415 -124.470 340.910 -124.445 ;
        RECT 336.415 -124.565 340.260 -124.470 ;
        RECT 329.185 -124.760 331.395 -124.685 ;
        RECT 329.185 -125.005 335.630 -124.760 ;
        RECT 321.225 -127.990 321.395 -125.030 ;
        RECT 329.235 -127.090 329.405 -125.005 ;
        RECT 330.215 -127.090 330.385 -125.005 ;
        RECT 331.195 -125.255 335.630 -125.005 ;
        RECT 336.445 -125.195 336.670 -124.565 ;
        RECT 337.420 -125.180 337.645 -124.565 ;
        RECT 331.195 -127.090 331.365 -125.255 ;
        RECT 332.280 -126.085 332.450 -125.255 ;
        RECT 333.260 -126.085 333.430 -125.255 ;
        RECT 334.240 -126.085 334.410 -125.255 ;
        RECT 335.220 -126.085 335.390 -125.255 ;
        RECT 336.470 -128.145 336.640 -125.195 ;
        RECT 337.450 -128.145 337.620 -125.180 ;
        RECT 339.530 -125.185 339.755 -124.565 ;
        RECT 340.515 -124.595 340.910 -124.470 ;
        RECT 341.765 -124.520 342.825 -123.825 ;
        RECT 356.610 -123.995 367.165 -123.440 ;
        RECT 369.265 -123.620 369.595 -117.115 ;
        RECT 356.610 -124.205 367.685 -123.995 ;
        RECT 369.180 -124.185 369.600 -123.620 ;
        RECT 370.945 -123.765 371.275 -117.115 ;
        RECT 385.430 -118.150 386.040 -106.470 ;
        RECT 403.470 -106.540 414.025 -106.470 ;
        RECT 403.470 -106.575 414.545 -106.540 ;
        RECT 414.910 -106.575 415.220 -106.435 ;
        RECT 403.470 -106.750 415.220 -106.575 ;
        RECT 405.480 -106.785 406.610 -106.750 ;
        RECT 405.665 -106.820 406.610 -106.785 ;
        RECT 410.700 -106.835 415.220 -106.750 ;
        RECT 410.700 -106.870 414.545 -106.835 ;
        RECT 403.470 -107.065 405.680 -106.990 ;
        RECT 403.470 -107.310 409.915 -107.065 ;
        RECT 403.520 -109.395 403.690 -107.310 ;
        RECT 404.500 -109.395 404.670 -107.310 ;
        RECT 405.480 -107.560 409.915 -107.310 ;
        RECT 410.730 -107.500 410.955 -106.870 ;
        RECT 411.705 -107.485 411.930 -106.870 ;
        RECT 405.480 -109.395 405.650 -107.560 ;
        RECT 406.565 -108.390 406.735 -107.560 ;
        RECT 407.545 -108.390 407.715 -107.560 ;
        RECT 408.525 -108.390 408.695 -107.560 ;
        RECT 409.505 -108.390 409.675 -107.560 ;
        RECT 410.755 -110.450 410.925 -107.500 ;
        RECT 411.735 -110.450 411.905 -107.485 ;
        RECT 413.815 -107.490 414.040 -106.870 ;
        RECT 414.910 -106.905 415.220 -106.835 ;
        RECT 416.050 -106.935 419.450 -106.350 ;
        RECT 420.700 -106.775 420.890 -106.300 ;
        RECT 421.685 -106.765 421.875 -105.980 ;
        RECT 416.050 -106.965 416.540 -106.935 ;
        RECT 413.850 -110.450 414.020 -107.490 ;
        RECT 420.715 -109.240 420.885 -106.775 ;
        RECT 421.695 -109.240 421.865 -106.765 ;
        RECT 424.645 -106.880 424.895 -105.980 ;
        RECT 425.275 -106.865 425.525 -105.980 ;
        RECT 426.430 -106.790 426.645 -105.980 ;
        RECT 427.415 -106.780 427.630 -105.980 ;
        RECT 424.670 -109.240 424.840 -106.880 ;
        RECT 425.320 -109.240 425.490 -106.865 ;
        RECT 426.460 -108.240 426.630 -106.790 ;
        RECT 427.440 -108.240 427.610 -106.780 ;
        RECT 416.085 -116.925 418.095 -116.595 ;
        RECT 385.430 -118.760 388.590 -118.150 ;
        RECT 375.130 -122.150 375.300 -120.820 ;
        RECT 376.110 -122.150 376.280 -120.820 ;
        RECT 377.090 -122.150 377.260 -120.820 ;
        RECT 378.070 -122.150 378.240 -120.820 ;
        RECT 374.890 -122.645 378.480 -122.150 ;
        RECT 375.800 -123.595 376.660 -122.645 ;
        RECT 379.995 -123.050 380.165 -120.965 ;
        RECT 380.975 -123.050 381.145 -120.965 ;
        RECT 381.955 -122.800 382.125 -120.965 ;
        RECT 383.040 -122.800 383.210 -121.970 ;
        RECT 384.020 -122.800 384.190 -121.970 ;
        RECT 385.000 -122.800 385.170 -121.970 ;
        RECT 385.980 -122.800 386.150 -121.970 ;
        RECT 381.955 -123.050 386.390 -122.800 ;
        RECT 379.945 -123.295 386.390 -123.050 ;
        RECT 379.945 -123.365 382.155 -123.295 ;
        RECT 379.940 -123.510 382.155 -123.365 ;
        RECT 379.940 -123.595 383.030 -123.510 ;
        RECT 374.950 -123.765 385.505 -123.595 ;
        RECT 387.980 -123.740 388.590 -118.760 ;
        RECT 403.610 -121.805 403.780 -120.475 ;
        RECT 404.590 -121.805 404.760 -120.475 ;
        RECT 405.570 -121.805 405.740 -120.475 ;
        RECT 406.550 -121.805 406.720 -120.475 ;
        RECT 403.370 -122.300 406.960 -121.805 ;
        RECT 404.280 -123.250 405.140 -122.300 ;
        RECT 408.475 -122.705 408.645 -120.620 ;
        RECT 409.455 -122.705 409.625 -120.620 ;
        RECT 410.435 -122.455 410.605 -120.620 ;
        RECT 411.520 -122.455 411.690 -121.625 ;
        RECT 412.500 -122.455 412.670 -121.625 ;
        RECT 413.480 -122.455 413.650 -121.625 ;
        RECT 414.460 -122.455 414.630 -121.625 ;
        RECT 410.435 -122.705 414.870 -122.455 ;
        RECT 408.425 -122.950 414.870 -122.705 ;
        RECT 408.425 -123.020 410.635 -122.950 ;
        RECT 408.420 -123.165 410.635 -123.020 ;
        RECT 408.420 -123.250 411.510 -123.165 ;
        RECT 370.945 -124.095 385.505 -123.765 ;
        RECT 386.280 -123.970 386.675 -123.815 ;
        RECT 374.950 -124.150 385.505 -124.095 ;
        RECT 385.780 -124.150 386.675 -123.970 ;
        RECT 358.620 -124.240 359.750 -124.205 ;
        RECT 358.805 -124.275 359.750 -124.240 ;
        RECT 363.840 -124.325 367.685 -124.205 ;
        RECT 356.610 -124.520 358.820 -124.445 ;
        RECT 341.765 -124.660 342.460 -124.520 ;
        RECT 356.610 -124.765 363.055 -124.520 ;
        RECT 339.565 -128.145 339.735 -125.185 ;
        RECT 356.660 -126.850 356.830 -124.765 ;
        RECT 357.640 -126.850 357.810 -124.765 ;
        RECT 358.620 -125.015 363.055 -124.765 ;
        RECT 363.870 -124.955 364.095 -124.325 ;
        RECT 364.845 -124.940 365.070 -124.325 ;
        RECT 358.620 -126.850 358.790 -125.015 ;
        RECT 359.705 -125.845 359.875 -125.015 ;
        RECT 360.685 -125.845 360.855 -125.015 ;
        RECT 361.665 -125.845 361.835 -125.015 ;
        RECT 362.645 -125.845 362.815 -125.015 ;
        RECT 363.895 -127.905 364.065 -124.955 ;
        RECT 364.875 -127.905 365.045 -124.940 ;
        RECT 366.955 -124.945 367.180 -124.325 ;
        RECT 374.950 -124.360 386.675 -124.150 ;
        RECT 376.960 -124.395 378.090 -124.360 ;
        RECT 377.145 -124.430 378.090 -124.395 ;
        RECT 382.180 -124.385 386.675 -124.360 ;
        RECT 382.180 -124.480 386.025 -124.385 ;
        RECT 374.950 -124.675 377.160 -124.600 ;
        RECT 374.950 -124.920 381.395 -124.675 ;
        RECT 366.990 -127.905 367.160 -124.945 ;
        RECT 375.000 -127.005 375.170 -124.920 ;
        RECT 375.980 -127.005 376.150 -124.920 ;
        RECT 376.960 -125.170 381.395 -124.920 ;
        RECT 382.210 -125.110 382.435 -124.480 ;
        RECT 383.185 -125.095 383.410 -124.480 ;
        RECT 376.960 -127.005 377.130 -125.170 ;
        RECT 378.045 -126.000 378.215 -125.170 ;
        RECT 379.025 -126.000 379.195 -125.170 ;
        RECT 380.005 -126.000 380.175 -125.170 ;
        RECT 380.985 -126.000 381.155 -125.170 ;
        RECT 382.235 -128.060 382.405 -125.110 ;
        RECT 383.215 -128.060 383.385 -125.095 ;
        RECT 385.295 -125.100 385.520 -124.480 ;
        RECT 386.280 -124.510 386.675 -124.385 ;
        RECT 387.530 -124.435 388.590 -123.740 ;
        RECT 403.430 -123.805 413.985 -123.250 ;
        RECT 416.085 -123.430 416.415 -116.925 ;
        RECT 403.430 -124.015 414.505 -123.805 ;
        RECT 416.000 -123.995 416.420 -123.430 ;
        RECT 417.765 -123.575 418.095 -116.925 ;
        RECT 432.250 -117.960 432.860 -105.975 ;
        RECT 432.250 -118.570 435.410 -117.960 ;
        RECT 421.950 -121.960 422.120 -120.630 ;
        RECT 422.930 -121.960 423.100 -120.630 ;
        RECT 423.910 -121.960 424.080 -120.630 ;
        RECT 424.890 -121.960 425.060 -120.630 ;
        RECT 421.710 -122.455 425.300 -121.960 ;
        RECT 422.620 -123.405 423.480 -122.455 ;
        RECT 426.815 -122.860 426.985 -120.775 ;
        RECT 427.795 -122.860 427.965 -120.775 ;
        RECT 428.775 -122.610 428.945 -120.775 ;
        RECT 429.860 -122.610 430.030 -121.780 ;
        RECT 430.840 -122.610 431.010 -121.780 ;
        RECT 431.820 -122.610 431.990 -121.780 ;
        RECT 432.800 -122.610 432.970 -121.780 ;
        RECT 428.775 -122.860 433.210 -122.610 ;
        RECT 426.765 -123.105 433.210 -122.860 ;
        RECT 426.765 -123.175 428.975 -123.105 ;
        RECT 426.760 -123.320 428.975 -123.175 ;
        RECT 426.760 -123.405 429.850 -123.320 ;
        RECT 421.770 -123.575 432.325 -123.405 ;
        RECT 434.800 -123.550 435.410 -118.570 ;
        RECT 417.765 -123.905 432.325 -123.575 ;
        RECT 433.100 -123.780 433.495 -123.625 ;
        RECT 421.770 -123.960 432.325 -123.905 ;
        RECT 432.600 -123.960 433.495 -123.780 ;
        RECT 405.440 -124.050 406.570 -124.015 ;
        RECT 405.625 -124.085 406.570 -124.050 ;
        RECT 410.660 -124.135 414.505 -124.015 ;
        RECT 403.430 -124.330 405.640 -124.255 ;
        RECT 387.530 -124.575 388.225 -124.435 ;
        RECT 403.430 -124.575 409.875 -124.330 ;
        RECT 385.330 -128.060 385.500 -125.100 ;
        RECT 403.480 -126.660 403.650 -124.575 ;
        RECT 404.460 -126.660 404.630 -124.575 ;
        RECT 405.440 -124.825 409.875 -124.575 ;
        RECT 410.690 -124.765 410.915 -124.135 ;
        RECT 411.665 -124.750 411.890 -124.135 ;
        RECT 405.440 -126.660 405.610 -124.825 ;
        RECT 406.525 -125.655 406.695 -124.825 ;
        RECT 407.505 -125.655 407.675 -124.825 ;
        RECT 408.485 -125.655 408.655 -124.825 ;
        RECT 409.465 -125.655 409.635 -124.825 ;
        RECT 410.715 -127.715 410.885 -124.765 ;
        RECT 411.695 -127.715 411.865 -124.750 ;
        RECT 413.775 -124.755 414.000 -124.135 ;
        RECT 421.770 -124.170 433.495 -123.960 ;
        RECT 423.780 -124.205 424.910 -124.170 ;
        RECT 423.965 -124.240 424.910 -124.205 ;
        RECT 429.000 -124.195 433.495 -124.170 ;
        RECT 429.000 -124.290 432.845 -124.195 ;
        RECT 421.770 -124.485 423.980 -124.410 ;
        RECT 421.770 -124.730 428.215 -124.485 ;
        RECT 413.810 -127.715 413.980 -124.755 ;
        RECT 421.820 -126.815 421.990 -124.730 ;
        RECT 422.800 -126.815 422.970 -124.730 ;
        RECT 423.780 -124.980 428.215 -124.730 ;
        RECT 429.030 -124.920 429.255 -124.290 ;
        RECT 430.005 -124.905 430.230 -124.290 ;
        RECT 423.780 -126.815 423.950 -124.980 ;
        RECT 424.865 -125.810 425.035 -124.980 ;
        RECT 425.845 -125.810 426.015 -124.980 ;
        RECT 426.825 -125.810 426.995 -124.980 ;
        RECT 427.805 -125.810 427.975 -124.980 ;
        RECT 429.055 -127.870 429.225 -124.920 ;
        RECT 430.035 -127.870 430.205 -124.905 ;
        RECT 432.115 -124.910 432.340 -124.290 ;
        RECT 433.100 -124.320 433.495 -124.195 ;
        RECT 434.350 -124.245 435.410 -123.550 ;
        RECT 434.350 -124.385 435.045 -124.245 ;
        RECT 432.150 -127.870 432.320 -124.910 ;
        RECT 61.985 -136.350 70.995 -136.325 ;
        RECT 75.485 -136.350 83.350 -136.325 ;
        RECT 36.685 -137.245 36.915 -136.635 ;
        RECT 57.225 -136.665 83.350 -136.350 ;
        RECT 5.975 -137.780 8.940 -137.590 ;
        RECT 18.040 -137.780 21.005 -137.590 ;
        RECT 31.655 -137.780 36.915 -137.245 ;
        RECT -113.875 -137.955 -100.865 -137.910 ;
        RECT -37.670 -138.745 37.140 -137.780 ;
        RECT 479.145 -141.695 493.990 -79.080 ;
        RECT 416.665 -156.540 493.990 -141.695 ;
        RECT 416.665 -163.245 431.510 -156.540 ;
        RECT 129.615 -164.350 435.355 -163.245 ;
        RECT 34.475 -168.160 435.355 -164.350 ;
        RECT -127.845 -170.685 -127.605 -169.855 ;
        RECT -130.080 -170.855 -127.605 -170.685 ;
        RECT -127.845 -171.865 -127.605 -170.855 ;
        RECT -130.080 -172.035 -127.605 -171.865 ;
        RECT -127.845 -173.045 -127.605 -172.035 ;
        RECT -130.080 -173.215 -127.605 -173.045 ;
        RECT -127.845 -174.225 -127.605 -173.215 ;
        RECT -130.080 -174.395 -127.605 -174.225 ;
        RECT -127.845 -175.345 -127.605 -174.395 ;
        RECT -127.245 -175.345 -126.915 -170.405 ;
        RECT 34.475 -173.930 38.285 -168.160 ;
        RECT 129.615 -168.760 435.355 -168.160 ;
        RECT -36.670 -173.985 40.630 -173.930 ;
        RECT -48.325 -174.165 40.630 -173.985 ;
        RECT -127.845 -175.405 -126.915 -175.345 ;
        RECT -130.080 -175.575 -126.915 -175.405 ;
        RECT -127.845 -175.640 -126.915 -175.575 ;
        RECT -127.845 -176.585 -127.605 -175.640 ;
        RECT -130.080 -176.755 -127.605 -176.585 ;
        RECT -127.845 -177.730 -127.605 -176.755 ;
        RECT -127.245 -177.300 -126.915 -175.640 ;
        RECT -73.450 -174.430 40.630 -174.165 ;
        RECT -73.450 -174.480 -47.325 -174.430 ;
        RECT -73.450 -174.505 -65.585 -174.480 ;
        RECT -61.095 -174.505 -52.085 -174.480 ;
        RECT -73.450 -177.300 -73.005 -174.505 ;
        RECT -72.205 -175.960 -72.035 -174.505 ;
        RECT -71.225 -175.960 -71.055 -174.505 ;
        RECT -70.245 -175.960 -70.075 -174.505 ;
        RECT -68.020 -175.960 -67.850 -174.505 ;
        RECT -67.040 -175.960 -66.870 -174.505 ;
        RECT -66.060 -175.960 -65.890 -174.505 ;
        RECT -58.705 -175.960 -58.535 -174.505 ;
        RECT -57.725 -175.960 -57.555 -174.505 ;
        RECT -56.745 -175.960 -56.575 -174.505 ;
        RECT -54.520 -175.960 -54.350 -174.505 ;
        RECT -53.540 -175.960 -53.370 -174.505 ;
        RECT -52.560 -175.960 -52.390 -174.505 ;
        RECT -40.415 -175.050 -40.190 -174.430 ;
        RECT -38.305 -175.045 -38.080 -174.430 ;
        RECT -127.245 -177.730 -73.005 -177.300 ;
        RECT -127.845 -177.765 -73.005 -177.730 ;
        RECT -130.080 -177.935 -73.005 -177.765 ;
        RECT -127.845 -178.025 -73.005 -177.935 ;
        RECT -40.395 -178.010 -40.225 -175.050 ;
        RECT -38.280 -178.010 -38.110 -175.045 ;
        RECT -37.330 -175.060 -37.105 -174.430 ;
        RECT -36.680 -174.895 40.630 -174.430 ;
        RECT -37.300 -178.010 -37.130 -175.060 ;
        RECT -29.855 -175.430 -24.595 -174.895 ;
        RECT -29.855 -176.075 -29.655 -175.430 ;
        RECT -28.910 -176.075 -28.680 -175.430 ;
        RECT -27.920 -176.055 -27.690 -175.430 ;
        RECT -29.855 -176.990 -29.685 -176.075 ;
        RECT -28.875 -176.990 -28.705 -176.075 ;
        RECT -27.895 -176.990 -27.725 -176.055 ;
        RECT -27.355 -176.075 -27.125 -175.430 ;
        RECT -26.375 -176.050 -26.145 -175.430 ;
        RECT -27.325 -176.990 -27.155 -176.075 ;
        RECT -26.345 -176.990 -26.175 -176.050 ;
        RECT -25.810 -176.100 -25.580 -175.430 ;
        RECT -24.825 -176.040 -24.595 -175.430 ;
        RECT -25.780 -176.990 -25.610 -176.100 ;
        RECT -24.800 -176.990 -24.630 -176.040 ;
        RECT -127.845 -178.885 -127.605 -178.025 ;
        RECT -127.245 -178.365 -73.005 -178.025 ;
        RECT -127.245 -178.415 -107.090 -178.365 ;
        RECT -127.245 -178.660 -116.905 -178.415 ;
        RECT -127.245 -178.885 -126.915 -178.660 ;
        RECT -127.845 -178.945 -126.915 -178.885 ;
        RECT -130.080 -179.115 -126.915 -178.945 ;
        RECT -127.845 -179.180 -126.915 -179.115 ;
        RECT -127.845 -180.065 -127.605 -179.180 ;
        RECT -127.245 -180.065 -126.915 -179.180 ;
        RECT -127.845 -180.125 -126.915 -180.065 ;
        RECT -130.080 -180.295 -126.915 -180.125 ;
        RECT -127.845 -180.360 -126.915 -180.295 ;
        RECT -127.845 -181.255 -127.605 -180.360 ;
        RECT -127.245 -181.255 -126.915 -180.360 ;
        RECT -127.845 -181.300 -126.915 -181.255 ;
        RECT -118.265 -181.300 -116.905 -178.660 ;
        RECT -110.200 -179.895 -110.030 -178.415 ;
        RECT -109.220 -179.895 -109.050 -178.415 ;
        RECT -108.240 -179.895 -108.070 -178.415 ;
        RECT -107.260 -179.895 -107.090 -178.415 ;
        RECT -104.575 -178.435 -103.350 -178.365 ;
        RECT -104.550 -179.895 -104.380 -178.435 ;
        RECT -103.570 -179.895 -103.400 -178.435 ;
        RECT -100.465 -178.675 -93.830 -178.365 ;
        RECT -100.465 -178.950 -93.810 -178.675 ;
        RECT -100.205 -181.005 -100.035 -178.950 ;
        RECT -99.225 -181.005 -99.055 -178.950 ;
        RECT -98.245 -179.170 -93.810 -178.950 ;
        RECT -98.245 -181.005 -98.075 -179.170 ;
        RECT -97.160 -180.000 -96.990 -179.170 ;
        RECT -96.180 -180.000 -96.010 -179.170 ;
        RECT -95.200 -180.000 -95.030 -179.170 ;
        RECT -94.220 -180.000 -94.050 -179.170 ;
        RECT -127.845 -181.305 -116.905 -181.300 ;
        RECT -130.080 -181.475 -116.905 -181.305 ;
        RECT -127.845 -181.550 -116.905 -181.475 ;
        RECT -127.845 -182.455 -127.605 -181.550 ;
        RECT -127.245 -182.455 -116.905 -181.550 ;
        RECT -127.845 -182.485 -116.905 -182.455 ;
        RECT -130.080 -182.655 -116.905 -182.485 ;
        RECT -127.845 -182.660 -116.905 -182.655 ;
        RECT -127.845 -182.750 -126.915 -182.660 ;
        RECT -127.845 -183.605 -127.605 -182.750 ;
        RECT -127.245 -183.605 -126.915 -182.750 ;
        RECT -127.845 -183.665 -126.915 -183.605 ;
        RECT -130.080 -183.835 -126.915 -183.665 ;
        RECT -127.845 -183.900 -126.915 -183.835 ;
        RECT -127.845 -184.790 -127.605 -183.900 ;
        RECT -127.245 -184.790 -126.915 -183.900 ;
        RECT -127.845 -184.845 -126.915 -184.790 ;
        RECT -130.080 -185.015 -126.915 -184.845 ;
        RECT -127.845 -185.085 -126.915 -185.015 ;
        RECT -127.845 -185.960 -127.605 -185.085 ;
        RECT -127.245 -185.960 -126.915 -185.085 ;
        RECT -127.845 -186.025 -126.915 -185.960 ;
        RECT -130.080 -186.195 -126.915 -186.025 ;
        RECT -127.845 -186.255 -126.915 -186.195 ;
        RECT -127.845 -187.130 -127.605 -186.255 ;
        RECT -127.245 -186.605 -126.915 -186.255 ;
        RECT -118.265 -186.605 -116.905 -182.660 ;
        RECT -73.450 -182.980 -73.005 -178.365 ;
        RECT -23.220 -179.080 -22.645 -174.895 ;
        RECT -15.785 -175.085 -12.820 -174.895 ;
        RECT -17.355 -175.430 -12.095 -175.085 ;
        RECT -17.355 -176.075 -17.155 -175.430 ;
        RECT -16.410 -176.075 -16.180 -175.430 ;
        RECT -15.420 -176.055 -15.190 -175.430 ;
        RECT -17.355 -176.990 -17.185 -176.075 ;
        RECT -16.375 -176.990 -16.205 -176.075 ;
        RECT -15.395 -176.990 -15.225 -176.055 ;
        RECT -14.855 -176.075 -14.625 -175.430 ;
        RECT -13.875 -176.050 -13.645 -175.430 ;
        RECT -14.825 -176.990 -14.655 -176.075 ;
        RECT -13.845 -176.990 -13.675 -176.050 ;
        RECT -13.310 -176.100 -13.080 -175.430 ;
        RECT -12.325 -176.040 -12.095 -175.430 ;
        RECT -13.280 -176.990 -13.110 -176.100 ;
        RECT -12.300 -176.990 -12.130 -176.040 ;
        RECT -23.245 -179.760 -22.630 -179.080 ;
        RECT -10.380 -179.255 -9.810 -174.895 ;
        RECT -3.205 -175.085 -0.240 -174.895 ;
        RECT -4.855 -175.430 0.405 -175.085 ;
        RECT -4.855 -176.075 -4.655 -175.430 ;
        RECT -3.910 -176.075 -3.680 -175.430 ;
        RECT -2.920 -176.055 -2.690 -175.430 ;
        RECT -4.855 -176.990 -4.685 -176.075 ;
        RECT -3.875 -176.990 -3.705 -176.075 ;
        RECT -2.895 -176.990 -2.725 -176.055 ;
        RECT -2.355 -176.075 -2.125 -175.430 ;
        RECT -1.375 -176.050 -1.145 -175.430 ;
        RECT -2.325 -176.990 -2.155 -176.075 ;
        RECT -1.345 -176.990 -1.175 -176.050 ;
        RECT -0.810 -176.100 -0.580 -175.430 ;
        RECT 0.175 -176.040 0.405 -175.430 ;
        RECT -0.780 -176.990 -0.610 -176.100 ;
        RECT 0.200 -176.990 0.370 -176.040 ;
        RECT 2.030 -179.255 2.605 -174.895 ;
        RECT 9.465 -175.085 12.430 -174.895 ;
        RECT 21.530 -175.085 24.495 -174.895 ;
        RECT 7.645 -175.430 12.905 -175.085 ;
        RECT 7.645 -176.075 7.845 -175.430 ;
        RECT 8.590 -176.075 8.820 -175.430 ;
        RECT 9.580 -176.055 9.810 -175.430 ;
        RECT 7.645 -176.990 7.815 -176.075 ;
        RECT 8.625 -176.990 8.795 -176.075 ;
        RECT 9.605 -176.990 9.775 -176.055 ;
        RECT 10.145 -176.075 10.375 -175.430 ;
        RECT 11.125 -176.050 11.355 -175.430 ;
        RECT 10.175 -176.990 10.345 -176.075 ;
        RECT 11.155 -176.990 11.325 -176.050 ;
        RECT 11.690 -176.100 11.920 -175.430 ;
        RECT 12.675 -176.040 12.905 -175.430 ;
        RECT 20.145 -175.430 25.405 -175.085 ;
        RECT 11.720 -176.990 11.890 -176.100 ;
        RECT 12.700 -176.990 12.870 -176.040 ;
        RECT 20.145 -176.075 20.345 -175.430 ;
        RECT 21.090 -176.075 21.320 -175.430 ;
        RECT 22.080 -176.055 22.310 -175.430 ;
        RECT 20.145 -176.990 20.315 -176.075 ;
        RECT 21.125 -176.990 21.295 -176.075 ;
        RECT 22.105 -176.990 22.275 -176.055 ;
        RECT 22.645 -176.075 22.875 -175.430 ;
        RECT 23.625 -176.050 23.855 -175.430 ;
        RECT 22.675 -176.990 22.845 -176.075 ;
        RECT 23.655 -176.990 23.825 -176.050 ;
        RECT 24.190 -176.100 24.420 -175.430 ;
        RECT 25.175 -176.040 25.405 -175.430 ;
        RECT 35.145 -175.430 40.405 -174.895 ;
        RECT 24.220 -176.990 24.390 -176.100 ;
        RECT 25.200 -176.990 25.370 -176.040 ;
        RECT 35.145 -176.075 35.345 -175.430 ;
        RECT 36.090 -176.075 36.320 -175.430 ;
        RECT 37.080 -176.055 37.310 -175.430 ;
        RECT 35.145 -176.990 35.315 -176.075 ;
        RECT 36.125 -176.990 36.295 -176.075 ;
        RECT 37.105 -176.990 37.275 -176.055 ;
        RECT 37.645 -176.075 37.875 -175.430 ;
        RECT 38.625 -176.050 38.855 -175.430 ;
        RECT 37.675 -176.990 37.845 -176.075 ;
        RECT 38.655 -176.990 38.825 -176.050 ;
        RECT 39.190 -176.100 39.420 -175.430 ;
        RECT 40.175 -176.040 40.405 -175.430 ;
        RECT 129.615 -175.705 135.130 -168.760 ;
        RECT 39.220 -176.990 39.390 -176.100 ;
        RECT 40.200 -176.990 40.370 -176.040 ;
        RECT -10.410 -179.935 -9.795 -179.255 ;
        RECT 2.005 -179.935 2.620 -179.255 ;
        RECT -71.715 -182.965 -71.545 -181.510 ;
        RECT -70.735 -182.965 -70.565 -181.510 ;
        RECT -69.755 -182.965 -69.585 -181.510 ;
        RECT -63.000 -182.965 -62.830 -181.510 ;
        RECT -62.020 -182.965 -61.850 -181.510 ;
        RECT -61.040 -182.965 -60.870 -181.510 ;
        RECT -58.215 -182.965 -58.045 -181.510 ;
        RECT -57.235 -182.965 -57.065 -181.510 ;
        RECT -56.255 -182.965 -56.085 -181.510 ;
        RECT -49.500 -182.965 -49.330 -181.510 ;
        RECT -48.520 -182.965 -48.350 -181.510 ;
        RECT -47.540 -182.965 -47.370 -181.510 ;
        RECT -45.090 -182.965 -44.920 -181.510 ;
        RECT -44.110 -182.965 -43.940 -181.510 ;
        RECT -43.130 -182.965 -42.960 -181.510 ;
        RECT 2.000 -182.025 2.615 -182.020 ;
        RECT -72.015 -182.980 -69.540 -182.965 ;
        RECT -63.305 -182.970 -56.040 -182.965 ;
        RECT -73.450 -182.990 -67.930 -182.980 ;
        RECT -63.305 -182.990 -54.475 -182.970 ;
        RECT -49.805 -182.990 -42.915 -182.965 ;
        RECT -92.025 -186.360 -91.855 -184.275 ;
        RECT -91.045 -186.360 -90.875 -184.275 ;
        RECT -90.065 -186.110 -89.895 -184.275 ;
        RECT -88.980 -186.110 -88.810 -185.280 ;
        RECT -88.000 -186.110 -87.830 -185.280 ;
        RECT -87.020 -186.110 -86.850 -185.280 ;
        RECT -86.040 -186.110 -85.870 -185.280 ;
        RECT -90.065 -186.360 -85.630 -186.110 ;
        RECT -84.790 -186.170 -84.620 -183.220 ;
        RECT -127.245 -187.120 -116.905 -186.605 ;
        RECT -92.075 -186.605 -85.630 -186.360 ;
        RECT -92.075 -186.680 -89.865 -186.605 ;
        RECT -84.815 -186.800 -84.590 -186.170 ;
        RECT -83.810 -186.185 -83.640 -183.220 ;
        RECT -81.695 -186.180 -81.525 -183.220 ;
        RECT -73.450 -183.305 -42.915 -182.990 ;
        RECT -73.450 -183.320 -67.930 -183.305 ;
        RECT -56.840 -183.310 -54.475 -183.305 ;
        RECT -83.840 -186.800 -83.615 -186.185 ;
        RECT -81.730 -186.800 -81.505 -186.180 ;
        RECT -89.880 -186.885 -88.935 -186.850 ;
        RECT -90.065 -186.920 -88.935 -186.885 ;
        RECT -84.845 -186.920 -81.000 -186.800 ;
        RECT -92.075 -187.120 -81.000 -186.920 ;
        RECT -127.245 -187.130 -81.000 -187.120 ;
        RECT -127.845 -187.205 -81.520 -187.130 ;
        RECT -130.080 -187.375 -81.520 -187.205 ;
        RECT -127.845 -187.425 -81.520 -187.375 ;
        RECT -127.845 -188.385 -127.605 -187.425 ;
        RECT -130.080 -188.555 -127.605 -188.385 ;
        RECT -127.845 -189.625 -127.605 -188.555 ;
        RECT -130.080 -189.795 -127.605 -189.625 ;
        RECT -127.845 -190.755 -127.605 -189.795 ;
        RECT -127.245 -187.685 -81.520 -187.425 ;
        RECT -127.245 -187.965 -94.200 -187.685 ;
        RECT -127.245 -190.755 -126.915 -187.965 ;
        RECT -118.265 -188.115 -94.200 -187.965 ;
        RECT -118.265 -188.280 -94.250 -188.115 ;
        RECT -109.965 -188.465 -103.520 -188.280 ;
        RECT -109.915 -190.550 -109.745 -188.465 ;
        RECT -108.935 -190.550 -108.765 -188.465 ;
        RECT -107.955 -188.715 -103.520 -188.465 ;
        RECT -107.955 -190.550 -107.785 -188.715 ;
        RECT -106.870 -189.545 -106.700 -188.715 ;
        RECT -105.890 -189.545 -105.720 -188.715 ;
        RECT -104.910 -189.545 -104.740 -188.715 ;
        RECT -103.930 -189.545 -103.760 -188.715 ;
        RECT -101.050 -189.575 -100.880 -188.280 ;
        RECT -100.070 -189.575 -99.900 -188.280 ;
        RECT -99.090 -189.575 -98.920 -188.280 ;
        RECT -98.110 -189.575 -97.940 -188.280 ;
        RECT -95.400 -189.575 -95.230 -188.280 ;
        RECT -94.420 -189.575 -94.250 -188.280 ;
        RECT -91.225 -188.635 -90.365 -187.685 ;
        RECT -87.085 -187.770 -83.995 -187.685 ;
        RECT -87.085 -187.915 -84.870 -187.770 ;
        RECT -87.080 -187.985 -84.870 -187.915 ;
        RECT -87.080 -188.230 -80.635 -187.985 ;
        RECT -92.135 -189.130 -88.545 -188.635 ;
        RECT -91.895 -190.460 -91.725 -189.130 ;
        RECT -90.915 -190.460 -90.745 -189.130 ;
        RECT -89.935 -190.460 -89.765 -189.130 ;
        RECT -88.955 -190.460 -88.785 -189.130 ;
        RECT -87.030 -190.315 -86.860 -188.230 ;
        RECT -86.050 -190.315 -85.880 -188.230 ;
        RECT -85.070 -188.480 -80.635 -188.230 ;
        RECT -85.070 -190.315 -84.900 -188.480 ;
        RECT -83.985 -189.310 -83.815 -188.480 ;
        RECT -83.005 -189.310 -82.835 -188.480 ;
        RECT -82.025 -189.310 -81.855 -188.480 ;
        RECT -81.045 -189.310 -80.875 -188.480 ;
        RECT -127.845 -190.805 -126.915 -190.755 ;
        RECT -130.080 -190.975 -126.915 -190.805 ;
        RECT -127.845 -191.050 -126.915 -190.975 ;
        RECT -127.845 -191.910 -127.605 -191.050 ;
        RECT -127.245 -191.910 -126.915 -191.050 ;
        RECT -127.845 -191.985 -126.915 -191.910 ;
        RECT -130.080 -192.155 -126.915 -191.985 ;
        RECT -127.845 -192.205 -126.915 -192.155 ;
        RECT -127.845 -193.090 -127.605 -192.205 ;
        RECT -127.245 -193.090 -126.915 -192.205 ;
        RECT -127.845 -193.165 -126.915 -193.090 ;
        RECT -130.080 -193.335 -126.915 -193.165 ;
        RECT -127.845 -193.385 -126.915 -193.335 ;
        RECT -127.845 -194.265 -127.605 -193.385 ;
        RECT -127.245 -194.265 -126.915 -193.385 ;
        RECT -127.845 -194.345 -126.915 -194.265 ;
        RECT -130.080 -194.515 -126.915 -194.345 ;
        RECT -127.845 -194.560 -126.915 -194.515 ;
        RECT -127.845 -195.460 -127.605 -194.560 ;
        RECT -127.245 -195.460 -126.915 -194.560 ;
        RECT -127.845 -195.525 -126.915 -195.460 ;
        RECT -130.080 -195.695 -126.915 -195.525 ;
        RECT -127.845 -195.755 -126.915 -195.695 ;
        RECT -127.845 -196.605 -127.605 -195.755 ;
        RECT -127.245 -196.605 -126.915 -195.755 ;
        RECT -127.845 -196.705 -126.915 -196.605 ;
        RECT -130.080 -196.875 -126.915 -196.705 ;
        RECT -127.845 -196.900 -126.915 -196.875 ;
        RECT -127.845 -197.885 -127.605 -196.900 ;
        RECT -130.080 -198.055 -127.605 -197.885 ;
        RECT -127.845 -199.065 -127.605 -198.055 ;
        RECT -130.080 -199.235 -127.605 -199.065 ;
        RECT -127.845 -199.635 -127.605 -199.235 ;
        RECT -127.245 -199.635 -126.915 -196.900 ;
        RECT -71.140 -191.800 -70.375 -183.320 ;
        RECT -31.550 -184.050 -31.380 -182.595 ;
        RECT -30.570 -184.050 -30.400 -182.595 ;
        RECT -29.590 -184.050 -29.420 -182.595 ;
        RECT -10.415 -182.875 -9.800 -182.195 ;
        RECT 2.000 -182.335 3.530 -182.025 ;
        RECT -23.250 -183.595 -22.635 -182.915 ;
        RECT -31.595 -184.390 -29.120 -184.050 ;
        RECT -31.515 -186.340 -31.075 -184.390 ;
        RECT -30.600 -186.340 -30.160 -184.390 ;
        RECT -29.690 -186.340 -29.250 -184.390 ;
        RECT -34.080 -186.355 -28.560 -186.340 ;
        RECT -23.225 -186.355 -22.650 -183.595 ;
        RECT -17.470 -186.355 -15.105 -186.350 ;
        RECT -10.395 -186.355 -9.820 -182.875 ;
        RECT -4.120 -186.355 -3.505 -186.245 ;
        RECT -34.080 -186.670 -3.505 -186.355 ;
        RECT -34.080 -186.680 -28.560 -186.670 ;
        RECT -67.080 -191.240 -66.910 -189.155 ;
        RECT -66.100 -191.240 -65.930 -189.155 ;
        RECT -65.120 -190.990 -64.950 -189.155 ;
        RECT -64.035 -190.990 -63.865 -190.160 ;
        RECT -63.055 -190.990 -62.885 -190.160 ;
        RECT -62.075 -190.990 -61.905 -190.160 ;
        RECT -61.095 -190.990 -60.925 -190.160 ;
        RECT -65.120 -191.240 -60.685 -190.990 ;
        RECT -59.845 -191.050 -59.675 -188.100 ;
        RECT -67.130 -191.485 -60.685 -191.240 ;
        RECT -67.130 -191.560 -64.920 -191.485 ;
        RECT -59.870 -191.680 -59.645 -191.050 ;
        RECT -58.865 -191.065 -58.695 -188.100 ;
        RECT -56.750 -191.060 -56.580 -188.100 ;
        RECT -58.895 -191.680 -58.670 -191.065 ;
        RECT -56.785 -191.680 -56.560 -191.060 ;
        RECT -64.935 -191.765 -63.990 -191.730 ;
        RECT -65.120 -191.800 -63.990 -191.765 ;
        RECT -59.900 -191.800 -56.055 -191.680 ;
        RECT -71.140 -192.010 -56.055 -191.800 ;
        RECT -71.140 -192.565 -56.575 -192.010 ;
        RECT -71.140 -198.800 -70.375 -192.565 ;
        RECT -66.280 -193.515 -65.420 -192.565 ;
        RECT -62.140 -192.650 -59.050 -192.565 ;
        RECT -62.140 -192.795 -59.925 -192.650 ;
        RECT -62.135 -192.865 -59.925 -192.795 ;
        RECT -62.135 -193.110 -55.690 -192.865 ;
        RECT -67.190 -194.010 -63.600 -193.515 ;
        RECT -66.950 -195.340 -66.780 -194.010 ;
        RECT -65.970 -195.340 -65.800 -194.010 ;
        RECT -64.990 -195.340 -64.820 -194.010 ;
        RECT -64.010 -195.340 -63.840 -194.010 ;
        RECT -62.085 -195.195 -61.915 -193.110 ;
        RECT -61.105 -195.195 -60.935 -193.110 ;
        RECT -60.125 -193.360 -55.690 -193.110 ;
        RECT -60.125 -195.195 -59.955 -193.360 ;
        RECT -59.040 -194.190 -58.870 -193.360 ;
        RECT -58.060 -194.190 -57.890 -193.360 ;
        RECT -57.080 -194.190 -56.910 -193.360 ;
        RECT -56.100 -194.190 -55.930 -193.360 ;
        RECT -34.080 -195.155 -33.635 -186.680 ;
        RECT -32.645 -186.695 -30.170 -186.680 ;
        RECT -23.935 -186.690 -15.105 -186.670 ;
        RECT -23.935 -186.695 -16.670 -186.690 ;
        RECT -10.435 -186.695 -3.505 -186.670 ;
        RECT -32.345 -188.150 -32.175 -186.695 ;
        RECT -31.365 -188.150 -31.195 -186.695 ;
        RECT -30.385 -188.150 -30.215 -186.695 ;
        RECT -23.630 -188.150 -23.460 -186.695 ;
        RECT -22.650 -188.150 -22.480 -186.695 ;
        RECT -21.670 -188.150 -21.500 -186.695 ;
        RECT -18.845 -188.150 -18.675 -186.695 ;
        RECT -17.865 -188.150 -17.695 -186.695 ;
        RECT -16.885 -188.150 -16.715 -186.695 ;
        RECT -10.130 -188.150 -9.960 -186.695 ;
        RECT -9.150 -188.150 -8.980 -186.695 ;
        RECT -8.170 -188.150 -8.000 -186.695 ;
        RECT -5.720 -188.150 -5.550 -186.695 ;
        RECT -4.740 -188.150 -4.570 -186.695 ;
        RECT -4.120 -186.925 -3.505 -186.695 ;
        RECT -2.650 -186.375 -2.035 -186.240 ;
        RECT 2.025 -186.375 2.600 -182.335 ;
        RECT 12.240 -186.375 12.855 -186.305 ;
        RECT -2.650 -186.770 12.855 -186.375 ;
        RECT -2.650 -186.775 -0.875 -186.770 ;
        RECT -2.650 -186.920 -1.880 -186.775 ;
        RECT -3.760 -188.150 -3.590 -186.925 ;
        RECT -2.050 -188.235 -1.880 -186.920 ;
        RECT -1.070 -188.235 -0.900 -186.775 ;
        RECT 1.640 -188.235 1.810 -186.770 ;
        RECT 2.620 -188.235 2.790 -186.770 ;
        RECT 3.600 -188.235 3.770 -186.770 ;
        RECT 4.580 -188.235 4.750 -186.770 ;
        RECT 6.375 -186.970 10.810 -186.770 ;
        RECT 6.615 -187.800 6.785 -186.970 ;
        RECT 7.595 -187.800 7.765 -186.970 ;
        RECT 8.575 -187.800 8.745 -186.970 ;
        RECT 9.555 -187.800 9.725 -186.970 ;
        RECT 10.640 -188.805 10.810 -186.970 ;
        RECT 11.620 -188.805 11.790 -186.770 ;
        RECT 12.240 -186.985 12.855 -186.770 ;
        RECT 14.185 -186.485 14.800 -186.300 ;
        RECT 20.325 -186.410 20.940 -186.185 ;
        RECT 18.635 -186.485 20.940 -186.410 ;
        RECT 14.185 -186.730 20.940 -186.485 ;
        RECT 14.185 -186.980 18.835 -186.730 ;
        RECT 12.600 -188.805 12.770 -186.985 ;
        RECT 14.640 -187.810 14.810 -186.980 ;
        RECT 15.620 -187.810 15.790 -186.980 ;
        RECT 16.600 -187.810 16.770 -186.980 ;
        RECT 17.580 -187.810 17.750 -186.980 ;
        RECT 18.665 -188.815 18.835 -186.980 ;
        RECT 19.645 -188.815 19.815 -186.730 ;
        RECT 20.325 -186.865 20.940 -186.730 ;
        RECT 22.330 -186.340 22.945 -186.175 ;
        RECT 22.330 -186.365 26.810 -186.340 ;
        RECT 29.110 -186.365 29.725 -186.200 ;
        RECT 22.330 -186.705 29.725 -186.365 ;
        RECT 22.330 -186.730 23.935 -186.705 ;
        RECT 26.450 -186.710 29.725 -186.705 ;
        RECT 22.330 -186.855 22.945 -186.730 ;
        RECT 20.625 -188.815 20.795 -186.865 ;
        RECT 22.760 -188.190 22.930 -186.855 ;
        RECT 23.740 -188.190 23.910 -186.730 ;
        RECT 26.450 -188.190 26.620 -186.710 ;
        RECT 27.430 -188.190 27.600 -186.710 ;
        RECT 28.410 -188.190 28.580 -186.710 ;
        RECT 29.110 -186.880 29.725 -186.710 ;
        RECT 35.190 -186.340 35.805 -186.205 ;
        RECT 35.190 -186.685 40.455 -186.340 ;
        RECT 29.390 -188.190 29.560 -186.880 ;
        RECT 35.190 -186.885 35.805 -186.685 ;
        RECT 35.195 -187.330 35.395 -186.885 ;
        RECT 36.140 -187.330 36.370 -186.685 ;
        RECT 37.130 -187.310 37.360 -186.685 ;
        RECT 35.195 -188.245 35.365 -187.330 ;
        RECT 36.175 -188.245 36.345 -187.330 ;
        RECT 37.155 -188.245 37.325 -187.310 ;
        RECT 37.695 -187.330 37.925 -186.685 ;
        RECT 38.675 -187.305 38.905 -186.685 ;
        RECT 37.725 -188.245 37.895 -187.330 ;
        RECT 38.705 -188.245 38.875 -187.305 ;
        RECT 39.240 -187.355 39.470 -186.685 ;
        RECT 40.225 -187.295 40.455 -186.685 ;
        RECT 39.270 -188.245 39.440 -187.355 ;
        RECT 40.250 -188.245 40.420 -187.295 ;
        RECT 101.355 -188.015 127.480 -187.700 ;
        RECT 106.115 -188.040 115.125 -188.015 ;
        RECT 119.615 -188.040 127.480 -188.015 ;
        RECT 138.280 -188.020 138.450 -186.690 ;
        RECT 139.260 -188.020 139.430 -186.690 ;
        RECT 140.240 -188.020 140.410 -186.690 ;
        RECT 141.220 -188.020 141.390 -186.690 ;
        RECT 106.420 -189.495 106.590 -188.040 ;
        RECT 107.400 -189.495 107.570 -188.040 ;
        RECT 108.380 -189.495 108.550 -188.040 ;
        RECT 110.605 -189.495 110.775 -188.040 ;
        RECT 111.585 -189.495 111.755 -188.040 ;
        RECT 112.565 -189.495 112.735 -188.040 ;
        RECT 119.920 -189.495 120.090 -188.040 ;
        RECT 120.900 -189.495 121.070 -188.040 ;
        RECT 121.880 -189.495 122.050 -188.040 ;
        RECT 124.105 -189.495 124.275 -188.040 ;
        RECT 125.085 -189.495 125.255 -188.040 ;
        RECT 126.065 -189.495 126.235 -188.040 ;
        RECT 127.035 -188.340 127.480 -188.040 ;
        RECT 138.040 -188.340 141.630 -188.020 ;
        RECT 127.035 -188.515 141.630 -188.340 ;
        RECT 127.035 -189.465 139.810 -188.515 ;
        RECT 143.145 -188.920 143.315 -186.835 ;
        RECT 144.125 -188.920 144.295 -186.835 ;
        RECT 145.105 -188.670 145.275 -186.835 ;
        RECT 146.190 -188.670 146.360 -187.840 ;
        RECT 147.170 -188.670 147.340 -187.840 ;
        RECT 148.150 -188.670 148.320 -187.840 ;
        RECT 149.130 -188.670 149.300 -187.840 ;
        RECT 180.480 -188.075 180.650 -186.745 ;
        RECT 181.460 -188.075 181.630 -186.745 ;
        RECT 182.440 -188.075 182.610 -186.745 ;
        RECT 183.420 -188.075 183.590 -186.745 ;
        RECT 180.240 -188.570 183.830 -188.075 ;
        RECT 145.105 -188.920 149.540 -188.670 ;
        RECT 143.095 -189.165 149.540 -188.920 ;
        RECT 143.095 -189.235 145.305 -189.165 ;
        RECT 155.330 -189.195 167.490 -188.845 ;
        RECT 143.090 -189.380 145.305 -189.235 ;
        RECT 143.090 -189.465 146.180 -189.380 ;
        RECT 153.495 -189.455 167.490 -189.195 ;
        RECT 153.495 -189.460 162.260 -189.455 ;
        RECT 127.035 -189.810 148.655 -189.465 ;
        RECT -32.835 -195.155 -32.665 -193.700 ;
        RECT -31.855 -195.155 -31.685 -193.700 ;
        RECT -30.875 -195.155 -30.705 -193.700 ;
        RECT -28.650 -195.155 -28.480 -193.700 ;
        RECT -27.670 -195.155 -27.500 -193.700 ;
        RECT -26.690 -195.155 -26.520 -193.700 ;
        RECT -19.335 -195.155 -19.165 -193.700 ;
        RECT -18.355 -195.155 -18.185 -193.700 ;
        RECT -17.375 -195.155 -17.205 -193.700 ;
        RECT -15.150 -195.155 -14.980 -193.700 ;
        RECT -14.170 -195.155 -14.000 -193.700 ;
        RECT -13.190 -195.155 -13.020 -193.700 ;
        RECT -34.080 -195.180 -26.215 -195.155 ;
        RECT -21.725 -195.180 -12.715 -195.155 ;
        RECT -34.080 -195.495 -7.955 -195.180 ;
        RECT 90.385 -195.445 90.555 -192.445 ;
        RECT 91.365 -195.365 91.535 -192.445 ;
        RECT -34.080 -198.690 -33.635 -195.495 ;
        RECT -53.060 -198.800 -33.635 -198.690 ;
        RECT -127.845 -199.715 -126.915 -199.635 ;
        RECT -130.080 -199.885 -126.915 -199.715 ;
        RECT -127.845 -199.930 -126.915 -199.885 ;
        RECT -127.845 -200.795 -127.605 -199.930 ;
        RECT -127.245 -200.795 -126.915 -199.930 ;
        RECT -127.845 -200.895 -126.915 -200.795 ;
        RECT -130.080 -201.065 -126.915 -200.895 ;
        RECT -127.845 -201.090 -126.915 -201.065 ;
        RECT -127.845 -202.000 -127.605 -201.090 ;
        RECT -127.245 -202.000 -126.915 -201.090 ;
        RECT -127.845 -202.075 -126.915 -202.000 ;
        RECT -130.080 -202.245 -126.915 -202.075 ;
        RECT -127.845 -202.295 -126.915 -202.245 ;
        RECT -73.450 -199.115 -33.635 -198.800 ;
        RECT -73.450 -199.140 -65.585 -199.115 ;
        RECT -61.095 -199.140 -52.085 -199.115 ;
        RECT -73.450 -202.265 -73.005 -199.140 ;
        RECT -72.205 -200.595 -72.035 -199.140 ;
        RECT -71.225 -200.595 -71.055 -199.140 ;
        RECT -70.245 -200.595 -70.075 -199.140 ;
        RECT -68.020 -200.595 -67.850 -199.140 ;
        RECT -67.040 -200.595 -66.870 -199.140 ;
        RECT -66.060 -200.595 -65.890 -199.140 ;
        RECT -58.705 -200.595 -58.535 -199.140 ;
        RECT -57.725 -200.595 -57.555 -199.140 ;
        RECT -56.745 -200.595 -56.575 -199.140 ;
        RECT -54.520 -200.595 -54.350 -199.140 ;
        RECT -53.540 -200.595 -53.370 -199.140 ;
        RECT -52.560 -200.595 -52.390 -199.140 ;
        RECT -40.280 -199.720 -40.055 -199.115 ;
        RECT -38.170 -199.715 -37.945 -199.115 ;
        RECT -127.845 -203.255 -127.605 -202.295 ;
        RECT -130.080 -203.355 -127.605 -203.255 ;
        RECT -127.245 -203.355 -126.915 -202.295 ;
        RECT -111.185 -203.100 -73.000 -202.265 ;
        RECT -40.260 -202.680 -40.090 -199.720 ;
        RECT -38.145 -202.680 -37.975 -199.715 ;
        RECT -37.195 -199.730 -36.970 -199.115 ;
        RECT -34.080 -199.690 -33.635 -199.115 ;
        RECT -37.165 -202.680 -36.995 -199.730 ;
        RECT -34.080 -200.135 -33.630 -199.690 ;
        RECT -32.640 -200.135 -31.295 -195.495 ;
        RECT -29.910 -200.135 -28.565 -195.495 ;
        RECT -25.525 -200.135 -24.180 -195.495 ;
        RECT -21.215 -200.135 -19.870 -195.495 ;
        RECT -16.700 -200.135 -15.355 -195.495 ;
        RECT -11.545 -200.135 -10.200 -195.495 ;
        RECT 90.340 -196.005 90.605 -195.445 ;
        RECT 91.320 -196.005 91.585 -195.365 ;
        RECT 90.340 -196.670 94.680 -196.005 ;
        RECT 96.990 -196.500 97.160 -195.045 ;
        RECT 97.970 -196.500 98.140 -195.045 ;
        RECT 98.950 -196.500 99.120 -195.045 ;
        RECT 101.400 -196.500 101.570 -195.045 ;
        RECT 102.380 -196.500 102.550 -195.045 ;
        RECT 103.360 -196.500 103.530 -195.045 ;
        RECT 110.115 -196.500 110.285 -195.045 ;
        RECT 111.095 -196.500 111.265 -195.045 ;
        RECT 112.075 -196.500 112.245 -195.045 ;
        RECT 114.900 -196.500 115.070 -195.045 ;
        RECT 115.880 -196.500 116.050 -195.045 ;
        RECT 116.860 -196.500 117.030 -195.045 ;
        RECT 123.615 -196.500 123.785 -195.045 ;
        RECT 124.595 -196.500 124.765 -195.045 ;
        RECT 125.575 -196.500 125.745 -195.045 ;
        RECT 96.945 -196.525 103.835 -196.500 ;
        RECT 110.070 -196.505 117.335 -196.500 ;
        RECT 108.505 -196.525 117.335 -196.505 ;
        RECT 123.570 -196.515 126.045 -196.500 ;
        RECT 127.035 -196.515 127.480 -189.810 ;
        RECT 138.100 -190.020 148.655 -189.810 ;
        RECT 153.495 -189.780 155.520 -189.460 ;
        RECT 150.680 -189.830 151.170 -189.815 ;
        RECT 153.495 -189.830 154.080 -189.780 ;
        RECT 138.100 -190.055 149.175 -190.020 ;
        RECT 149.540 -190.055 149.850 -189.915 ;
        RECT 138.100 -190.230 149.850 -190.055 ;
        RECT 140.110 -190.265 141.240 -190.230 ;
        RECT 140.295 -190.300 141.240 -190.265 ;
        RECT 145.330 -190.315 149.850 -190.230 ;
        RECT 145.330 -190.350 149.175 -190.315 ;
        RECT 138.100 -190.545 140.310 -190.470 ;
        RECT 138.100 -190.790 144.545 -190.545 ;
        RECT 138.150 -192.875 138.320 -190.790 ;
        RECT 139.130 -192.875 139.300 -190.790 ;
        RECT 140.110 -191.040 144.545 -190.790 ;
        RECT 145.360 -190.980 145.585 -190.350 ;
        RECT 146.335 -190.965 146.560 -190.350 ;
        RECT 140.110 -192.875 140.280 -191.040 ;
        RECT 141.195 -191.870 141.365 -191.040 ;
        RECT 142.175 -191.870 142.345 -191.040 ;
        RECT 143.155 -191.870 143.325 -191.040 ;
        RECT 144.135 -191.870 144.305 -191.040 ;
        RECT 145.385 -193.930 145.555 -190.980 ;
        RECT 146.365 -193.930 146.535 -190.965 ;
        RECT 148.445 -190.970 148.670 -190.350 ;
        RECT 149.540 -190.385 149.850 -190.315 ;
        RECT 150.680 -190.415 154.080 -189.830 ;
        RECT 155.330 -190.255 155.520 -189.780 ;
        RECT 156.315 -190.245 156.505 -189.460 ;
        RECT 150.680 -190.445 151.170 -190.415 ;
        RECT 148.480 -193.930 148.650 -190.970 ;
        RECT 155.345 -192.720 155.515 -190.255 ;
        RECT 156.325 -192.720 156.495 -190.245 ;
        RECT 159.275 -190.360 159.525 -189.460 ;
        RECT 159.905 -190.345 160.155 -189.460 ;
        RECT 161.060 -190.270 161.275 -189.460 ;
        RECT 162.045 -190.260 162.260 -189.460 ;
        RECT 166.880 -189.520 167.490 -189.455 ;
        RECT 181.150 -189.520 182.010 -188.570 ;
        RECT 185.345 -188.975 185.515 -186.890 ;
        RECT 186.325 -188.975 186.495 -186.890 ;
        RECT 187.305 -188.725 187.475 -186.890 ;
        RECT 188.390 -188.725 188.560 -187.895 ;
        RECT 189.370 -188.725 189.540 -187.895 ;
        RECT 190.350 -188.725 190.520 -187.895 ;
        RECT 191.330 -188.725 191.500 -187.895 ;
        RECT 224.795 -188.270 224.965 -186.940 ;
        RECT 225.775 -188.270 225.945 -186.940 ;
        RECT 226.755 -188.270 226.925 -186.940 ;
        RECT 227.735 -188.270 227.905 -186.940 ;
        RECT 224.555 -188.690 228.145 -188.270 ;
        RECT 187.305 -188.975 191.740 -188.725 ;
        RECT 204.390 -188.765 228.145 -188.690 ;
        RECT 204.390 -188.900 226.325 -188.765 ;
        RECT 185.295 -189.220 191.740 -188.975 ;
        RECT 185.295 -189.290 187.505 -189.220 ;
        RECT 197.530 -189.250 226.325 -188.900 ;
        RECT 229.660 -189.170 229.830 -187.085 ;
        RECT 230.640 -189.170 230.810 -187.085 ;
        RECT 231.620 -188.920 231.790 -187.085 ;
        RECT 232.705 -188.920 232.875 -188.090 ;
        RECT 233.685 -188.920 233.855 -188.090 ;
        RECT 234.665 -188.920 234.835 -188.090 ;
        RECT 235.645 -188.920 235.815 -188.090 ;
        RECT 270.785 -188.100 270.955 -186.770 ;
        RECT 271.765 -188.100 271.935 -186.770 ;
        RECT 272.745 -188.100 272.915 -186.770 ;
        RECT 273.725 -188.100 273.895 -186.770 ;
        RECT 270.545 -188.440 274.135 -188.100 ;
        RECT 248.645 -188.595 274.135 -188.440 ;
        RECT 231.620 -189.170 236.055 -188.920 ;
        RECT 248.645 -189.095 272.315 -188.595 ;
        RECT 275.650 -189.000 275.820 -186.915 ;
        RECT 276.630 -189.000 276.800 -186.915 ;
        RECT 277.610 -188.750 277.780 -186.915 ;
        RECT 314.555 -187.770 314.725 -186.440 ;
        RECT 315.535 -187.770 315.705 -186.440 ;
        RECT 316.515 -187.770 316.685 -186.440 ;
        RECT 317.495 -187.770 317.665 -186.440 ;
        RECT 278.695 -188.750 278.865 -187.920 ;
        RECT 279.675 -188.750 279.845 -187.920 ;
        RECT 280.655 -188.750 280.825 -187.920 ;
        RECT 281.635 -188.750 281.805 -187.920 ;
        RECT 314.315 -187.955 317.905 -187.770 ;
        RECT 294.560 -188.265 317.905 -187.955 ;
        RECT 277.610 -189.000 282.045 -188.750 ;
        RECT 294.560 -188.925 316.085 -188.265 ;
        RECT 319.420 -188.670 319.590 -186.585 ;
        RECT 320.400 -188.670 320.570 -186.585 ;
        RECT 321.380 -188.420 321.550 -186.585 ;
        RECT 322.465 -188.420 322.635 -187.590 ;
        RECT 323.445 -188.420 323.615 -187.590 ;
        RECT 324.425 -188.420 324.595 -187.590 ;
        RECT 325.405 -188.420 325.575 -187.590 ;
        RECT 360.320 -187.685 360.490 -186.355 ;
        RECT 361.300 -187.685 361.470 -186.355 ;
        RECT 362.280 -187.685 362.450 -186.355 ;
        RECT 363.260 -187.685 363.430 -186.355 ;
        RECT 360.080 -188.060 363.670 -187.685 ;
        RECT 338.295 -188.180 363.670 -188.060 ;
        RECT 321.380 -188.670 325.815 -188.420 ;
        RECT 338.295 -188.595 361.850 -188.180 ;
        RECT 365.185 -188.585 365.355 -186.500 ;
        RECT 366.165 -188.585 366.335 -186.500 ;
        RECT 367.145 -188.335 367.315 -186.500 ;
        RECT 407.140 -187.495 407.310 -186.165 ;
        RECT 408.120 -187.495 408.290 -186.165 ;
        RECT 409.100 -187.495 409.270 -186.165 ;
        RECT 410.080 -187.495 410.250 -186.165 ;
        RECT 368.230 -188.335 368.400 -187.505 ;
        RECT 369.210 -188.335 369.380 -187.505 ;
        RECT 370.190 -188.335 370.360 -187.505 ;
        RECT 371.170 -188.335 371.340 -187.505 ;
        RECT 406.900 -187.715 410.490 -187.495 ;
        RECT 384.105 -187.990 410.490 -187.715 ;
        RECT 367.145 -188.585 371.580 -188.335 ;
        RECT 384.105 -188.510 408.670 -187.990 ;
        RECT 412.005 -188.395 412.175 -186.310 ;
        RECT 412.985 -188.395 413.155 -186.310 ;
        RECT 413.965 -188.145 414.135 -186.310 ;
        RECT 415.050 -188.145 415.220 -187.315 ;
        RECT 416.030 -188.145 416.200 -187.315 ;
        RECT 417.010 -188.145 417.180 -187.315 ;
        RECT 417.990 -188.145 418.160 -187.315 ;
        RECT 413.965 -188.395 418.400 -188.145 ;
        RECT 432.980 -188.320 435.355 -168.760 ;
        RECT 185.290 -189.435 187.505 -189.290 ;
        RECT 185.290 -189.520 188.380 -189.435 ;
        RECT 195.695 -189.515 226.325 -189.250 ;
        RECT 229.610 -189.415 236.055 -189.170 ;
        RECT 229.610 -189.485 231.820 -189.415 ;
        RECT 241.845 -189.445 272.315 -189.095 ;
        RECT 275.600 -189.245 282.045 -189.000 ;
        RECT 287.835 -189.215 316.085 -188.925 ;
        RECT 319.370 -188.915 325.815 -188.670 ;
        RECT 319.370 -188.985 321.580 -188.915 ;
        RECT 331.605 -188.945 361.850 -188.595 ;
        RECT 365.135 -188.830 371.580 -188.585 ;
        RECT 365.135 -188.900 367.345 -188.830 ;
        RECT 377.370 -188.860 408.670 -188.510 ;
        RECT 411.955 -188.640 418.400 -188.395 ;
        RECT 411.955 -188.710 414.165 -188.640 ;
        RECT 424.190 -188.670 436.350 -188.320 ;
        RECT 319.365 -189.130 321.580 -188.985 ;
        RECT 329.770 -189.130 361.850 -188.945 ;
        RECT 365.130 -189.045 367.345 -188.900 ;
        RECT 375.535 -188.940 408.670 -188.860 ;
        RECT 411.950 -188.855 414.165 -188.710 ;
        RECT 411.950 -188.940 415.040 -188.855 ;
        RECT 422.355 -188.930 436.350 -188.670 ;
        RECT 422.355 -188.935 431.120 -188.930 ;
        RECT 365.130 -189.130 368.220 -189.045 ;
        RECT 375.535 -189.125 417.515 -188.940 ;
        RECT 319.365 -189.215 322.455 -189.130 ;
        RECT 329.770 -189.210 370.695 -189.130 ;
        RECT 275.600 -189.315 277.810 -189.245 ;
        RECT 287.835 -189.275 324.930 -189.215 ;
        RECT 166.880 -190.075 190.855 -189.520 ;
        RECT 195.695 -189.835 197.720 -189.515 ;
        RECT 192.880 -189.885 193.370 -189.870 ;
        RECT 195.695 -189.885 196.280 -189.835 ;
        RECT 166.880 -190.110 191.375 -190.075 ;
        RECT 191.740 -190.110 192.050 -189.970 ;
        RECT 159.300 -192.720 159.470 -190.360 ;
        RECT 159.950 -192.720 160.120 -190.345 ;
        RECT 161.090 -191.720 161.260 -190.270 ;
        RECT 162.070 -191.720 162.240 -190.260 ;
        RECT 166.880 -190.285 192.050 -190.110 ;
        RECT 121.960 -196.525 127.480 -196.515 ;
        RECT 96.945 -196.840 127.480 -196.525 ;
        RECT 108.505 -196.845 110.870 -196.840 ;
        RECT 109.455 -197.940 110.615 -196.845 ;
        RECT 121.960 -196.855 127.480 -196.840 ;
        RECT 109.165 -198.260 111.375 -197.940 ;
        RECT -34.080 -200.450 -7.955 -200.135 ;
        RECT -34.080 -200.475 -26.215 -200.450 ;
        RECT -21.725 -200.475 -12.715 -200.450 ;
        RECT -130.080 -203.425 -126.915 -203.355 ;
        RECT -127.845 -203.650 -126.915 -203.425 ;
        RECT -127.845 -204.435 -127.605 -203.650 ;
        RECT -130.080 -204.605 -127.605 -204.435 ;
        RECT -127.845 -205.085 -127.605 -204.605 ;
        RECT -130.080 -205.255 -127.605 -205.085 ;
        RECT -127.845 -206.265 -127.605 -205.255 ;
        RECT -130.080 -206.295 -127.605 -206.265 ;
        RECT -127.245 -206.295 -126.915 -203.650 ;
        RECT -109.335 -203.795 -105.425 -203.100 ;
        RECT -103.545 -203.730 -100.955 -203.100 ;
        RECT -109.635 -204.460 -105.295 -203.795 ;
        RECT -103.620 -204.075 -100.850 -203.730 ;
        RECT -99.100 -203.735 -96.335 -203.100 ;
        RECT -99.100 -203.940 -96.325 -203.735 ;
        RECT -109.635 -205.020 -109.370 -204.460 ;
        RECT -130.080 -206.435 -126.915 -206.295 ;
        RECT -127.845 -206.590 -126.915 -206.435 ;
        RECT -127.845 -207.445 -127.605 -206.590 ;
        RECT -130.080 -207.615 -127.605 -207.445 ;
        RECT -127.245 -207.595 -126.915 -206.590 ;
        RECT -109.590 -208.020 -109.420 -205.020 ;
        RECT -108.655 -205.100 -108.390 -204.460 ;
        RECT -103.595 -204.710 -103.355 -204.075 ;
        RECT -108.610 -208.020 -108.440 -205.100 ;
        RECT -103.560 -206.665 -103.390 -204.710 ;
        RECT -102.610 -204.740 -102.370 -204.075 ;
        RECT -99.095 -204.080 -96.325 -203.940 ;
        RECT -99.070 -204.715 -98.830 -204.080 ;
        RECT -102.580 -206.665 -102.410 -204.740 ;
        RECT -99.035 -206.670 -98.865 -204.715 ;
        RECT -98.085 -204.745 -97.845 -204.080 ;
        RECT -98.055 -206.670 -97.885 -204.745 ;
        RECT -73.450 -207.615 -73.005 -203.100 ;
        RECT -71.715 -207.600 -71.545 -206.145 ;
        RECT -70.735 -207.600 -70.565 -206.145 ;
        RECT -69.755 -207.600 -69.585 -206.145 ;
        RECT -63.000 -207.600 -62.830 -206.145 ;
        RECT -62.020 -207.600 -61.850 -206.145 ;
        RECT -61.040 -207.600 -60.870 -206.145 ;
        RECT -58.215 -207.600 -58.045 -206.145 ;
        RECT -57.235 -207.600 -57.065 -206.145 ;
        RECT -56.255 -207.600 -56.085 -206.145 ;
        RECT -49.500 -207.600 -49.330 -206.145 ;
        RECT -48.520 -207.600 -48.350 -206.145 ;
        RECT -47.540 -207.600 -47.370 -206.145 ;
        RECT -45.090 -207.600 -44.920 -206.145 ;
        RECT -44.110 -207.600 -43.940 -206.145 ;
        RECT -43.130 -207.600 -42.960 -206.145 ;
        RECT -72.015 -207.615 -69.540 -207.600 ;
        RECT -63.305 -207.605 -56.040 -207.600 ;
        RECT -73.450 -207.625 -67.930 -207.615 ;
        RECT -63.305 -207.625 -54.475 -207.605 ;
        RECT -49.805 -207.625 -42.915 -207.600 ;
        RECT -73.450 -207.940 -42.915 -207.625 ;
        RECT -73.450 -207.955 -67.930 -207.940 ;
        RECT -56.840 -207.945 -54.475 -207.940 ;
        RECT -92.025 -211.360 -91.855 -209.275 ;
        RECT -91.045 -211.360 -90.875 -209.275 ;
        RECT -90.065 -211.110 -89.895 -209.275 ;
        RECT -88.980 -211.110 -88.810 -210.280 ;
        RECT -88.000 -211.110 -87.830 -210.280 ;
        RECT -87.020 -211.110 -86.850 -210.280 ;
        RECT -86.040 -211.110 -85.870 -210.280 ;
        RECT -90.065 -211.360 -85.630 -211.110 ;
        RECT -84.790 -211.170 -84.620 -208.220 ;
        RECT -92.075 -211.605 -85.630 -211.360 ;
        RECT -92.075 -211.680 -89.865 -211.605 ;
        RECT -84.815 -211.800 -84.590 -211.170 ;
        RECT -83.810 -211.185 -83.640 -208.220 ;
        RECT -81.695 -211.180 -81.525 -208.220 ;
        RECT -34.080 -208.950 -33.635 -200.475 ;
        RECT -32.835 -201.930 -32.665 -200.475 ;
        RECT -31.855 -201.930 -31.685 -200.475 ;
        RECT -30.875 -201.930 -30.705 -200.475 ;
        RECT -28.650 -201.930 -28.480 -200.475 ;
        RECT -27.670 -201.930 -27.500 -200.475 ;
        RECT -26.690 -201.930 -26.520 -200.475 ;
        RECT -19.335 -201.930 -19.165 -200.475 ;
        RECT -18.355 -201.930 -18.185 -200.475 ;
        RECT -17.375 -201.930 -17.205 -200.475 ;
        RECT -15.150 -201.930 -14.980 -200.475 ;
        RECT -14.170 -201.930 -14.000 -200.475 ;
        RECT -13.190 -201.930 -13.020 -200.475 ;
        RECT 109.215 -200.845 109.385 -198.260 ;
        RECT 110.195 -200.845 110.365 -198.260 ;
        RECT 111.175 -200.845 111.345 -198.260 ;
        RECT -32.345 -208.935 -32.175 -207.480 ;
        RECT -31.365 -208.935 -31.195 -207.480 ;
        RECT -30.385 -208.935 -30.215 -207.480 ;
        RECT -23.630 -208.935 -23.460 -207.480 ;
        RECT -22.650 -208.935 -22.480 -207.480 ;
        RECT -21.670 -208.935 -21.500 -207.480 ;
        RECT -18.845 -208.935 -18.675 -207.480 ;
        RECT -17.865 -208.935 -17.695 -207.480 ;
        RECT -16.885 -208.935 -16.715 -207.480 ;
        RECT -10.130 -208.935 -9.960 -207.480 ;
        RECT -9.150 -208.935 -8.980 -207.480 ;
        RECT -8.170 -208.935 -8.000 -207.480 ;
        RECT -5.720 -208.935 -5.550 -207.480 ;
        RECT -4.740 -208.935 -4.570 -207.480 ;
        RECT -3.760 -208.705 -3.590 -207.480 ;
        RECT -4.120 -208.935 -3.505 -208.705 ;
        RECT -2.050 -208.710 -1.880 -207.395 ;
        RECT -32.645 -208.950 -30.170 -208.935 ;
        RECT -23.935 -208.940 -16.670 -208.935 ;
        RECT -34.080 -208.960 -28.560 -208.950 ;
        RECT -23.935 -208.960 -15.105 -208.940 ;
        RECT -10.435 -208.960 -3.505 -208.935 ;
        RECT -34.080 -209.275 -3.505 -208.960 ;
        RECT -34.080 -209.290 -28.560 -209.275 ;
        RECT -83.840 -211.800 -83.615 -211.185 ;
        RECT -81.730 -211.800 -81.505 -211.180 ;
        RECT -89.880 -211.885 -88.935 -211.850 ;
        RECT -90.065 -211.920 -88.935 -211.885 ;
        RECT -84.845 -211.920 -81.000 -211.800 ;
        RECT -98.245 -212.130 -81.000 -211.920 ;
        RECT -23.225 -212.035 -22.650 -209.275 ;
        RECT -17.470 -209.280 -15.105 -209.275 ;
        RECT -98.245 -212.685 -81.520 -212.130 ;
        RECT -98.245 -212.780 -90.365 -212.685 ;
        RECT -98.245 -217.755 -97.385 -212.780 ;
        RECT -91.225 -213.635 -90.365 -212.780 ;
        RECT -87.085 -212.770 -83.995 -212.685 ;
        RECT -23.250 -212.715 -22.635 -212.035 ;
        RECT -10.395 -212.755 -9.820 -209.275 ;
        RECT -4.120 -209.385 -3.505 -209.275 ;
        RECT -2.650 -208.855 -1.880 -208.710 ;
        RECT -1.070 -208.855 -0.900 -207.395 ;
        RECT -2.650 -208.860 -0.875 -208.855 ;
        RECT 1.640 -208.860 1.810 -207.395 ;
        RECT 2.620 -208.860 2.790 -207.395 ;
        RECT 3.600 -208.860 3.770 -207.395 ;
        RECT 4.580 -208.860 4.750 -207.395 ;
        RECT 6.615 -208.660 6.785 -207.830 ;
        RECT 7.595 -208.660 7.765 -207.830 ;
        RECT 8.575 -208.660 8.745 -207.830 ;
        RECT 9.555 -208.660 9.725 -207.830 ;
        RECT 10.640 -208.660 10.810 -206.825 ;
        RECT 6.375 -208.860 10.810 -208.660 ;
        RECT 11.620 -208.860 11.790 -206.825 ;
        RECT 12.600 -208.645 12.770 -206.825 ;
        RECT 12.240 -208.860 12.855 -208.645 ;
        RECT 14.640 -208.650 14.810 -207.820 ;
        RECT 15.620 -208.650 15.790 -207.820 ;
        RECT 16.600 -208.650 16.770 -207.820 ;
        RECT 17.580 -208.650 17.750 -207.820 ;
        RECT 18.665 -208.650 18.835 -206.815 ;
        RECT -2.650 -209.255 12.855 -208.860 ;
        RECT -2.650 -209.390 -2.035 -209.255 ;
        RECT -87.085 -212.915 -84.870 -212.770 ;
        RECT -87.080 -212.985 -84.870 -212.915 ;
        RECT -87.080 -213.230 -80.635 -212.985 ;
        RECT -92.135 -214.130 -88.545 -213.635 ;
        RECT -91.895 -215.460 -91.725 -214.130 ;
        RECT -90.915 -215.460 -90.745 -214.130 ;
        RECT -89.935 -215.460 -89.765 -214.130 ;
        RECT -88.955 -215.460 -88.785 -214.130 ;
        RECT -87.030 -215.315 -86.860 -213.230 ;
        RECT -86.050 -215.315 -85.880 -213.230 ;
        RECT -85.070 -213.480 -80.635 -213.230 ;
        RECT -10.415 -213.435 -9.800 -212.755 ;
        RECT 2.025 -213.295 2.600 -209.255 ;
        RECT 12.240 -209.325 12.855 -209.255 ;
        RECT 14.185 -208.900 18.835 -208.650 ;
        RECT 19.645 -208.900 19.815 -206.815 ;
        RECT 20.625 -208.765 20.795 -206.815 ;
        RECT 90.360 -207.130 90.530 -205.175 ;
        RECT 91.340 -207.100 91.510 -205.175 ;
        RECT 20.325 -208.900 20.940 -208.765 ;
        RECT 22.760 -208.775 22.930 -207.440 ;
        RECT 14.185 -209.145 20.940 -208.900 ;
        RECT 14.185 -209.330 14.800 -209.145 ;
        RECT 18.635 -209.220 20.940 -209.145 ;
        RECT 20.325 -209.445 20.940 -209.220 ;
        RECT 22.330 -208.900 22.945 -208.775 ;
        RECT 23.740 -208.900 23.910 -207.440 ;
        RECT 22.330 -208.925 23.935 -208.900 ;
        RECT 26.450 -208.920 26.620 -207.440 ;
        RECT 27.430 -208.920 27.600 -207.440 ;
        RECT 28.410 -208.920 28.580 -207.440 ;
        RECT 29.390 -208.750 29.560 -207.440 ;
        RECT 35.195 -208.300 35.365 -207.385 ;
        RECT 36.175 -208.300 36.345 -207.385 ;
        RECT 35.195 -208.745 35.395 -208.300 ;
        RECT 29.110 -208.920 29.725 -208.750 ;
        RECT 26.450 -208.925 29.725 -208.920 ;
        RECT 22.330 -209.265 29.725 -208.925 ;
        RECT 22.330 -209.290 26.810 -209.265 ;
        RECT 22.330 -209.455 22.945 -209.290 ;
        RECT 29.110 -209.430 29.725 -209.265 ;
        RECT 35.190 -208.945 35.805 -208.745 ;
        RECT 36.140 -208.945 36.370 -208.300 ;
        RECT 37.155 -208.320 37.325 -207.385 ;
        RECT 37.725 -208.300 37.895 -207.385 ;
        RECT 37.130 -208.945 37.360 -208.320 ;
        RECT 37.695 -208.945 37.925 -208.300 ;
        RECT 38.705 -208.325 38.875 -207.385 ;
        RECT 39.270 -208.275 39.440 -207.385 ;
        RECT 38.675 -208.945 38.905 -208.325 ;
        RECT 39.240 -208.945 39.470 -208.275 ;
        RECT 40.250 -208.335 40.420 -207.385 ;
        RECT 90.325 -207.765 90.565 -207.130 ;
        RECT 91.310 -207.765 91.550 -207.100 ;
        RECT 95.090 -207.130 95.260 -205.175 ;
        RECT 96.070 -207.100 96.240 -205.175 ;
        RECT 95.055 -207.765 95.295 -207.130 ;
        RECT 96.040 -207.765 96.280 -207.100 ;
        RECT 98.445 -207.765 98.875 -207.725 ;
        RECT 86.210 -207.825 98.875 -207.765 ;
        RECT 99.670 -207.825 99.840 -206.345 ;
        RECT 100.650 -207.825 100.820 -206.345 ;
        RECT 101.630 -207.825 101.800 -206.345 ;
        RECT 102.610 -207.825 102.780 -206.345 ;
        RECT 104.045 -207.805 104.360 -207.735 ;
        RECT 105.320 -207.805 105.490 -206.345 ;
        RECT 106.300 -207.805 106.470 -206.345 ;
        RECT 107.450 -207.765 107.820 -207.735 ;
        RECT 108.965 -207.765 109.135 -206.310 ;
        RECT 109.945 -207.765 110.115 -206.310 ;
        RECT 110.925 -207.630 111.095 -206.310 ;
        RECT 113.365 -207.630 113.535 -203.455 ;
        RECT 114.345 -207.630 114.515 -203.455 ;
        RECT 115.365 -207.630 115.535 -203.455 ;
        RECT 116.345 -207.630 116.515 -203.455 ;
        RECT 118.365 -207.630 118.535 -203.455 ;
        RECT 119.345 -207.630 119.515 -203.455 ;
        RECT 120.365 -207.630 120.535 -203.455 ;
        RECT 121.345 -207.630 121.515 -203.455 ;
        RECT 123.365 -207.630 123.535 -203.455 ;
        RECT 124.345 -207.630 124.515 -203.455 ;
        RECT 125.365 -207.630 125.535 -203.455 ;
        RECT 126.345 -207.630 126.515 -203.455 ;
        RECT 127.035 -207.630 127.480 -196.855 ;
        RECT 150.715 -200.405 152.725 -200.075 ;
        RECT 138.240 -205.285 138.410 -203.955 ;
        RECT 139.220 -205.285 139.390 -203.955 ;
        RECT 140.200 -205.285 140.370 -203.955 ;
        RECT 141.180 -205.285 141.350 -203.955 ;
        RECT 138.000 -205.780 141.590 -205.285 ;
        RECT 138.910 -206.730 139.770 -205.780 ;
        RECT 143.105 -206.185 143.275 -204.100 ;
        RECT 144.085 -206.185 144.255 -204.100 ;
        RECT 145.065 -205.935 145.235 -204.100 ;
        RECT 146.150 -205.935 146.320 -205.105 ;
        RECT 147.130 -205.935 147.300 -205.105 ;
        RECT 148.110 -205.935 148.280 -205.105 ;
        RECT 149.090 -205.935 149.260 -205.105 ;
        RECT 145.065 -206.185 149.500 -205.935 ;
        RECT 143.055 -206.430 149.500 -206.185 ;
        RECT 143.055 -206.500 145.265 -206.430 ;
        RECT 143.050 -206.645 145.265 -206.500 ;
        RECT 143.050 -206.730 146.140 -206.645 ;
        RECT 138.060 -207.285 148.615 -206.730 ;
        RECT 150.715 -206.910 151.045 -200.405 ;
        RECT 138.060 -207.495 149.135 -207.285 ;
        RECT 150.630 -207.475 151.050 -206.910 ;
        RECT 152.395 -207.055 152.725 -200.405 ;
        RECT 166.880 -201.440 167.490 -190.285 ;
        RECT 182.310 -190.320 183.440 -190.285 ;
        RECT 182.495 -190.355 183.440 -190.320 ;
        RECT 187.530 -190.370 192.050 -190.285 ;
        RECT 187.530 -190.405 191.375 -190.370 ;
        RECT 180.300 -190.600 182.510 -190.525 ;
        RECT 180.300 -190.845 186.745 -190.600 ;
        RECT 180.350 -192.930 180.520 -190.845 ;
        RECT 181.330 -192.930 181.500 -190.845 ;
        RECT 182.310 -191.095 186.745 -190.845 ;
        RECT 187.560 -191.035 187.785 -190.405 ;
        RECT 188.535 -191.020 188.760 -190.405 ;
        RECT 182.310 -192.930 182.480 -191.095 ;
        RECT 183.395 -191.925 183.565 -191.095 ;
        RECT 184.375 -191.925 184.545 -191.095 ;
        RECT 185.355 -191.925 185.525 -191.095 ;
        RECT 186.335 -191.925 186.505 -191.095 ;
        RECT 187.585 -193.985 187.755 -191.035 ;
        RECT 188.565 -193.985 188.735 -191.020 ;
        RECT 190.645 -191.025 190.870 -190.405 ;
        RECT 191.740 -190.440 192.050 -190.370 ;
        RECT 192.880 -190.470 196.280 -189.885 ;
        RECT 197.530 -190.310 197.720 -189.835 ;
        RECT 198.515 -190.300 198.705 -189.515 ;
        RECT 192.880 -190.500 193.370 -190.470 ;
        RECT 190.680 -193.985 190.850 -191.025 ;
        RECT 197.545 -192.775 197.715 -190.310 ;
        RECT 198.525 -192.775 198.695 -190.300 ;
        RECT 201.475 -190.415 201.725 -189.515 ;
        RECT 202.105 -190.400 202.355 -189.515 ;
        RECT 203.260 -190.325 203.475 -189.515 ;
        RECT 204.245 -189.715 226.325 -189.515 ;
        RECT 229.605 -189.630 231.820 -189.485 ;
        RECT 240.010 -189.545 272.315 -189.445 ;
        RECT 275.595 -189.460 277.810 -189.315 ;
        RECT 275.595 -189.545 278.685 -189.460 ;
        RECT 286.000 -189.540 324.930 -189.275 ;
        RECT 229.605 -189.715 232.695 -189.630 ;
        RECT 240.010 -189.710 281.160 -189.545 ;
        RECT 204.245 -189.960 235.170 -189.715 ;
        RECT 204.245 -190.315 204.460 -189.960 ;
        RECT 201.500 -192.775 201.670 -190.415 ;
        RECT 202.150 -192.775 202.320 -190.400 ;
        RECT 203.290 -191.775 203.460 -190.325 ;
        RECT 204.270 -191.775 204.440 -190.315 ;
        RECT 192.915 -200.460 194.925 -200.130 ;
        RECT 166.880 -202.050 170.040 -201.440 ;
        RECT 156.580 -205.440 156.750 -204.110 ;
        RECT 157.560 -205.440 157.730 -204.110 ;
        RECT 158.540 -205.440 158.710 -204.110 ;
        RECT 159.520 -205.440 159.690 -204.110 ;
        RECT 156.340 -205.935 159.930 -205.440 ;
        RECT 157.250 -206.885 158.110 -205.935 ;
        RECT 161.445 -206.340 161.615 -204.255 ;
        RECT 162.425 -206.340 162.595 -204.255 ;
        RECT 163.405 -206.090 163.575 -204.255 ;
        RECT 164.490 -206.090 164.660 -205.260 ;
        RECT 165.470 -206.090 165.640 -205.260 ;
        RECT 166.450 -206.090 166.620 -205.260 ;
        RECT 167.430 -206.090 167.600 -205.260 ;
        RECT 163.405 -206.340 167.840 -206.090 ;
        RECT 161.395 -206.585 167.840 -206.340 ;
        RECT 161.395 -206.655 163.605 -206.585 ;
        RECT 161.390 -206.800 163.605 -206.655 ;
        RECT 161.390 -206.885 164.480 -206.800 ;
        RECT 156.400 -207.055 166.955 -206.885 ;
        RECT 169.430 -207.030 170.040 -202.050 ;
        RECT 180.440 -205.340 180.610 -204.010 ;
        RECT 181.420 -205.340 181.590 -204.010 ;
        RECT 182.400 -205.340 182.570 -204.010 ;
        RECT 183.380 -205.340 183.550 -204.010 ;
        RECT 180.200 -205.835 183.790 -205.340 ;
        RECT 181.110 -206.785 181.970 -205.835 ;
        RECT 185.305 -206.240 185.475 -204.155 ;
        RECT 186.285 -206.240 186.455 -204.155 ;
        RECT 187.265 -205.990 187.435 -204.155 ;
        RECT 188.350 -205.990 188.520 -205.160 ;
        RECT 189.330 -205.990 189.500 -205.160 ;
        RECT 190.310 -205.990 190.480 -205.160 ;
        RECT 191.290 -205.990 191.460 -205.160 ;
        RECT 187.265 -206.240 191.700 -205.990 ;
        RECT 185.255 -206.485 191.700 -206.240 ;
        RECT 185.255 -206.555 187.465 -206.485 ;
        RECT 185.250 -206.700 187.465 -206.555 ;
        RECT 185.250 -206.785 188.340 -206.700 ;
        RECT 152.395 -207.385 166.955 -207.055 ;
        RECT 167.730 -207.260 168.125 -207.105 ;
        RECT 156.400 -207.440 166.955 -207.385 ;
        RECT 167.230 -207.440 168.125 -207.260 ;
        RECT 140.070 -207.530 141.200 -207.495 ;
        RECT 140.255 -207.565 141.200 -207.530 ;
        RECT 145.290 -207.615 149.135 -207.495 ;
        RECT 110.925 -207.765 127.480 -207.630 ;
        RECT 107.450 -207.805 127.480 -207.765 ;
        RECT 104.045 -207.825 127.480 -207.805 ;
        RECT 86.210 -208.105 127.480 -207.825 ;
        RECT 138.060 -207.810 140.270 -207.735 ;
        RECT 138.060 -208.055 144.505 -207.810 ;
        RECT 86.210 -208.110 107.820 -208.105 ;
        RECT 40.225 -208.945 40.455 -208.335 ;
        RECT 35.190 -209.290 40.455 -208.945 ;
        RECT 35.190 -209.425 35.805 -209.290 ;
        RECT 86.210 -210.465 86.840 -208.110 ;
        RECT 98.445 -208.140 107.820 -208.110 ;
        RECT 98.445 -208.170 104.360 -208.140 ;
        RECT 107.450 -208.170 107.820 -208.140 ;
        RECT 111.035 -208.145 127.480 -208.105 ;
        RECT 98.445 -208.190 98.875 -208.170 ;
        RECT 104.045 -208.225 104.360 -208.170 ;
        RECT 138.110 -210.140 138.280 -208.055 ;
        RECT 139.090 -210.140 139.260 -208.055 ;
        RECT 140.070 -208.305 144.505 -208.055 ;
        RECT 145.320 -208.245 145.545 -207.615 ;
        RECT 146.295 -208.230 146.520 -207.615 ;
        RECT 140.070 -210.140 140.240 -208.305 ;
        RECT 141.155 -209.135 141.325 -208.305 ;
        RECT 142.135 -209.135 142.305 -208.305 ;
        RECT 143.115 -209.135 143.285 -208.305 ;
        RECT 144.095 -209.135 144.265 -208.305 ;
        RECT 67.865 -210.480 70.230 -210.475 ;
        RECT 81.320 -210.480 86.840 -210.465 ;
        RECT 56.305 -210.795 86.840 -210.480 ;
        RECT 56.305 -210.820 63.195 -210.795 ;
        RECT 67.865 -210.815 76.695 -210.795 ;
        RECT 81.320 -210.805 86.840 -210.795 ;
        RECT 69.430 -210.820 76.695 -210.815 ;
        RECT 82.930 -210.820 85.405 -210.805 ;
        RECT 56.350 -212.275 56.520 -210.820 ;
        RECT 57.330 -212.275 57.500 -210.820 ;
        RECT 58.310 -212.275 58.480 -210.820 ;
        RECT 60.760 -212.275 60.930 -210.820 ;
        RECT 61.740 -212.275 61.910 -210.820 ;
        RECT 62.720 -212.275 62.890 -210.820 ;
        RECT 69.475 -212.275 69.645 -210.820 ;
        RECT 70.455 -212.275 70.625 -210.820 ;
        RECT 71.435 -212.275 71.605 -210.820 ;
        RECT 74.260 -212.275 74.430 -210.820 ;
        RECT 75.240 -212.275 75.410 -210.820 ;
        RECT 76.220 -212.275 76.390 -210.820 ;
        RECT 82.975 -212.275 83.145 -210.820 ;
        RECT 83.955 -212.275 84.125 -210.820 ;
        RECT 84.935 -212.275 85.105 -210.820 ;
        RECT -85.070 -215.315 -84.900 -213.480 ;
        RECT -83.985 -214.310 -83.815 -213.480 ;
        RECT -83.005 -214.310 -82.835 -213.480 ;
        RECT -82.025 -214.310 -81.855 -213.480 ;
        RECT -81.045 -214.310 -80.875 -213.480 ;
        RECT 2.000 -213.605 3.530 -213.295 ;
        RECT 2.000 -213.610 2.615 -213.605 ;
        RECT -23.245 -216.550 -22.630 -215.870 ;
        RECT -10.410 -216.375 -9.795 -215.695 ;
        RECT 2.005 -216.375 2.620 -215.695 ;
        RECT -98.255 -218.190 -97.375 -217.755 ;
        RECT -111.275 -220.530 -111.105 -219.070 ;
        RECT -110.295 -220.450 -110.125 -219.070 ;
        RECT -107.585 -220.450 -107.415 -219.070 ;
        RECT -106.605 -220.450 -106.435 -219.070 ;
        RECT -105.625 -220.450 -105.455 -219.070 ;
        RECT -104.645 -220.450 -104.475 -219.070 ;
        RECT -29.855 -219.555 -29.685 -218.640 ;
        RECT -28.875 -219.555 -28.705 -218.640 ;
        RECT -29.855 -220.200 -29.655 -219.555 ;
        RECT -28.910 -220.200 -28.680 -219.555 ;
        RECT -27.895 -219.575 -27.725 -218.640 ;
        RECT -27.325 -219.555 -27.155 -218.640 ;
        RECT -27.920 -220.200 -27.690 -219.575 ;
        RECT -27.355 -220.200 -27.125 -219.555 ;
        RECT -26.345 -219.580 -26.175 -218.640 ;
        RECT -25.780 -219.530 -25.610 -218.640 ;
        RECT -26.375 -220.200 -26.145 -219.580 ;
        RECT -25.810 -220.200 -25.580 -219.530 ;
        RECT -24.800 -219.590 -24.630 -218.640 ;
        RECT -24.825 -220.200 -24.595 -219.590 ;
        RECT -110.385 -220.530 -97.375 -220.450 ;
        RECT -111.325 -220.865 -97.375 -220.530 ;
        RECT -29.855 -220.735 -24.595 -220.200 ;
        RECT -23.220 -220.735 -22.645 -216.550 ;
        RECT -17.355 -219.555 -17.185 -218.640 ;
        RECT -16.375 -219.555 -16.205 -218.640 ;
        RECT -17.355 -220.200 -17.155 -219.555 ;
        RECT -16.410 -220.200 -16.180 -219.555 ;
        RECT -15.395 -219.575 -15.225 -218.640 ;
        RECT -14.825 -219.555 -14.655 -218.640 ;
        RECT -15.420 -220.200 -15.190 -219.575 ;
        RECT -14.855 -220.200 -14.625 -219.555 ;
        RECT -13.845 -219.580 -13.675 -218.640 ;
        RECT -13.280 -219.530 -13.110 -218.640 ;
        RECT -13.875 -220.200 -13.645 -219.580 ;
        RECT -13.310 -220.200 -13.080 -219.530 ;
        RECT -12.300 -219.590 -12.130 -218.640 ;
        RECT -12.325 -220.200 -12.095 -219.590 ;
        RECT -17.355 -220.545 -12.095 -220.200 ;
        RECT -15.785 -220.735 -12.820 -220.545 ;
        RECT -10.380 -220.735 -9.810 -216.375 ;
        RECT -4.855 -219.555 -4.685 -218.640 ;
        RECT -3.875 -219.555 -3.705 -218.640 ;
        RECT -4.855 -220.200 -4.655 -219.555 ;
        RECT -3.910 -220.200 -3.680 -219.555 ;
        RECT -2.895 -219.575 -2.725 -218.640 ;
        RECT -2.325 -219.555 -2.155 -218.640 ;
        RECT -2.920 -220.200 -2.690 -219.575 ;
        RECT -2.355 -220.200 -2.125 -219.555 ;
        RECT -1.345 -219.580 -1.175 -218.640 ;
        RECT -0.780 -219.530 -0.610 -218.640 ;
        RECT -1.375 -220.200 -1.145 -219.580 ;
        RECT -0.810 -220.200 -0.580 -219.530 ;
        RECT 0.200 -219.590 0.370 -218.640 ;
        RECT 0.175 -220.200 0.405 -219.590 ;
        RECT -4.855 -220.545 0.405 -220.200 ;
        RECT -3.205 -220.735 -0.240 -220.545 ;
        RECT 2.030 -220.735 2.605 -216.375 ;
        RECT 7.645 -219.555 7.815 -218.640 ;
        RECT 8.625 -219.555 8.795 -218.640 ;
        RECT 7.645 -220.200 7.845 -219.555 ;
        RECT 8.590 -220.200 8.820 -219.555 ;
        RECT 9.605 -219.575 9.775 -218.640 ;
        RECT 10.175 -219.555 10.345 -218.640 ;
        RECT 9.580 -220.200 9.810 -219.575 ;
        RECT 10.145 -220.200 10.375 -219.555 ;
        RECT 11.155 -219.580 11.325 -218.640 ;
        RECT 11.720 -219.530 11.890 -218.640 ;
        RECT 11.125 -220.200 11.355 -219.580 ;
        RECT 11.690 -220.200 11.920 -219.530 ;
        RECT 12.700 -219.590 12.870 -218.640 ;
        RECT 20.145 -219.555 20.315 -218.640 ;
        RECT 21.125 -219.555 21.295 -218.640 ;
        RECT 12.675 -220.200 12.905 -219.590 ;
        RECT 7.645 -220.545 12.905 -220.200 ;
        RECT 20.145 -220.200 20.345 -219.555 ;
        RECT 21.090 -220.200 21.320 -219.555 ;
        RECT 22.105 -219.575 22.275 -218.640 ;
        RECT 22.675 -219.555 22.845 -218.640 ;
        RECT 22.080 -220.200 22.310 -219.575 ;
        RECT 22.645 -220.200 22.875 -219.555 ;
        RECT 23.655 -219.580 23.825 -218.640 ;
        RECT 24.220 -219.530 24.390 -218.640 ;
        RECT 23.625 -220.200 23.855 -219.580 ;
        RECT 24.190 -220.200 24.420 -219.530 ;
        RECT 25.200 -219.590 25.370 -218.640 ;
        RECT 35.145 -219.555 35.315 -218.640 ;
        RECT 36.125 -219.555 36.295 -218.640 ;
        RECT 25.175 -220.200 25.405 -219.590 ;
        RECT 20.145 -220.545 25.405 -220.200 ;
        RECT 35.145 -220.200 35.345 -219.555 ;
        RECT 36.090 -220.200 36.320 -219.555 ;
        RECT 37.105 -219.575 37.275 -218.640 ;
        RECT 37.675 -219.555 37.845 -218.640 ;
        RECT 37.080 -220.200 37.310 -219.575 ;
        RECT 37.645 -220.200 37.875 -219.555 ;
        RECT 38.655 -219.580 38.825 -218.640 ;
        RECT 39.220 -219.530 39.390 -218.640 ;
        RECT 38.625 -220.200 38.855 -219.580 ;
        RECT 39.190 -220.200 39.420 -219.530 ;
        RECT 40.200 -219.590 40.370 -218.640 ;
        RECT 65.780 -219.280 65.950 -217.825 ;
        RECT 66.760 -219.280 66.930 -217.825 ;
        RECT 67.740 -219.280 67.910 -217.825 ;
        RECT 69.965 -219.280 70.135 -217.825 ;
        RECT 70.945 -219.280 71.115 -217.825 ;
        RECT 71.925 -219.280 72.095 -217.825 ;
        RECT 79.280 -219.280 79.450 -217.825 ;
        RECT 80.260 -219.280 80.430 -217.825 ;
        RECT 81.240 -219.280 81.410 -217.825 ;
        RECT 83.465 -219.280 83.635 -217.825 ;
        RECT 84.445 -219.280 84.615 -217.825 ;
        RECT 85.425 -219.280 85.595 -217.825 ;
        RECT 86.395 -219.280 86.840 -210.805 ;
        RECT 145.345 -211.195 145.515 -208.245 ;
        RECT 146.325 -211.195 146.495 -208.230 ;
        RECT 148.405 -208.235 148.630 -207.615 ;
        RECT 156.400 -207.650 168.125 -207.440 ;
        RECT 158.410 -207.685 159.540 -207.650 ;
        RECT 158.595 -207.720 159.540 -207.685 ;
        RECT 163.630 -207.675 168.125 -207.650 ;
        RECT 163.630 -207.770 167.475 -207.675 ;
        RECT 156.400 -207.965 158.610 -207.890 ;
        RECT 156.400 -208.210 162.845 -207.965 ;
        RECT 148.440 -211.195 148.610 -208.235 ;
        RECT 156.450 -210.295 156.620 -208.210 ;
        RECT 157.430 -210.295 157.600 -208.210 ;
        RECT 158.410 -208.460 162.845 -208.210 ;
        RECT 163.660 -208.400 163.885 -207.770 ;
        RECT 164.635 -208.385 164.860 -207.770 ;
        RECT 158.410 -210.295 158.580 -208.460 ;
        RECT 159.495 -209.290 159.665 -208.460 ;
        RECT 160.475 -209.290 160.645 -208.460 ;
        RECT 161.455 -209.290 161.625 -208.460 ;
        RECT 162.435 -209.290 162.605 -208.460 ;
        RECT 163.685 -211.350 163.855 -208.400 ;
        RECT 164.665 -211.350 164.835 -208.385 ;
        RECT 166.745 -208.390 166.970 -207.770 ;
        RECT 167.730 -207.800 168.125 -207.675 ;
        RECT 168.980 -207.725 170.040 -207.030 ;
        RECT 180.260 -207.340 190.815 -206.785 ;
        RECT 192.915 -206.965 193.245 -200.460 ;
        RECT 180.260 -207.550 191.335 -207.340 ;
        RECT 192.830 -207.530 193.250 -206.965 ;
        RECT 194.595 -207.110 194.925 -200.460 ;
        RECT 209.080 -201.495 209.690 -189.960 ;
        RECT 224.615 -190.270 235.170 -189.960 ;
        RECT 240.010 -190.030 242.035 -189.710 ;
        RECT 237.195 -190.080 237.685 -190.065 ;
        RECT 240.010 -190.080 240.595 -190.030 ;
        RECT 224.615 -190.305 235.690 -190.270 ;
        RECT 236.055 -190.305 236.365 -190.165 ;
        RECT 224.615 -190.480 236.365 -190.305 ;
        RECT 226.625 -190.515 227.755 -190.480 ;
        RECT 226.810 -190.550 227.755 -190.515 ;
        RECT 231.845 -190.565 236.365 -190.480 ;
        RECT 231.845 -190.600 235.690 -190.565 ;
        RECT 224.615 -190.795 226.825 -190.720 ;
        RECT 224.615 -191.040 231.060 -190.795 ;
        RECT 224.665 -193.125 224.835 -191.040 ;
        RECT 225.645 -193.125 225.815 -191.040 ;
        RECT 226.625 -191.290 231.060 -191.040 ;
        RECT 231.875 -191.230 232.100 -190.600 ;
        RECT 232.850 -191.215 233.075 -190.600 ;
        RECT 226.625 -193.125 226.795 -191.290 ;
        RECT 227.710 -192.120 227.880 -191.290 ;
        RECT 228.690 -192.120 228.860 -191.290 ;
        RECT 229.670 -192.120 229.840 -191.290 ;
        RECT 230.650 -192.120 230.820 -191.290 ;
        RECT 231.900 -194.180 232.070 -191.230 ;
        RECT 232.880 -194.180 233.050 -191.215 ;
        RECT 234.960 -191.220 235.185 -190.600 ;
        RECT 236.055 -190.635 236.365 -190.565 ;
        RECT 237.195 -190.665 240.595 -190.080 ;
        RECT 241.845 -190.505 242.035 -190.030 ;
        RECT 242.830 -190.495 243.020 -189.710 ;
        RECT 237.195 -190.695 237.685 -190.665 ;
        RECT 234.995 -194.180 235.165 -191.220 ;
        RECT 241.860 -192.970 242.030 -190.505 ;
        RECT 242.840 -192.970 243.010 -190.495 ;
        RECT 245.790 -190.610 246.040 -189.710 ;
        RECT 246.420 -190.595 246.670 -189.710 ;
        RECT 247.575 -190.520 247.790 -189.710 ;
        RECT 248.560 -190.010 281.160 -189.710 ;
        RECT 286.000 -189.860 288.025 -189.540 ;
        RECT 283.185 -189.910 283.675 -189.895 ;
        RECT 286.000 -189.910 286.585 -189.860 ;
        RECT 248.560 -190.510 248.775 -190.010 ;
        RECT 245.815 -192.970 245.985 -190.610 ;
        RECT 246.465 -192.970 246.635 -190.595 ;
        RECT 247.605 -191.970 247.775 -190.520 ;
        RECT 248.585 -191.970 248.755 -190.510 ;
        RECT 237.230 -200.655 239.240 -200.325 ;
        RECT 209.080 -202.105 212.240 -201.495 ;
        RECT 198.780 -205.495 198.950 -204.165 ;
        RECT 199.760 -205.495 199.930 -204.165 ;
        RECT 200.740 -205.495 200.910 -204.165 ;
        RECT 201.720 -205.495 201.890 -204.165 ;
        RECT 198.540 -205.990 202.130 -205.495 ;
        RECT 199.450 -206.940 200.310 -205.990 ;
        RECT 203.645 -206.395 203.815 -204.310 ;
        RECT 204.625 -206.395 204.795 -204.310 ;
        RECT 205.605 -206.145 205.775 -204.310 ;
        RECT 206.690 -206.145 206.860 -205.315 ;
        RECT 207.670 -206.145 207.840 -205.315 ;
        RECT 208.650 -206.145 208.820 -205.315 ;
        RECT 209.630 -206.145 209.800 -205.315 ;
        RECT 205.605 -206.395 210.040 -206.145 ;
        RECT 203.595 -206.640 210.040 -206.395 ;
        RECT 203.595 -206.710 205.805 -206.640 ;
        RECT 203.590 -206.855 205.805 -206.710 ;
        RECT 203.590 -206.940 206.680 -206.855 ;
        RECT 198.600 -207.110 209.155 -206.940 ;
        RECT 211.630 -207.085 212.240 -202.105 ;
        RECT 224.755 -205.535 224.925 -204.205 ;
        RECT 225.735 -205.535 225.905 -204.205 ;
        RECT 226.715 -205.535 226.885 -204.205 ;
        RECT 227.695 -205.535 227.865 -204.205 ;
        RECT 224.515 -206.030 228.105 -205.535 ;
        RECT 225.425 -206.980 226.285 -206.030 ;
        RECT 229.620 -206.435 229.790 -204.350 ;
        RECT 230.600 -206.435 230.770 -204.350 ;
        RECT 231.580 -206.185 231.750 -204.350 ;
        RECT 232.665 -206.185 232.835 -205.355 ;
        RECT 233.645 -206.185 233.815 -205.355 ;
        RECT 234.625 -206.185 234.795 -205.355 ;
        RECT 235.605 -206.185 235.775 -205.355 ;
        RECT 231.580 -206.435 236.015 -206.185 ;
        RECT 229.570 -206.680 236.015 -206.435 ;
        RECT 229.570 -206.750 231.780 -206.680 ;
        RECT 229.565 -206.895 231.780 -206.750 ;
        RECT 229.565 -206.980 232.655 -206.895 ;
        RECT 194.595 -207.440 209.155 -207.110 ;
        RECT 209.930 -207.315 210.325 -207.160 ;
        RECT 198.600 -207.495 209.155 -207.440 ;
        RECT 209.430 -207.495 210.325 -207.315 ;
        RECT 182.270 -207.585 183.400 -207.550 ;
        RECT 182.455 -207.620 183.400 -207.585 ;
        RECT 187.490 -207.670 191.335 -207.550 ;
        RECT 168.980 -207.865 169.675 -207.725 ;
        RECT 180.260 -207.865 182.470 -207.790 ;
        RECT 180.260 -208.110 186.705 -207.865 ;
        RECT 166.780 -211.350 166.950 -208.390 ;
        RECT 180.310 -210.195 180.480 -208.110 ;
        RECT 181.290 -210.195 181.460 -208.110 ;
        RECT 182.270 -208.360 186.705 -208.110 ;
        RECT 187.520 -208.300 187.745 -207.670 ;
        RECT 188.495 -208.285 188.720 -207.670 ;
        RECT 182.270 -210.195 182.440 -208.360 ;
        RECT 183.355 -209.190 183.525 -208.360 ;
        RECT 184.335 -209.190 184.505 -208.360 ;
        RECT 185.315 -209.190 185.485 -208.360 ;
        RECT 186.295 -209.190 186.465 -208.360 ;
        RECT 187.545 -211.250 187.715 -208.300 ;
        RECT 188.525 -211.250 188.695 -208.285 ;
        RECT 190.605 -208.290 190.830 -207.670 ;
        RECT 198.600 -207.705 210.325 -207.495 ;
        RECT 200.610 -207.740 201.740 -207.705 ;
        RECT 200.795 -207.775 201.740 -207.740 ;
        RECT 205.830 -207.730 210.325 -207.705 ;
        RECT 205.830 -207.825 209.675 -207.730 ;
        RECT 198.600 -208.020 200.810 -207.945 ;
        RECT 198.600 -208.265 205.045 -208.020 ;
        RECT 190.640 -211.250 190.810 -208.290 ;
        RECT 198.650 -210.350 198.820 -208.265 ;
        RECT 199.630 -210.350 199.800 -208.265 ;
        RECT 200.610 -208.515 205.045 -208.265 ;
        RECT 205.860 -208.455 206.085 -207.825 ;
        RECT 206.835 -208.440 207.060 -207.825 ;
        RECT 200.610 -210.350 200.780 -208.515 ;
        RECT 201.695 -209.345 201.865 -208.515 ;
        RECT 202.675 -209.345 202.845 -208.515 ;
        RECT 203.655 -209.345 203.825 -208.515 ;
        RECT 204.635 -209.345 204.805 -208.515 ;
        RECT 205.885 -211.405 206.055 -208.455 ;
        RECT 206.865 -211.405 207.035 -208.440 ;
        RECT 208.945 -208.445 209.170 -207.825 ;
        RECT 209.930 -207.855 210.325 -207.730 ;
        RECT 211.180 -207.780 212.240 -207.085 ;
        RECT 224.575 -207.535 235.130 -206.980 ;
        RECT 237.230 -207.160 237.560 -200.655 ;
        RECT 224.575 -207.745 235.650 -207.535 ;
        RECT 237.145 -207.725 237.565 -207.160 ;
        RECT 238.910 -207.305 239.240 -200.655 ;
        RECT 253.395 -201.690 254.005 -190.010 ;
        RECT 270.605 -190.100 281.160 -190.010 ;
        RECT 270.605 -190.135 281.680 -190.100 ;
        RECT 282.045 -190.135 282.355 -189.995 ;
        RECT 270.605 -190.310 282.355 -190.135 ;
        RECT 272.615 -190.345 273.745 -190.310 ;
        RECT 272.800 -190.380 273.745 -190.345 ;
        RECT 277.835 -190.395 282.355 -190.310 ;
        RECT 277.835 -190.430 281.680 -190.395 ;
        RECT 270.605 -190.625 272.815 -190.550 ;
        RECT 270.605 -190.870 277.050 -190.625 ;
        RECT 270.655 -192.955 270.825 -190.870 ;
        RECT 271.635 -192.955 271.805 -190.870 ;
        RECT 272.615 -191.120 277.050 -190.870 ;
        RECT 277.865 -191.060 278.090 -190.430 ;
        RECT 278.840 -191.045 279.065 -190.430 ;
        RECT 272.615 -192.955 272.785 -191.120 ;
        RECT 273.700 -191.950 273.870 -191.120 ;
        RECT 274.680 -191.950 274.850 -191.120 ;
        RECT 275.660 -191.950 275.830 -191.120 ;
        RECT 276.640 -191.950 276.810 -191.120 ;
        RECT 277.890 -194.010 278.060 -191.060 ;
        RECT 278.870 -194.010 279.040 -191.045 ;
        RECT 280.950 -191.050 281.175 -190.430 ;
        RECT 282.045 -190.465 282.355 -190.395 ;
        RECT 283.185 -190.495 286.585 -189.910 ;
        RECT 287.835 -190.335 288.025 -189.860 ;
        RECT 288.820 -190.325 289.010 -189.540 ;
        RECT 283.185 -190.525 283.675 -190.495 ;
        RECT 280.985 -194.010 281.155 -191.050 ;
        RECT 287.850 -192.800 288.020 -190.335 ;
        RECT 288.830 -192.800 289.000 -190.325 ;
        RECT 291.780 -190.440 292.030 -189.540 ;
        RECT 292.410 -190.425 292.660 -189.540 ;
        RECT 293.565 -190.350 293.780 -189.540 ;
        RECT 294.550 -189.770 324.930 -189.540 ;
        RECT 329.770 -189.530 331.795 -189.210 ;
        RECT 326.955 -189.580 327.445 -189.565 ;
        RECT 329.770 -189.580 330.355 -189.530 ;
        RECT 294.550 -189.805 325.450 -189.770 ;
        RECT 325.815 -189.805 326.125 -189.665 ;
        RECT 294.550 -189.850 326.125 -189.805 ;
        RECT 294.550 -190.340 294.765 -189.850 ;
        RECT 291.805 -192.800 291.975 -190.440 ;
        RECT 292.455 -192.800 292.625 -190.425 ;
        RECT 293.595 -191.800 293.765 -190.350 ;
        RECT 294.575 -191.800 294.745 -190.340 ;
        RECT 283.220 -200.485 285.230 -200.155 ;
        RECT 253.395 -202.300 256.555 -201.690 ;
        RECT 243.095 -205.690 243.265 -204.360 ;
        RECT 244.075 -205.690 244.245 -204.360 ;
        RECT 245.055 -205.690 245.225 -204.360 ;
        RECT 246.035 -205.690 246.205 -204.360 ;
        RECT 242.855 -206.185 246.445 -205.690 ;
        RECT 243.765 -207.135 244.625 -206.185 ;
        RECT 247.960 -206.590 248.130 -204.505 ;
        RECT 248.940 -206.590 249.110 -204.505 ;
        RECT 249.920 -206.340 250.090 -204.505 ;
        RECT 251.005 -206.340 251.175 -205.510 ;
        RECT 251.985 -206.340 252.155 -205.510 ;
        RECT 252.965 -206.340 253.135 -205.510 ;
        RECT 253.945 -206.340 254.115 -205.510 ;
        RECT 249.920 -206.590 254.355 -206.340 ;
        RECT 247.910 -206.835 254.355 -206.590 ;
        RECT 247.910 -206.905 250.120 -206.835 ;
        RECT 247.905 -207.050 250.120 -206.905 ;
        RECT 247.905 -207.135 250.995 -207.050 ;
        RECT 242.915 -207.305 253.470 -207.135 ;
        RECT 255.945 -207.280 256.555 -202.300 ;
        RECT 270.745 -205.365 270.915 -204.035 ;
        RECT 271.725 -205.365 271.895 -204.035 ;
        RECT 272.705 -205.365 272.875 -204.035 ;
        RECT 273.685 -205.365 273.855 -204.035 ;
        RECT 270.505 -205.860 274.095 -205.365 ;
        RECT 271.415 -206.810 272.275 -205.860 ;
        RECT 275.610 -206.265 275.780 -204.180 ;
        RECT 276.590 -206.265 276.760 -204.180 ;
        RECT 277.570 -206.015 277.740 -204.180 ;
        RECT 278.655 -206.015 278.825 -205.185 ;
        RECT 279.635 -206.015 279.805 -205.185 ;
        RECT 280.615 -206.015 280.785 -205.185 ;
        RECT 281.595 -206.015 281.765 -205.185 ;
        RECT 277.570 -206.265 282.005 -206.015 ;
        RECT 275.560 -206.510 282.005 -206.265 ;
        RECT 275.560 -206.580 277.770 -206.510 ;
        RECT 275.555 -206.725 277.770 -206.580 ;
        RECT 275.555 -206.810 278.645 -206.725 ;
        RECT 238.910 -207.635 253.470 -207.305 ;
        RECT 254.245 -207.510 254.640 -207.355 ;
        RECT 242.915 -207.690 253.470 -207.635 ;
        RECT 253.745 -207.690 254.640 -207.510 ;
        RECT 226.585 -207.780 227.715 -207.745 ;
        RECT 211.180 -207.920 211.875 -207.780 ;
        RECT 226.770 -207.815 227.715 -207.780 ;
        RECT 231.805 -207.865 235.650 -207.745 ;
        RECT 224.575 -208.060 226.785 -207.985 ;
        RECT 224.575 -208.305 231.020 -208.060 ;
        RECT 208.980 -211.405 209.150 -208.445 ;
        RECT 224.625 -210.390 224.795 -208.305 ;
        RECT 225.605 -210.390 225.775 -208.305 ;
        RECT 226.585 -208.555 231.020 -208.305 ;
        RECT 231.835 -208.495 232.060 -207.865 ;
        RECT 232.810 -208.480 233.035 -207.865 ;
        RECT 226.585 -210.390 226.755 -208.555 ;
        RECT 227.670 -209.385 227.840 -208.555 ;
        RECT 228.650 -209.385 228.820 -208.555 ;
        RECT 229.630 -209.385 229.800 -208.555 ;
        RECT 230.610 -209.385 230.780 -208.555 ;
        RECT 231.860 -211.445 232.030 -208.495 ;
        RECT 232.840 -211.445 233.010 -208.480 ;
        RECT 234.920 -208.485 235.145 -207.865 ;
        RECT 242.915 -207.900 254.640 -207.690 ;
        RECT 244.925 -207.935 246.055 -207.900 ;
        RECT 245.110 -207.970 246.055 -207.935 ;
        RECT 250.145 -207.925 254.640 -207.900 ;
        RECT 250.145 -208.020 253.990 -207.925 ;
        RECT 242.915 -208.215 245.125 -208.140 ;
        RECT 242.915 -208.460 249.360 -208.215 ;
        RECT 234.955 -211.445 235.125 -208.485 ;
        RECT 242.965 -210.545 243.135 -208.460 ;
        RECT 243.945 -210.545 244.115 -208.460 ;
        RECT 244.925 -208.710 249.360 -208.460 ;
        RECT 250.175 -208.650 250.400 -208.020 ;
        RECT 251.150 -208.635 251.375 -208.020 ;
        RECT 244.925 -210.545 245.095 -208.710 ;
        RECT 246.010 -209.540 246.180 -208.710 ;
        RECT 246.990 -209.540 247.160 -208.710 ;
        RECT 247.970 -209.540 248.140 -208.710 ;
        RECT 248.950 -209.540 249.120 -208.710 ;
        RECT 250.200 -211.600 250.370 -208.650 ;
        RECT 251.180 -211.600 251.350 -208.635 ;
        RECT 253.260 -208.640 253.485 -208.020 ;
        RECT 254.245 -208.050 254.640 -207.925 ;
        RECT 255.495 -207.975 256.555 -207.280 ;
        RECT 270.565 -207.365 281.120 -206.810 ;
        RECT 283.220 -206.990 283.550 -200.485 ;
        RECT 270.565 -207.575 281.640 -207.365 ;
        RECT 283.135 -207.555 283.555 -206.990 ;
        RECT 284.900 -207.135 285.230 -200.485 ;
        RECT 299.385 -201.520 299.995 -189.850 ;
        RECT 314.375 -189.980 326.125 -189.850 ;
        RECT 316.385 -190.015 317.515 -189.980 ;
        RECT 316.570 -190.050 317.515 -190.015 ;
        RECT 321.605 -190.065 326.125 -189.980 ;
        RECT 321.605 -190.100 325.450 -190.065 ;
        RECT 314.375 -190.295 316.585 -190.220 ;
        RECT 314.375 -190.540 320.820 -190.295 ;
        RECT 314.425 -192.625 314.595 -190.540 ;
        RECT 315.405 -192.625 315.575 -190.540 ;
        RECT 316.385 -190.790 320.820 -190.540 ;
        RECT 321.635 -190.730 321.860 -190.100 ;
        RECT 322.610 -190.715 322.835 -190.100 ;
        RECT 316.385 -192.625 316.555 -190.790 ;
        RECT 317.470 -191.620 317.640 -190.790 ;
        RECT 318.450 -191.620 318.620 -190.790 ;
        RECT 319.430 -191.620 319.600 -190.790 ;
        RECT 320.410 -191.620 320.580 -190.790 ;
        RECT 321.660 -193.680 321.830 -190.730 ;
        RECT 322.640 -193.680 322.810 -190.715 ;
        RECT 324.720 -190.720 324.945 -190.100 ;
        RECT 325.815 -190.135 326.125 -190.065 ;
        RECT 326.955 -190.165 330.355 -189.580 ;
        RECT 331.605 -190.005 331.795 -189.530 ;
        RECT 332.590 -189.995 332.780 -189.210 ;
        RECT 326.955 -190.195 327.445 -190.165 ;
        RECT 324.755 -193.680 324.925 -190.720 ;
        RECT 331.620 -192.470 331.790 -190.005 ;
        RECT 332.600 -192.470 332.770 -189.995 ;
        RECT 335.550 -190.110 335.800 -189.210 ;
        RECT 336.180 -190.095 336.430 -189.210 ;
        RECT 337.335 -190.020 337.550 -189.210 ;
        RECT 338.295 -189.380 370.695 -189.210 ;
        RECT 338.320 -190.010 338.535 -189.380 ;
        RECT 335.575 -192.470 335.745 -190.110 ;
        RECT 336.225 -192.470 336.395 -190.095 ;
        RECT 337.365 -191.470 337.535 -190.020 ;
        RECT 338.345 -191.470 338.515 -190.010 ;
        RECT 326.990 -200.155 329.000 -199.825 ;
        RECT 299.385 -202.130 302.545 -201.520 ;
        RECT 289.085 -205.520 289.255 -204.190 ;
        RECT 290.065 -205.520 290.235 -204.190 ;
        RECT 291.045 -205.520 291.215 -204.190 ;
        RECT 292.025 -205.520 292.195 -204.190 ;
        RECT 288.845 -206.015 292.435 -205.520 ;
        RECT 289.755 -206.965 290.615 -206.015 ;
        RECT 293.950 -206.420 294.120 -204.335 ;
        RECT 294.930 -206.420 295.100 -204.335 ;
        RECT 295.910 -206.170 296.080 -204.335 ;
        RECT 296.995 -206.170 297.165 -205.340 ;
        RECT 297.975 -206.170 298.145 -205.340 ;
        RECT 298.955 -206.170 299.125 -205.340 ;
        RECT 299.935 -206.170 300.105 -205.340 ;
        RECT 295.910 -206.420 300.345 -206.170 ;
        RECT 293.900 -206.665 300.345 -206.420 ;
        RECT 293.900 -206.735 296.110 -206.665 ;
        RECT 293.895 -206.880 296.110 -206.735 ;
        RECT 293.895 -206.965 296.985 -206.880 ;
        RECT 288.905 -207.135 299.460 -206.965 ;
        RECT 301.935 -207.110 302.545 -202.130 ;
        RECT 314.515 -205.035 314.685 -203.705 ;
        RECT 315.495 -205.035 315.665 -203.705 ;
        RECT 316.475 -205.035 316.645 -203.705 ;
        RECT 317.455 -205.035 317.625 -203.705 ;
        RECT 314.275 -205.530 317.865 -205.035 ;
        RECT 315.185 -206.480 316.045 -205.530 ;
        RECT 319.380 -205.935 319.550 -203.850 ;
        RECT 320.360 -205.935 320.530 -203.850 ;
        RECT 321.340 -205.685 321.510 -203.850 ;
        RECT 322.425 -205.685 322.595 -204.855 ;
        RECT 323.405 -205.685 323.575 -204.855 ;
        RECT 324.385 -205.685 324.555 -204.855 ;
        RECT 325.365 -205.685 325.535 -204.855 ;
        RECT 321.340 -205.935 325.775 -205.685 ;
        RECT 319.330 -206.180 325.775 -205.935 ;
        RECT 319.330 -206.250 321.540 -206.180 ;
        RECT 319.325 -206.395 321.540 -206.250 ;
        RECT 319.325 -206.480 322.415 -206.395 ;
        RECT 284.900 -207.465 299.460 -207.135 ;
        RECT 300.235 -207.340 300.630 -207.185 ;
        RECT 288.905 -207.520 299.460 -207.465 ;
        RECT 299.735 -207.520 300.630 -207.340 ;
        RECT 272.575 -207.610 273.705 -207.575 ;
        RECT 272.760 -207.645 273.705 -207.610 ;
        RECT 277.795 -207.695 281.640 -207.575 ;
        RECT 270.565 -207.890 272.775 -207.815 ;
        RECT 255.495 -208.115 256.190 -207.975 ;
        RECT 270.565 -208.135 277.010 -207.890 ;
        RECT 253.295 -211.600 253.465 -208.640 ;
        RECT 270.615 -210.220 270.785 -208.135 ;
        RECT 271.595 -210.220 271.765 -208.135 ;
        RECT 272.575 -208.385 277.010 -208.135 ;
        RECT 277.825 -208.325 278.050 -207.695 ;
        RECT 278.800 -208.310 279.025 -207.695 ;
        RECT 272.575 -210.220 272.745 -208.385 ;
        RECT 273.660 -209.215 273.830 -208.385 ;
        RECT 274.640 -209.215 274.810 -208.385 ;
        RECT 275.620 -209.215 275.790 -208.385 ;
        RECT 276.600 -209.215 276.770 -208.385 ;
        RECT 277.850 -211.275 278.020 -208.325 ;
        RECT 278.830 -211.275 279.000 -208.310 ;
        RECT 280.910 -208.315 281.135 -207.695 ;
        RECT 288.905 -207.730 300.630 -207.520 ;
        RECT 290.915 -207.765 292.045 -207.730 ;
        RECT 291.100 -207.800 292.045 -207.765 ;
        RECT 296.135 -207.755 300.630 -207.730 ;
        RECT 296.135 -207.850 299.980 -207.755 ;
        RECT 288.905 -208.045 291.115 -207.970 ;
        RECT 288.905 -208.290 295.350 -208.045 ;
        RECT 280.945 -211.275 281.115 -208.315 ;
        RECT 288.955 -210.375 289.125 -208.290 ;
        RECT 289.935 -210.375 290.105 -208.290 ;
        RECT 290.915 -208.540 295.350 -208.290 ;
        RECT 296.165 -208.480 296.390 -207.850 ;
        RECT 297.140 -208.465 297.365 -207.850 ;
        RECT 290.915 -210.375 291.085 -208.540 ;
        RECT 292.000 -209.370 292.170 -208.540 ;
        RECT 292.980 -209.370 293.150 -208.540 ;
        RECT 293.960 -209.370 294.130 -208.540 ;
        RECT 294.940 -209.370 295.110 -208.540 ;
        RECT 296.190 -211.430 296.360 -208.480 ;
        RECT 297.170 -211.430 297.340 -208.465 ;
        RECT 299.250 -208.470 299.475 -207.850 ;
        RECT 300.235 -207.880 300.630 -207.755 ;
        RECT 301.485 -207.805 302.545 -207.110 ;
        RECT 314.335 -207.035 324.890 -206.480 ;
        RECT 326.990 -206.660 327.320 -200.155 ;
        RECT 314.335 -207.245 325.410 -207.035 ;
        RECT 326.905 -207.225 327.325 -206.660 ;
        RECT 328.670 -206.805 329.000 -200.155 ;
        RECT 343.155 -201.190 343.765 -189.380 ;
        RECT 360.140 -189.685 370.695 -189.380 ;
        RECT 375.535 -189.445 377.560 -189.125 ;
        RECT 372.720 -189.495 373.210 -189.480 ;
        RECT 375.535 -189.495 376.120 -189.445 ;
        RECT 360.140 -189.720 371.215 -189.685 ;
        RECT 371.580 -189.720 371.890 -189.580 ;
        RECT 360.140 -189.895 371.890 -189.720 ;
        RECT 362.150 -189.930 363.280 -189.895 ;
        RECT 362.335 -189.965 363.280 -189.930 ;
        RECT 367.370 -189.980 371.890 -189.895 ;
        RECT 367.370 -190.015 371.215 -189.980 ;
        RECT 360.140 -190.210 362.350 -190.135 ;
        RECT 360.140 -190.455 366.585 -190.210 ;
        RECT 360.190 -192.540 360.360 -190.455 ;
        RECT 361.170 -192.540 361.340 -190.455 ;
        RECT 362.150 -190.705 366.585 -190.455 ;
        RECT 367.400 -190.645 367.625 -190.015 ;
        RECT 368.375 -190.630 368.600 -190.015 ;
        RECT 362.150 -192.540 362.320 -190.705 ;
        RECT 363.235 -191.535 363.405 -190.705 ;
        RECT 364.215 -191.535 364.385 -190.705 ;
        RECT 365.195 -191.535 365.365 -190.705 ;
        RECT 366.175 -191.535 366.345 -190.705 ;
        RECT 367.425 -193.595 367.595 -190.645 ;
        RECT 368.405 -193.595 368.575 -190.630 ;
        RECT 370.485 -190.635 370.710 -190.015 ;
        RECT 371.580 -190.050 371.890 -189.980 ;
        RECT 372.720 -190.080 376.120 -189.495 ;
        RECT 377.370 -189.920 377.560 -189.445 ;
        RECT 378.355 -189.910 378.545 -189.125 ;
        RECT 372.720 -190.110 373.210 -190.080 ;
        RECT 370.520 -193.595 370.690 -190.635 ;
        RECT 377.385 -192.385 377.555 -189.920 ;
        RECT 378.365 -192.385 378.535 -189.910 ;
        RECT 381.315 -190.025 381.565 -189.125 ;
        RECT 381.945 -190.010 382.195 -189.125 ;
        RECT 383.100 -189.935 383.315 -189.125 ;
        RECT 384.085 -189.425 417.515 -189.125 ;
        RECT 422.355 -189.255 424.380 -188.935 ;
        RECT 419.540 -189.305 420.030 -189.290 ;
        RECT 422.355 -189.305 422.940 -189.255 ;
        RECT 384.085 -189.925 384.300 -189.425 ;
        RECT 381.340 -192.385 381.510 -190.025 ;
        RECT 381.990 -192.385 382.160 -190.010 ;
        RECT 383.130 -191.385 383.300 -189.935 ;
        RECT 384.110 -191.385 384.280 -189.925 ;
        RECT 372.755 -200.070 374.765 -199.740 ;
        RECT 343.155 -201.800 346.315 -201.190 ;
        RECT 332.855 -205.190 333.025 -203.860 ;
        RECT 333.835 -205.190 334.005 -203.860 ;
        RECT 334.815 -205.190 334.985 -203.860 ;
        RECT 335.795 -205.190 335.965 -203.860 ;
        RECT 332.615 -205.685 336.205 -205.190 ;
        RECT 333.525 -206.635 334.385 -205.685 ;
        RECT 337.720 -206.090 337.890 -204.005 ;
        RECT 338.700 -206.090 338.870 -204.005 ;
        RECT 339.680 -205.840 339.850 -204.005 ;
        RECT 340.765 -205.840 340.935 -205.010 ;
        RECT 341.745 -205.840 341.915 -205.010 ;
        RECT 342.725 -205.840 342.895 -205.010 ;
        RECT 343.705 -205.840 343.875 -205.010 ;
        RECT 339.680 -206.090 344.115 -205.840 ;
        RECT 337.670 -206.335 344.115 -206.090 ;
        RECT 337.670 -206.405 339.880 -206.335 ;
        RECT 337.665 -206.550 339.880 -206.405 ;
        RECT 337.665 -206.635 340.755 -206.550 ;
        RECT 332.675 -206.805 343.230 -206.635 ;
        RECT 345.705 -206.780 346.315 -201.800 ;
        RECT 360.280 -204.950 360.450 -203.620 ;
        RECT 361.260 -204.950 361.430 -203.620 ;
        RECT 362.240 -204.950 362.410 -203.620 ;
        RECT 363.220 -204.950 363.390 -203.620 ;
        RECT 360.040 -205.445 363.630 -204.950 ;
        RECT 360.950 -206.395 361.810 -205.445 ;
        RECT 365.145 -205.850 365.315 -203.765 ;
        RECT 366.125 -205.850 366.295 -203.765 ;
        RECT 367.105 -205.600 367.275 -203.765 ;
        RECT 368.190 -205.600 368.360 -204.770 ;
        RECT 369.170 -205.600 369.340 -204.770 ;
        RECT 370.150 -205.600 370.320 -204.770 ;
        RECT 371.130 -205.600 371.300 -204.770 ;
        RECT 367.105 -205.850 371.540 -205.600 ;
        RECT 365.095 -206.095 371.540 -205.850 ;
        RECT 365.095 -206.165 367.305 -206.095 ;
        RECT 365.090 -206.310 367.305 -206.165 ;
        RECT 365.090 -206.395 368.180 -206.310 ;
        RECT 328.670 -207.135 343.230 -206.805 ;
        RECT 344.005 -207.010 344.400 -206.855 ;
        RECT 332.675 -207.190 343.230 -207.135 ;
        RECT 343.505 -207.190 344.400 -207.010 ;
        RECT 316.345 -207.280 317.475 -207.245 ;
        RECT 316.530 -207.315 317.475 -207.280 ;
        RECT 321.565 -207.365 325.410 -207.245 ;
        RECT 314.335 -207.560 316.545 -207.485 ;
        RECT 314.335 -207.805 320.780 -207.560 ;
        RECT 301.485 -207.945 302.180 -207.805 ;
        RECT 299.285 -211.430 299.455 -208.470 ;
        RECT 314.385 -209.890 314.555 -207.805 ;
        RECT 315.365 -209.890 315.535 -207.805 ;
        RECT 316.345 -208.055 320.780 -207.805 ;
        RECT 321.595 -207.995 321.820 -207.365 ;
        RECT 322.570 -207.980 322.795 -207.365 ;
        RECT 316.345 -209.890 316.515 -208.055 ;
        RECT 317.430 -208.885 317.600 -208.055 ;
        RECT 318.410 -208.885 318.580 -208.055 ;
        RECT 319.390 -208.885 319.560 -208.055 ;
        RECT 320.370 -208.885 320.540 -208.055 ;
        RECT 321.620 -210.945 321.790 -207.995 ;
        RECT 322.600 -210.945 322.770 -207.980 ;
        RECT 324.680 -207.985 324.905 -207.365 ;
        RECT 332.675 -207.400 344.400 -207.190 ;
        RECT 334.685 -207.435 335.815 -207.400 ;
        RECT 334.870 -207.470 335.815 -207.435 ;
        RECT 339.905 -207.425 344.400 -207.400 ;
        RECT 339.905 -207.520 343.750 -207.425 ;
        RECT 332.675 -207.715 334.885 -207.640 ;
        RECT 332.675 -207.960 339.120 -207.715 ;
        RECT 324.715 -210.945 324.885 -207.985 ;
        RECT 332.725 -210.045 332.895 -207.960 ;
        RECT 333.705 -210.045 333.875 -207.960 ;
        RECT 334.685 -208.210 339.120 -207.960 ;
        RECT 339.935 -208.150 340.160 -207.520 ;
        RECT 340.910 -208.135 341.135 -207.520 ;
        RECT 334.685 -210.045 334.855 -208.210 ;
        RECT 335.770 -209.040 335.940 -208.210 ;
        RECT 336.750 -209.040 336.920 -208.210 ;
        RECT 337.730 -209.040 337.900 -208.210 ;
        RECT 338.710 -209.040 338.880 -208.210 ;
        RECT 339.960 -211.100 340.130 -208.150 ;
        RECT 340.940 -211.100 341.110 -208.135 ;
        RECT 343.020 -208.140 343.245 -207.520 ;
        RECT 344.005 -207.550 344.400 -207.425 ;
        RECT 345.255 -207.475 346.315 -206.780 ;
        RECT 360.100 -206.950 370.655 -206.395 ;
        RECT 372.755 -206.575 373.085 -200.070 ;
        RECT 360.100 -207.160 371.175 -206.950 ;
        RECT 372.670 -207.140 373.090 -206.575 ;
        RECT 374.435 -206.720 374.765 -200.070 ;
        RECT 388.920 -201.105 389.530 -189.425 ;
        RECT 406.960 -189.495 417.515 -189.425 ;
        RECT 406.960 -189.530 418.035 -189.495 ;
        RECT 418.400 -189.530 418.710 -189.390 ;
        RECT 406.960 -189.705 418.710 -189.530 ;
        RECT 408.970 -189.740 410.100 -189.705 ;
        RECT 409.155 -189.775 410.100 -189.740 ;
        RECT 414.190 -189.790 418.710 -189.705 ;
        RECT 414.190 -189.825 418.035 -189.790 ;
        RECT 406.960 -190.020 409.170 -189.945 ;
        RECT 406.960 -190.265 413.405 -190.020 ;
        RECT 407.010 -192.350 407.180 -190.265 ;
        RECT 407.990 -192.350 408.160 -190.265 ;
        RECT 408.970 -190.515 413.405 -190.265 ;
        RECT 414.220 -190.455 414.445 -189.825 ;
        RECT 415.195 -190.440 415.420 -189.825 ;
        RECT 408.970 -192.350 409.140 -190.515 ;
        RECT 410.055 -191.345 410.225 -190.515 ;
        RECT 411.035 -191.345 411.205 -190.515 ;
        RECT 412.015 -191.345 412.185 -190.515 ;
        RECT 412.995 -191.345 413.165 -190.515 ;
        RECT 414.245 -193.405 414.415 -190.455 ;
        RECT 415.225 -193.405 415.395 -190.440 ;
        RECT 417.305 -190.445 417.530 -189.825 ;
        RECT 418.400 -189.860 418.710 -189.790 ;
        RECT 419.540 -189.890 422.940 -189.305 ;
        RECT 424.190 -189.730 424.380 -189.255 ;
        RECT 425.175 -189.720 425.365 -188.935 ;
        RECT 419.540 -189.920 420.030 -189.890 ;
        RECT 417.340 -193.405 417.510 -190.445 ;
        RECT 424.205 -192.195 424.375 -189.730 ;
        RECT 425.185 -192.195 425.355 -189.720 ;
        RECT 428.135 -189.835 428.385 -188.935 ;
        RECT 428.765 -189.820 429.015 -188.935 ;
        RECT 429.920 -189.745 430.135 -188.935 ;
        RECT 430.905 -189.735 431.120 -188.935 ;
        RECT 428.160 -192.195 428.330 -189.835 ;
        RECT 428.810 -192.195 428.980 -189.820 ;
        RECT 429.950 -191.195 430.120 -189.745 ;
        RECT 430.930 -191.195 431.100 -189.735 ;
        RECT 419.575 -199.880 421.585 -199.550 ;
        RECT 388.920 -201.715 392.080 -201.105 ;
        RECT 378.620 -205.105 378.790 -203.775 ;
        RECT 379.600 -205.105 379.770 -203.775 ;
        RECT 380.580 -205.105 380.750 -203.775 ;
        RECT 381.560 -205.105 381.730 -203.775 ;
        RECT 378.380 -205.600 381.970 -205.105 ;
        RECT 379.290 -206.550 380.150 -205.600 ;
        RECT 383.485 -206.005 383.655 -203.920 ;
        RECT 384.465 -206.005 384.635 -203.920 ;
        RECT 385.445 -205.755 385.615 -203.920 ;
        RECT 386.530 -205.755 386.700 -204.925 ;
        RECT 387.510 -205.755 387.680 -204.925 ;
        RECT 388.490 -205.755 388.660 -204.925 ;
        RECT 389.470 -205.755 389.640 -204.925 ;
        RECT 385.445 -206.005 389.880 -205.755 ;
        RECT 383.435 -206.250 389.880 -206.005 ;
        RECT 383.435 -206.320 385.645 -206.250 ;
        RECT 383.430 -206.465 385.645 -206.320 ;
        RECT 383.430 -206.550 386.520 -206.465 ;
        RECT 378.440 -206.720 388.995 -206.550 ;
        RECT 391.470 -206.695 392.080 -201.715 ;
        RECT 407.100 -204.760 407.270 -203.430 ;
        RECT 408.080 -204.760 408.250 -203.430 ;
        RECT 409.060 -204.760 409.230 -203.430 ;
        RECT 410.040 -204.760 410.210 -203.430 ;
        RECT 406.860 -205.255 410.450 -204.760 ;
        RECT 407.770 -206.205 408.630 -205.255 ;
        RECT 411.965 -205.660 412.135 -203.575 ;
        RECT 412.945 -205.660 413.115 -203.575 ;
        RECT 413.925 -205.410 414.095 -203.575 ;
        RECT 415.010 -205.410 415.180 -204.580 ;
        RECT 415.990 -205.410 416.160 -204.580 ;
        RECT 416.970 -205.410 417.140 -204.580 ;
        RECT 417.950 -205.410 418.120 -204.580 ;
        RECT 413.925 -205.660 418.360 -205.410 ;
        RECT 411.915 -205.905 418.360 -205.660 ;
        RECT 411.915 -205.975 414.125 -205.905 ;
        RECT 411.910 -206.120 414.125 -205.975 ;
        RECT 411.910 -206.205 415.000 -206.120 ;
        RECT 374.435 -207.050 388.995 -206.720 ;
        RECT 389.770 -206.925 390.165 -206.770 ;
        RECT 378.440 -207.105 388.995 -207.050 ;
        RECT 389.270 -207.105 390.165 -206.925 ;
        RECT 362.110 -207.195 363.240 -207.160 ;
        RECT 362.295 -207.230 363.240 -207.195 ;
        RECT 367.330 -207.280 371.175 -207.160 ;
        RECT 360.100 -207.475 362.310 -207.400 ;
        RECT 345.255 -207.615 345.950 -207.475 ;
        RECT 360.100 -207.720 366.545 -207.475 ;
        RECT 343.055 -211.100 343.225 -208.140 ;
        RECT 360.150 -209.805 360.320 -207.720 ;
        RECT 361.130 -209.805 361.300 -207.720 ;
        RECT 362.110 -207.970 366.545 -207.720 ;
        RECT 367.360 -207.910 367.585 -207.280 ;
        RECT 368.335 -207.895 368.560 -207.280 ;
        RECT 362.110 -209.805 362.280 -207.970 ;
        RECT 363.195 -208.800 363.365 -207.970 ;
        RECT 364.175 -208.800 364.345 -207.970 ;
        RECT 365.155 -208.800 365.325 -207.970 ;
        RECT 366.135 -208.800 366.305 -207.970 ;
        RECT 367.385 -210.860 367.555 -207.910 ;
        RECT 368.365 -210.860 368.535 -207.895 ;
        RECT 370.445 -207.900 370.670 -207.280 ;
        RECT 378.440 -207.315 390.165 -207.105 ;
        RECT 380.450 -207.350 381.580 -207.315 ;
        RECT 380.635 -207.385 381.580 -207.350 ;
        RECT 385.670 -207.340 390.165 -207.315 ;
        RECT 385.670 -207.435 389.515 -207.340 ;
        RECT 378.440 -207.630 380.650 -207.555 ;
        RECT 378.440 -207.875 384.885 -207.630 ;
        RECT 370.480 -210.860 370.650 -207.900 ;
        RECT 378.490 -209.960 378.660 -207.875 ;
        RECT 379.470 -209.960 379.640 -207.875 ;
        RECT 380.450 -208.125 384.885 -207.875 ;
        RECT 385.700 -208.065 385.925 -207.435 ;
        RECT 386.675 -208.050 386.900 -207.435 ;
        RECT 380.450 -209.960 380.620 -208.125 ;
        RECT 381.535 -208.955 381.705 -208.125 ;
        RECT 382.515 -208.955 382.685 -208.125 ;
        RECT 383.495 -208.955 383.665 -208.125 ;
        RECT 384.475 -208.955 384.645 -208.125 ;
        RECT 385.725 -211.015 385.895 -208.065 ;
        RECT 386.705 -211.015 386.875 -208.050 ;
        RECT 388.785 -208.055 389.010 -207.435 ;
        RECT 389.770 -207.465 390.165 -207.340 ;
        RECT 391.020 -207.390 392.080 -206.695 ;
        RECT 406.920 -206.760 417.475 -206.205 ;
        RECT 419.575 -206.385 419.905 -199.880 ;
        RECT 406.920 -206.970 417.995 -206.760 ;
        RECT 419.490 -206.950 419.910 -206.385 ;
        RECT 421.255 -206.530 421.585 -199.880 ;
        RECT 435.740 -200.915 436.350 -188.930 ;
        RECT 435.740 -201.525 438.900 -200.915 ;
        RECT 425.440 -204.915 425.610 -203.585 ;
        RECT 426.420 -204.915 426.590 -203.585 ;
        RECT 427.400 -204.915 427.570 -203.585 ;
        RECT 428.380 -204.915 428.550 -203.585 ;
        RECT 425.200 -205.410 428.790 -204.915 ;
        RECT 426.110 -206.360 426.970 -205.410 ;
        RECT 430.305 -205.815 430.475 -203.730 ;
        RECT 431.285 -205.815 431.455 -203.730 ;
        RECT 432.265 -205.565 432.435 -203.730 ;
        RECT 433.350 -205.565 433.520 -204.735 ;
        RECT 434.330 -205.565 434.500 -204.735 ;
        RECT 435.310 -205.565 435.480 -204.735 ;
        RECT 436.290 -205.565 436.460 -204.735 ;
        RECT 432.265 -205.815 436.700 -205.565 ;
        RECT 430.255 -206.060 436.700 -205.815 ;
        RECT 430.255 -206.130 432.465 -206.060 ;
        RECT 430.250 -206.275 432.465 -206.130 ;
        RECT 430.250 -206.360 433.340 -206.275 ;
        RECT 425.260 -206.530 435.815 -206.360 ;
        RECT 438.290 -206.505 438.900 -201.525 ;
        RECT 421.255 -206.860 435.815 -206.530 ;
        RECT 436.590 -206.735 436.985 -206.580 ;
        RECT 425.260 -206.915 435.815 -206.860 ;
        RECT 436.090 -206.915 436.985 -206.735 ;
        RECT 408.930 -207.005 410.060 -206.970 ;
        RECT 409.115 -207.040 410.060 -207.005 ;
        RECT 414.150 -207.090 417.995 -206.970 ;
        RECT 406.920 -207.285 409.130 -207.210 ;
        RECT 391.020 -207.530 391.715 -207.390 ;
        RECT 406.920 -207.530 413.365 -207.285 ;
        RECT 388.820 -211.015 388.990 -208.055 ;
        RECT 406.970 -209.615 407.140 -207.530 ;
        RECT 407.950 -209.615 408.120 -207.530 ;
        RECT 408.930 -207.780 413.365 -207.530 ;
        RECT 414.180 -207.720 414.405 -207.090 ;
        RECT 415.155 -207.705 415.380 -207.090 ;
        RECT 408.930 -209.615 409.100 -207.780 ;
        RECT 410.015 -208.610 410.185 -207.780 ;
        RECT 410.995 -208.610 411.165 -207.780 ;
        RECT 411.975 -208.610 412.145 -207.780 ;
        RECT 412.955 -208.610 413.125 -207.780 ;
        RECT 414.205 -210.670 414.375 -207.720 ;
        RECT 415.185 -210.670 415.355 -207.705 ;
        RECT 417.265 -207.710 417.490 -207.090 ;
        RECT 425.260 -207.125 436.985 -206.915 ;
        RECT 427.270 -207.160 428.400 -207.125 ;
        RECT 427.455 -207.195 428.400 -207.160 ;
        RECT 432.490 -207.150 436.985 -207.125 ;
        RECT 432.490 -207.245 436.335 -207.150 ;
        RECT 425.260 -207.440 427.470 -207.365 ;
        RECT 425.260 -207.685 431.705 -207.440 ;
        RECT 417.300 -210.670 417.470 -207.710 ;
        RECT 425.310 -209.770 425.480 -207.685 ;
        RECT 426.290 -209.770 426.460 -207.685 ;
        RECT 427.270 -207.935 431.705 -207.685 ;
        RECT 432.520 -207.875 432.745 -207.245 ;
        RECT 433.495 -207.860 433.720 -207.245 ;
        RECT 427.270 -209.770 427.440 -207.935 ;
        RECT 428.355 -208.765 428.525 -207.935 ;
        RECT 429.335 -208.765 429.505 -207.935 ;
        RECT 430.315 -208.765 430.485 -207.935 ;
        RECT 431.295 -208.765 431.465 -207.935 ;
        RECT 432.545 -210.825 432.715 -207.875 ;
        RECT 433.525 -210.825 433.695 -207.860 ;
        RECT 435.605 -207.865 435.830 -207.245 ;
        RECT 436.590 -207.275 436.985 -207.150 ;
        RECT 437.840 -207.200 438.900 -206.505 ;
        RECT 437.840 -207.340 438.535 -207.200 ;
        RECT 435.640 -210.825 435.810 -207.865 ;
        RECT 65.475 -219.305 74.485 -219.280 ;
        RECT 78.975 -219.305 86.840 -219.280 ;
        RECT 40.175 -220.200 40.405 -219.590 ;
        RECT 60.715 -219.620 86.840 -219.305 ;
        RECT 9.465 -220.735 12.430 -220.545 ;
        RECT 21.530 -220.735 24.495 -220.545 ;
        RECT 35.145 -220.735 40.405 -220.200 ;
        RECT -110.385 -220.910 -97.375 -220.865 ;
        RECT -34.180 -221.700 40.630 -220.735 ;
        RECT 479.145 -230.565 493.990 -156.540 ;
        RECT 416.665 -245.410 493.990 -230.565 ;
        RECT 416.665 -253.800 431.510 -245.410 ;
        RECT 133.130 -254.905 438.870 -253.800 ;
        RECT 37.990 -258.715 438.870 -254.905 ;
        RECT -136.945 -261.410 -136.705 -260.580 ;
        RECT -139.180 -261.580 -136.705 -261.410 ;
        RECT -136.945 -262.590 -136.705 -261.580 ;
        RECT -139.180 -262.760 -136.705 -262.590 ;
        RECT -136.945 -263.770 -136.705 -262.760 ;
        RECT -139.180 -263.940 -136.705 -263.770 ;
        RECT -136.945 -264.950 -136.705 -263.940 ;
        RECT -139.180 -265.120 -136.705 -264.950 ;
        RECT -136.945 -266.070 -136.705 -265.120 ;
        RECT -136.345 -266.070 -136.015 -261.130 ;
        RECT 37.990 -264.485 41.800 -258.715 ;
        RECT 133.130 -259.315 438.870 -258.715 ;
        RECT -33.155 -264.540 44.145 -264.485 ;
        RECT -44.810 -264.720 44.145 -264.540 ;
        RECT -136.945 -266.130 -136.015 -266.070 ;
        RECT -139.180 -266.300 -136.015 -266.130 ;
        RECT -136.945 -266.365 -136.015 -266.300 ;
        RECT -136.945 -267.310 -136.705 -266.365 ;
        RECT -139.180 -267.480 -136.705 -267.310 ;
        RECT -136.945 -268.455 -136.705 -267.480 ;
        RECT -136.345 -268.455 -136.015 -266.365 ;
        RECT -69.935 -264.985 44.145 -264.720 ;
        RECT -69.935 -265.035 -43.810 -264.985 ;
        RECT -69.935 -265.060 -62.070 -265.035 ;
        RECT -57.580 -265.060 -48.570 -265.035 ;
        RECT -69.935 -267.855 -69.490 -265.060 ;
        RECT -68.690 -266.515 -68.520 -265.060 ;
        RECT -67.710 -266.515 -67.540 -265.060 ;
        RECT -66.730 -266.515 -66.560 -265.060 ;
        RECT -64.505 -266.515 -64.335 -265.060 ;
        RECT -63.525 -266.515 -63.355 -265.060 ;
        RECT -62.545 -266.515 -62.375 -265.060 ;
        RECT -55.190 -266.515 -55.020 -265.060 ;
        RECT -54.210 -266.515 -54.040 -265.060 ;
        RECT -53.230 -266.515 -53.060 -265.060 ;
        RECT -51.005 -266.515 -50.835 -265.060 ;
        RECT -50.025 -266.515 -49.855 -265.060 ;
        RECT -49.045 -266.515 -48.875 -265.060 ;
        RECT -36.900 -265.605 -36.675 -264.985 ;
        RECT -34.790 -265.600 -34.565 -264.985 ;
        RECT -136.945 -268.490 -136.015 -268.455 ;
        RECT -139.180 -268.660 -136.015 -268.490 ;
        RECT -136.945 -268.750 -136.015 -268.660 ;
        RECT -136.945 -269.610 -136.705 -268.750 ;
        RECT -136.345 -269.040 -136.015 -268.750 ;
        RECT -114.750 -268.920 -69.490 -267.855 ;
        RECT -36.880 -268.565 -36.710 -265.605 ;
        RECT -34.765 -268.565 -34.595 -265.600 ;
        RECT -33.815 -265.615 -33.590 -264.985 ;
        RECT -33.165 -265.450 44.145 -264.985 ;
        RECT -33.785 -268.565 -33.615 -265.615 ;
        RECT -26.340 -265.985 -21.080 -265.450 ;
        RECT -26.340 -266.630 -26.140 -265.985 ;
        RECT -25.395 -266.630 -25.165 -265.985 ;
        RECT -24.405 -266.610 -24.175 -265.985 ;
        RECT -26.340 -267.545 -26.170 -266.630 ;
        RECT -25.360 -267.545 -25.190 -266.630 ;
        RECT -24.380 -267.545 -24.210 -266.610 ;
        RECT -23.840 -266.630 -23.610 -265.985 ;
        RECT -22.860 -266.605 -22.630 -265.985 ;
        RECT -23.810 -267.545 -23.640 -266.630 ;
        RECT -22.830 -267.545 -22.660 -266.605 ;
        RECT -22.295 -266.655 -22.065 -265.985 ;
        RECT -21.310 -266.595 -21.080 -265.985 ;
        RECT -22.265 -267.545 -22.095 -266.655 ;
        RECT -21.285 -267.545 -21.115 -266.595 ;
        RECT -114.750 -268.970 -103.575 -268.920 ;
        RECT -114.750 -269.040 -113.390 -268.970 ;
        RECT -136.345 -269.610 -113.390 -269.040 ;
        RECT -136.945 -269.670 -113.390 -269.610 ;
        RECT -139.180 -269.840 -113.390 -269.670 ;
        RECT -136.945 -269.905 -113.390 -269.840 ;
        RECT -136.945 -270.790 -136.705 -269.905 ;
        RECT -136.345 -270.400 -113.390 -269.905 ;
        RECT -136.345 -270.790 -136.015 -270.400 ;
        RECT -136.945 -270.850 -136.015 -270.790 ;
        RECT -139.180 -271.020 -136.015 -270.850 ;
        RECT -136.945 -271.085 -136.015 -271.020 ;
        RECT -136.945 -271.980 -136.705 -271.085 ;
        RECT -136.345 -271.980 -136.015 -271.085 ;
        RECT -136.945 -272.030 -136.015 -271.980 ;
        RECT -139.180 -272.200 -136.015 -272.030 ;
        RECT -136.945 -272.275 -136.015 -272.200 ;
        RECT -136.945 -273.180 -136.705 -272.275 ;
        RECT -136.345 -272.970 -136.015 -272.275 ;
        RECT -114.750 -272.970 -113.390 -270.400 ;
        RECT -106.685 -270.450 -106.515 -268.970 ;
        RECT -105.705 -270.450 -105.535 -268.970 ;
        RECT -104.725 -270.450 -104.555 -268.970 ;
        RECT -103.745 -270.450 -103.575 -268.970 ;
        RECT -101.060 -268.990 -99.835 -268.920 ;
        RECT -101.035 -270.450 -100.865 -268.990 ;
        RECT -100.055 -270.450 -99.885 -268.990 ;
        RECT -96.950 -269.230 -90.315 -268.920 ;
        RECT -96.950 -269.505 -90.295 -269.230 ;
        RECT -96.690 -271.560 -96.520 -269.505 ;
        RECT -95.710 -271.560 -95.540 -269.505 ;
        RECT -94.730 -269.725 -90.295 -269.505 ;
        RECT -94.730 -271.560 -94.560 -269.725 ;
        RECT -93.645 -270.555 -93.475 -269.725 ;
        RECT -92.665 -270.555 -92.495 -269.725 ;
        RECT -91.685 -270.555 -91.515 -269.725 ;
        RECT -90.705 -270.555 -90.535 -269.725 ;
        RECT -136.345 -273.180 -113.390 -272.970 ;
        RECT -136.945 -273.210 -113.390 -273.180 ;
        RECT -139.180 -273.380 -113.390 -273.210 ;
        RECT -136.945 -273.475 -113.390 -273.380 ;
        RECT -136.945 -274.330 -136.705 -273.475 ;
        RECT -136.345 -274.330 -113.390 -273.475 ;
        RECT -69.935 -273.535 -69.490 -268.920 ;
        RECT -19.705 -269.635 -19.130 -265.450 ;
        RECT -12.270 -265.640 -9.305 -265.450 ;
        RECT -13.840 -265.985 -8.580 -265.640 ;
        RECT -13.840 -266.630 -13.640 -265.985 ;
        RECT -12.895 -266.630 -12.665 -265.985 ;
        RECT -11.905 -266.610 -11.675 -265.985 ;
        RECT -13.840 -267.545 -13.670 -266.630 ;
        RECT -12.860 -267.545 -12.690 -266.630 ;
        RECT -11.880 -267.545 -11.710 -266.610 ;
        RECT -11.340 -266.630 -11.110 -265.985 ;
        RECT -10.360 -266.605 -10.130 -265.985 ;
        RECT -11.310 -267.545 -11.140 -266.630 ;
        RECT -10.330 -267.545 -10.160 -266.605 ;
        RECT -9.795 -266.655 -9.565 -265.985 ;
        RECT -8.810 -266.595 -8.580 -265.985 ;
        RECT -9.765 -267.545 -9.595 -266.655 ;
        RECT -8.785 -267.545 -8.615 -266.595 ;
        RECT -19.730 -270.315 -19.115 -269.635 ;
        RECT -6.865 -269.810 -6.295 -265.450 ;
        RECT 0.310 -265.640 3.275 -265.450 ;
        RECT -1.340 -265.985 3.920 -265.640 ;
        RECT -1.340 -266.630 -1.140 -265.985 ;
        RECT -0.395 -266.630 -0.165 -265.985 ;
        RECT 0.595 -266.610 0.825 -265.985 ;
        RECT -1.340 -267.545 -1.170 -266.630 ;
        RECT -0.360 -267.545 -0.190 -266.630 ;
        RECT 0.620 -267.545 0.790 -266.610 ;
        RECT 1.160 -266.630 1.390 -265.985 ;
        RECT 2.140 -266.605 2.370 -265.985 ;
        RECT 1.190 -267.545 1.360 -266.630 ;
        RECT 2.170 -267.545 2.340 -266.605 ;
        RECT 2.705 -266.655 2.935 -265.985 ;
        RECT 3.690 -266.595 3.920 -265.985 ;
        RECT 2.735 -267.545 2.905 -266.655 ;
        RECT 3.715 -267.545 3.885 -266.595 ;
        RECT 5.545 -269.810 6.120 -265.450 ;
        RECT 12.980 -265.640 15.945 -265.450 ;
        RECT 25.045 -265.640 28.010 -265.450 ;
        RECT 11.160 -265.985 16.420 -265.640 ;
        RECT 11.160 -266.630 11.360 -265.985 ;
        RECT 12.105 -266.630 12.335 -265.985 ;
        RECT 13.095 -266.610 13.325 -265.985 ;
        RECT 11.160 -267.545 11.330 -266.630 ;
        RECT 12.140 -267.545 12.310 -266.630 ;
        RECT 13.120 -267.545 13.290 -266.610 ;
        RECT 13.660 -266.630 13.890 -265.985 ;
        RECT 14.640 -266.605 14.870 -265.985 ;
        RECT 13.690 -267.545 13.860 -266.630 ;
        RECT 14.670 -267.545 14.840 -266.605 ;
        RECT 15.205 -266.655 15.435 -265.985 ;
        RECT 16.190 -266.595 16.420 -265.985 ;
        RECT 23.660 -265.985 28.920 -265.640 ;
        RECT 15.235 -267.545 15.405 -266.655 ;
        RECT 16.215 -267.545 16.385 -266.595 ;
        RECT 23.660 -266.630 23.860 -265.985 ;
        RECT 24.605 -266.630 24.835 -265.985 ;
        RECT 25.595 -266.610 25.825 -265.985 ;
        RECT 23.660 -267.545 23.830 -266.630 ;
        RECT 24.640 -267.545 24.810 -266.630 ;
        RECT 25.620 -267.545 25.790 -266.610 ;
        RECT 26.160 -266.630 26.390 -265.985 ;
        RECT 27.140 -266.605 27.370 -265.985 ;
        RECT 26.190 -267.545 26.360 -266.630 ;
        RECT 27.170 -267.545 27.340 -266.605 ;
        RECT 27.705 -266.655 27.935 -265.985 ;
        RECT 28.690 -266.595 28.920 -265.985 ;
        RECT 38.660 -265.985 43.920 -265.450 ;
        RECT 27.735 -267.545 27.905 -266.655 ;
        RECT 28.715 -267.545 28.885 -266.595 ;
        RECT 38.660 -266.630 38.860 -265.985 ;
        RECT 39.605 -266.630 39.835 -265.985 ;
        RECT 40.595 -266.610 40.825 -265.985 ;
        RECT 38.660 -267.545 38.830 -266.630 ;
        RECT 39.640 -267.545 39.810 -266.630 ;
        RECT 40.620 -267.545 40.790 -266.610 ;
        RECT 41.160 -266.630 41.390 -265.985 ;
        RECT 42.140 -266.605 42.370 -265.985 ;
        RECT 41.190 -267.545 41.360 -266.630 ;
        RECT 42.170 -267.545 42.340 -266.605 ;
        RECT 42.705 -266.655 42.935 -265.985 ;
        RECT 43.690 -266.595 43.920 -265.985 ;
        RECT 133.130 -266.260 138.645 -259.315 ;
        RECT 42.735 -267.545 42.905 -266.655 ;
        RECT 43.715 -267.545 43.885 -266.595 ;
        RECT -6.895 -270.490 -6.280 -269.810 ;
        RECT 5.520 -270.490 6.135 -269.810 ;
        RECT -68.200 -273.520 -68.030 -272.065 ;
        RECT -67.220 -273.520 -67.050 -272.065 ;
        RECT -66.240 -273.520 -66.070 -272.065 ;
        RECT -59.485 -273.520 -59.315 -272.065 ;
        RECT -58.505 -273.520 -58.335 -272.065 ;
        RECT -57.525 -273.520 -57.355 -272.065 ;
        RECT -54.700 -273.520 -54.530 -272.065 ;
        RECT -53.720 -273.520 -53.550 -272.065 ;
        RECT -52.740 -273.520 -52.570 -272.065 ;
        RECT -45.985 -273.520 -45.815 -272.065 ;
        RECT -45.005 -273.520 -44.835 -272.065 ;
        RECT -44.025 -273.520 -43.855 -272.065 ;
        RECT -41.575 -273.520 -41.405 -272.065 ;
        RECT -40.595 -273.520 -40.425 -272.065 ;
        RECT -39.615 -273.520 -39.445 -272.065 ;
        RECT 5.515 -272.580 6.130 -272.575 ;
        RECT -68.500 -273.535 -66.025 -273.520 ;
        RECT -59.790 -273.525 -52.525 -273.520 ;
        RECT -69.935 -273.545 -64.415 -273.535 ;
        RECT -59.790 -273.545 -50.960 -273.525 ;
        RECT -46.290 -273.545 -39.400 -273.520 ;
        RECT -136.945 -274.390 -136.015 -274.330 ;
        RECT -139.180 -274.560 -136.015 -274.390 ;
        RECT -136.945 -274.625 -136.015 -274.560 ;
        RECT -136.945 -275.515 -136.705 -274.625 ;
        RECT -136.345 -275.515 -136.015 -274.625 ;
        RECT -136.945 -275.570 -136.015 -275.515 ;
        RECT -139.180 -275.740 -136.015 -275.570 ;
        RECT -136.945 -275.810 -136.015 -275.740 ;
        RECT -136.945 -276.685 -136.705 -275.810 ;
        RECT -136.345 -276.640 -136.015 -275.810 ;
        RECT -114.750 -276.640 -113.390 -274.330 ;
        RECT -136.345 -276.685 -113.390 -276.640 ;
        RECT -136.945 -276.750 -113.390 -276.685 ;
        RECT -139.180 -276.920 -113.390 -276.750 ;
        RECT -88.510 -276.915 -88.340 -274.830 ;
        RECT -87.530 -276.915 -87.360 -274.830 ;
        RECT -86.550 -276.665 -86.380 -274.830 ;
        RECT -85.465 -276.665 -85.295 -275.835 ;
        RECT -84.485 -276.665 -84.315 -275.835 ;
        RECT -83.505 -276.665 -83.335 -275.835 ;
        RECT -82.525 -276.665 -82.355 -275.835 ;
        RECT -86.550 -276.915 -82.115 -276.665 ;
        RECT -81.275 -276.725 -81.105 -273.775 ;
        RECT -136.945 -276.980 -113.390 -276.920 ;
        RECT -136.945 -277.855 -136.705 -276.980 ;
        RECT -136.345 -277.675 -113.390 -276.980 ;
        RECT -88.560 -277.160 -82.115 -276.915 ;
        RECT -88.560 -277.235 -86.350 -277.160 ;
        RECT -81.300 -277.355 -81.075 -276.725 ;
        RECT -80.295 -276.740 -80.125 -273.775 ;
        RECT -78.180 -276.735 -78.010 -273.775 ;
        RECT -69.935 -273.860 -39.400 -273.545 ;
        RECT -69.935 -273.875 -64.415 -273.860 ;
        RECT -53.325 -273.865 -50.960 -273.860 ;
        RECT -80.325 -277.355 -80.100 -276.740 ;
        RECT -78.215 -277.355 -77.990 -276.735 ;
        RECT -86.365 -277.440 -85.420 -277.405 ;
        RECT -86.550 -277.475 -85.420 -277.440 ;
        RECT -81.330 -277.475 -77.485 -277.355 ;
        RECT -88.560 -277.675 -77.485 -277.475 ;
        RECT -136.345 -277.685 -77.485 -277.675 ;
        RECT -136.345 -277.855 -78.005 -277.685 ;
        RECT -136.945 -277.930 -78.005 -277.855 ;
        RECT -139.180 -278.000 -78.005 -277.930 ;
        RECT -139.180 -278.100 -136.015 -278.000 ;
        RECT -136.945 -278.150 -136.015 -278.100 ;
        RECT -136.945 -279.110 -136.705 -278.150 ;
        RECT -139.180 -279.280 -136.705 -279.110 ;
        RECT -136.945 -280.350 -136.705 -279.280 ;
        RECT -139.180 -280.520 -136.705 -280.350 ;
        RECT -136.945 -281.480 -136.705 -280.520 ;
        RECT -136.345 -281.480 -136.015 -278.150 ;
        RECT -114.750 -278.240 -78.005 -278.000 ;
        RECT -114.750 -278.670 -90.685 -278.240 ;
        RECT -114.750 -278.835 -90.735 -278.670 ;
        RECT -106.450 -279.020 -100.005 -278.835 ;
        RECT -106.400 -281.105 -106.230 -279.020 ;
        RECT -105.420 -281.105 -105.250 -279.020 ;
        RECT -104.440 -279.270 -100.005 -279.020 ;
        RECT -104.440 -281.105 -104.270 -279.270 ;
        RECT -103.355 -280.100 -103.185 -279.270 ;
        RECT -102.375 -280.100 -102.205 -279.270 ;
        RECT -101.395 -280.100 -101.225 -279.270 ;
        RECT -100.415 -280.100 -100.245 -279.270 ;
        RECT -97.535 -280.130 -97.365 -278.835 ;
        RECT -96.555 -280.130 -96.385 -278.835 ;
        RECT -95.575 -280.130 -95.405 -278.835 ;
        RECT -94.595 -280.130 -94.425 -278.835 ;
        RECT -91.885 -280.130 -91.715 -278.835 ;
        RECT -90.905 -280.130 -90.735 -278.835 ;
        RECT -87.710 -279.190 -86.850 -278.240 ;
        RECT -83.570 -278.325 -80.480 -278.240 ;
        RECT -83.570 -278.470 -81.355 -278.325 ;
        RECT -83.565 -278.540 -81.355 -278.470 ;
        RECT -83.565 -278.785 -77.120 -278.540 ;
        RECT -88.620 -279.685 -85.030 -279.190 ;
        RECT -88.380 -281.015 -88.210 -279.685 ;
        RECT -87.400 -281.015 -87.230 -279.685 ;
        RECT -86.420 -281.015 -86.250 -279.685 ;
        RECT -85.440 -281.015 -85.270 -279.685 ;
        RECT -83.515 -280.870 -83.345 -278.785 ;
        RECT -82.535 -280.870 -82.365 -278.785 ;
        RECT -81.555 -279.035 -77.120 -278.785 ;
        RECT -81.555 -280.870 -81.385 -279.035 ;
        RECT -80.470 -279.865 -80.300 -279.035 ;
        RECT -79.490 -279.865 -79.320 -279.035 ;
        RECT -78.510 -279.865 -78.340 -279.035 ;
        RECT -77.530 -279.865 -77.360 -279.035 ;
        RECT -136.945 -281.530 -136.015 -281.480 ;
        RECT -139.180 -281.700 -136.015 -281.530 ;
        RECT -136.945 -281.775 -136.015 -281.700 ;
        RECT -136.945 -282.635 -136.705 -281.775 ;
        RECT -136.345 -282.635 -136.015 -281.775 ;
        RECT -136.945 -282.710 -136.015 -282.635 ;
        RECT -139.180 -282.880 -136.015 -282.710 ;
        RECT -136.945 -282.930 -136.015 -282.880 ;
        RECT -136.945 -283.815 -136.705 -282.930 ;
        RECT -136.345 -283.815 -136.015 -282.930 ;
        RECT -136.945 -283.890 -136.015 -283.815 ;
        RECT -139.180 -284.060 -136.015 -283.890 ;
        RECT -136.945 -284.110 -136.015 -284.060 ;
        RECT -136.945 -284.990 -136.705 -284.110 ;
        RECT -136.345 -284.990 -136.015 -284.110 ;
        RECT -136.945 -285.070 -136.015 -284.990 ;
        RECT -139.180 -285.240 -136.015 -285.070 ;
        RECT -136.945 -285.285 -136.015 -285.240 ;
        RECT -136.945 -286.185 -136.705 -285.285 ;
        RECT -136.345 -286.185 -136.015 -285.285 ;
        RECT -136.945 -286.250 -136.015 -286.185 ;
        RECT -139.180 -286.420 -136.015 -286.250 ;
        RECT -136.945 -286.480 -136.015 -286.420 ;
        RECT -136.945 -287.330 -136.705 -286.480 ;
        RECT -136.345 -287.330 -136.015 -286.480 ;
        RECT -136.945 -287.430 -136.015 -287.330 ;
        RECT -139.180 -287.600 -136.015 -287.430 ;
        RECT -136.945 -287.625 -136.015 -287.600 ;
        RECT -136.945 -288.610 -136.705 -287.625 ;
        RECT -139.180 -288.780 -136.705 -288.610 ;
        RECT -136.945 -289.790 -136.705 -288.780 ;
        RECT -139.180 -289.960 -136.705 -289.790 ;
        RECT -136.945 -290.360 -136.705 -289.960 ;
        RECT -136.345 -290.360 -136.015 -287.625 ;
        RECT -67.625 -282.355 -66.860 -273.875 ;
        RECT -28.035 -274.605 -27.865 -273.150 ;
        RECT -27.055 -274.605 -26.885 -273.150 ;
        RECT -26.075 -274.605 -25.905 -273.150 ;
        RECT -6.900 -273.430 -6.285 -272.750 ;
        RECT 5.515 -272.890 7.045 -272.580 ;
        RECT -19.735 -274.150 -19.120 -273.470 ;
        RECT -28.080 -274.945 -25.605 -274.605 ;
        RECT -28.000 -276.895 -27.560 -274.945 ;
        RECT -27.085 -276.895 -26.645 -274.945 ;
        RECT -26.175 -276.895 -25.735 -274.945 ;
        RECT -30.565 -276.910 -25.045 -276.895 ;
        RECT -19.710 -276.910 -19.135 -274.150 ;
        RECT -13.955 -276.910 -11.590 -276.905 ;
        RECT -6.880 -276.910 -6.305 -273.430 ;
        RECT -0.605 -276.910 0.010 -276.800 ;
        RECT -30.565 -277.225 0.010 -276.910 ;
        RECT -30.565 -277.235 -25.045 -277.225 ;
        RECT -63.565 -281.795 -63.395 -279.710 ;
        RECT -62.585 -281.795 -62.415 -279.710 ;
        RECT -61.605 -281.545 -61.435 -279.710 ;
        RECT -60.520 -281.545 -60.350 -280.715 ;
        RECT -59.540 -281.545 -59.370 -280.715 ;
        RECT -58.560 -281.545 -58.390 -280.715 ;
        RECT -57.580 -281.545 -57.410 -280.715 ;
        RECT -61.605 -281.795 -57.170 -281.545 ;
        RECT -56.330 -281.605 -56.160 -278.655 ;
        RECT -63.615 -282.040 -57.170 -281.795 ;
        RECT -63.615 -282.115 -61.405 -282.040 ;
        RECT -56.355 -282.235 -56.130 -281.605 ;
        RECT -55.350 -281.620 -55.180 -278.655 ;
        RECT -53.235 -281.615 -53.065 -278.655 ;
        RECT -55.380 -282.235 -55.155 -281.620 ;
        RECT -53.270 -282.235 -53.045 -281.615 ;
        RECT -61.420 -282.320 -60.475 -282.285 ;
        RECT -61.605 -282.355 -60.475 -282.320 ;
        RECT -56.385 -282.355 -52.540 -282.235 ;
        RECT -67.625 -282.565 -52.540 -282.355 ;
        RECT -67.625 -283.120 -53.060 -282.565 ;
        RECT -67.625 -289.355 -66.860 -283.120 ;
        RECT -62.765 -284.070 -61.905 -283.120 ;
        RECT -58.625 -283.205 -55.535 -283.120 ;
        RECT -58.625 -283.350 -56.410 -283.205 ;
        RECT -58.620 -283.420 -56.410 -283.350 ;
        RECT -58.620 -283.665 -52.175 -283.420 ;
        RECT -63.675 -284.565 -60.085 -284.070 ;
        RECT -63.435 -285.895 -63.265 -284.565 ;
        RECT -62.455 -285.895 -62.285 -284.565 ;
        RECT -61.475 -285.895 -61.305 -284.565 ;
        RECT -60.495 -285.895 -60.325 -284.565 ;
        RECT -58.570 -285.750 -58.400 -283.665 ;
        RECT -57.590 -285.750 -57.420 -283.665 ;
        RECT -56.610 -283.915 -52.175 -283.665 ;
        RECT -56.610 -285.750 -56.440 -283.915 ;
        RECT -55.525 -284.745 -55.355 -283.915 ;
        RECT -54.545 -284.745 -54.375 -283.915 ;
        RECT -53.565 -284.745 -53.395 -283.915 ;
        RECT -52.585 -284.745 -52.415 -283.915 ;
        RECT -30.565 -285.710 -30.120 -277.235 ;
        RECT -29.130 -277.250 -26.655 -277.235 ;
        RECT -20.420 -277.245 -11.590 -277.225 ;
        RECT -20.420 -277.250 -13.155 -277.245 ;
        RECT -6.920 -277.250 0.010 -277.225 ;
        RECT -28.830 -278.705 -28.660 -277.250 ;
        RECT -27.850 -278.705 -27.680 -277.250 ;
        RECT -26.870 -278.705 -26.700 -277.250 ;
        RECT -20.115 -278.705 -19.945 -277.250 ;
        RECT -19.135 -278.705 -18.965 -277.250 ;
        RECT -18.155 -278.705 -17.985 -277.250 ;
        RECT -15.330 -278.705 -15.160 -277.250 ;
        RECT -14.350 -278.705 -14.180 -277.250 ;
        RECT -13.370 -278.705 -13.200 -277.250 ;
        RECT -6.615 -278.705 -6.445 -277.250 ;
        RECT -5.635 -278.705 -5.465 -277.250 ;
        RECT -4.655 -278.705 -4.485 -277.250 ;
        RECT -2.205 -278.705 -2.035 -277.250 ;
        RECT -1.225 -278.705 -1.055 -277.250 ;
        RECT -0.605 -277.480 0.010 -277.250 ;
        RECT 0.865 -276.930 1.480 -276.795 ;
        RECT 5.540 -276.930 6.115 -272.890 ;
        RECT 15.755 -276.930 16.370 -276.860 ;
        RECT 0.865 -277.325 16.370 -276.930 ;
        RECT 0.865 -277.330 2.640 -277.325 ;
        RECT 0.865 -277.475 1.635 -277.330 ;
        RECT -0.245 -278.705 -0.075 -277.480 ;
        RECT 1.465 -278.790 1.635 -277.475 ;
        RECT 2.445 -278.790 2.615 -277.330 ;
        RECT 5.155 -278.790 5.325 -277.325 ;
        RECT 6.135 -278.790 6.305 -277.325 ;
        RECT 7.115 -278.790 7.285 -277.325 ;
        RECT 8.095 -278.790 8.265 -277.325 ;
        RECT 9.890 -277.525 14.325 -277.325 ;
        RECT 10.130 -278.355 10.300 -277.525 ;
        RECT 11.110 -278.355 11.280 -277.525 ;
        RECT 12.090 -278.355 12.260 -277.525 ;
        RECT 13.070 -278.355 13.240 -277.525 ;
        RECT 14.155 -279.360 14.325 -277.525 ;
        RECT 15.135 -279.360 15.305 -277.325 ;
        RECT 15.755 -277.540 16.370 -277.325 ;
        RECT 17.700 -277.040 18.315 -276.855 ;
        RECT 23.840 -276.965 24.455 -276.740 ;
        RECT 22.150 -277.040 24.455 -276.965 ;
        RECT 17.700 -277.285 24.455 -277.040 ;
        RECT 17.700 -277.535 22.350 -277.285 ;
        RECT 16.115 -279.360 16.285 -277.540 ;
        RECT 18.155 -278.365 18.325 -277.535 ;
        RECT 19.135 -278.365 19.305 -277.535 ;
        RECT 20.115 -278.365 20.285 -277.535 ;
        RECT 21.095 -278.365 21.265 -277.535 ;
        RECT 22.180 -279.370 22.350 -277.535 ;
        RECT 23.160 -279.370 23.330 -277.285 ;
        RECT 23.840 -277.420 24.455 -277.285 ;
        RECT 25.845 -276.895 26.460 -276.730 ;
        RECT 25.845 -276.920 30.325 -276.895 ;
        RECT 32.625 -276.920 33.240 -276.755 ;
        RECT 25.845 -277.260 33.240 -276.920 ;
        RECT 25.845 -277.285 27.450 -277.260 ;
        RECT 29.965 -277.265 33.240 -277.260 ;
        RECT 25.845 -277.410 26.460 -277.285 ;
        RECT 24.140 -279.370 24.310 -277.420 ;
        RECT 26.275 -278.745 26.445 -277.410 ;
        RECT 27.255 -278.745 27.425 -277.285 ;
        RECT 29.965 -278.745 30.135 -277.265 ;
        RECT 30.945 -278.745 31.115 -277.265 ;
        RECT 31.925 -278.745 32.095 -277.265 ;
        RECT 32.625 -277.435 33.240 -277.265 ;
        RECT 38.705 -276.895 39.320 -276.760 ;
        RECT 38.705 -277.240 43.970 -276.895 ;
        RECT 32.905 -278.745 33.075 -277.435 ;
        RECT 38.705 -277.440 39.320 -277.240 ;
        RECT 38.710 -277.885 38.910 -277.440 ;
        RECT 39.655 -277.885 39.885 -277.240 ;
        RECT 40.645 -277.865 40.875 -277.240 ;
        RECT 38.710 -278.800 38.880 -277.885 ;
        RECT 39.690 -278.800 39.860 -277.885 ;
        RECT 40.670 -278.800 40.840 -277.865 ;
        RECT 41.210 -277.885 41.440 -277.240 ;
        RECT 42.190 -277.860 42.420 -277.240 ;
        RECT 41.240 -278.800 41.410 -277.885 ;
        RECT 42.220 -278.800 42.390 -277.860 ;
        RECT 42.755 -277.910 42.985 -277.240 ;
        RECT 43.740 -277.850 43.970 -277.240 ;
        RECT 42.785 -278.800 42.955 -277.910 ;
        RECT 43.765 -278.800 43.935 -277.850 ;
        RECT 104.870 -278.570 130.995 -278.255 ;
        RECT 109.630 -278.595 118.640 -278.570 ;
        RECT 123.130 -278.595 130.995 -278.570 ;
        RECT 141.795 -278.575 141.965 -277.245 ;
        RECT 142.775 -278.575 142.945 -277.245 ;
        RECT 143.755 -278.575 143.925 -277.245 ;
        RECT 144.735 -278.575 144.905 -277.245 ;
        RECT 109.935 -280.050 110.105 -278.595 ;
        RECT 110.915 -280.050 111.085 -278.595 ;
        RECT 111.895 -280.050 112.065 -278.595 ;
        RECT 114.120 -280.050 114.290 -278.595 ;
        RECT 115.100 -280.050 115.270 -278.595 ;
        RECT 116.080 -280.050 116.250 -278.595 ;
        RECT 123.435 -280.050 123.605 -278.595 ;
        RECT 124.415 -280.050 124.585 -278.595 ;
        RECT 125.395 -280.050 125.565 -278.595 ;
        RECT 127.620 -280.050 127.790 -278.595 ;
        RECT 128.600 -280.050 128.770 -278.595 ;
        RECT 129.580 -280.050 129.750 -278.595 ;
        RECT 130.550 -278.895 130.995 -278.595 ;
        RECT 141.555 -278.895 145.145 -278.575 ;
        RECT 130.550 -279.070 145.145 -278.895 ;
        RECT 130.550 -280.020 143.325 -279.070 ;
        RECT 146.660 -279.475 146.830 -277.390 ;
        RECT 147.640 -279.475 147.810 -277.390 ;
        RECT 148.620 -279.225 148.790 -277.390 ;
        RECT 149.705 -279.225 149.875 -278.395 ;
        RECT 150.685 -279.225 150.855 -278.395 ;
        RECT 151.665 -279.225 151.835 -278.395 ;
        RECT 152.645 -279.225 152.815 -278.395 ;
        RECT 183.995 -278.630 184.165 -277.300 ;
        RECT 184.975 -278.630 185.145 -277.300 ;
        RECT 185.955 -278.630 186.125 -277.300 ;
        RECT 186.935 -278.630 187.105 -277.300 ;
        RECT 183.755 -279.125 187.345 -278.630 ;
        RECT 148.620 -279.475 153.055 -279.225 ;
        RECT 146.610 -279.720 153.055 -279.475 ;
        RECT 146.610 -279.790 148.820 -279.720 ;
        RECT 158.845 -279.750 171.005 -279.400 ;
        RECT 146.605 -279.935 148.820 -279.790 ;
        RECT 146.605 -280.020 149.695 -279.935 ;
        RECT 157.010 -280.010 171.005 -279.750 ;
        RECT 157.010 -280.015 165.775 -280.010 ;
        RECT 130.550 -280.365 152.170 -280.020 ;
        RECT -29.320 -285.710 -29.150 -284.255 ;
        RECT -28.340 -285.710 -28.170 -284.255 ;
        RECT -27.360 -285.710 -27.190 -284.255 ;
        RECT -25.135 -285.710 -24.965 -284.255 ;
        RECT -24.155 -285.710 -23.985 -284.255 ;
        RECT -23.175 -285.710 -23.005 -284.255 ;
        RECT -15.820 -285.710 -15.650 -284.255 ;
        RECT -14.840 -285.710 -14.670 -284.255 ;
        RECT -13.860 -285.710 -13.690 -284.255 ;
        RECT -11.635 -285.710 -11.465 -284.255 ;
        RECT -10.655 -285.710 -10.485 -284.255 ;
        RECT -9.675 -285.710 -9.505 -284.255 ;
        RECT -30.565 -285.735 -22.700 -285.710 ;
        RECT -18.210 -285.735 -9.200 -285.710 ;
        RECT -30.565 -286.050 -4.440 -285.735 ;
        RECT 93.900 -286.000 94.070 -283.000 ;
        RECT 94.880 -285.920 95.050 -283.000 ;
        RECT -30.565 -289.245 -30.120 -286.050 ;
        RECT -49.545 -289.355 -30.120 -289.245 ;
        RECT -136.945 -290.440 -136.015 -290.360 ;
        RECT -139.180 -290.610 -136.015 -290.440 ;
        RECT -136.945 -290.655 -136.015 -290.610 ;
        RECT -136.945 -291.520 -136.705 -290.655 ;
        RECT -136.345 -291.520 -136.015 -290.655 ;
        RECT -136.945 -291.620 -136.015 -291.520 ;
        RECT -139.180 -291.790 -136.015 -291.620 ;
        RECT -136.945 -291.815 -136.015 -291.790 ;
        RECT -136.945 -292.725 -136.705 -291.815 ;
        RECT -136.345 -292.725 -136.015 -291.815 ;
        RECT -136.945 -292.800 -136.015 -292.725 ;
        RECT -139.180 -292.970 -136.015 -292.800 ;
        RECT -69.935 -289.670 -30.120 -289.355 ;
        RECT -69.935 -289.695 -62.070 -289.670 ;
        RECT -57.580 -289.695 -48.570 -289.670 ;
        RECT -69.935 -292.820 -69.490 -289.695 ;
        RECT -68.690 -291.150 -68.520 -289.695 ;
        RECT -67.710 -291.150 -67.540 -289.695 ;
        RECT -66.730 -291.150 -66.560 -289.695 ;
        RECT -64.505 -291.150 -64.335 -289.695 ;
        RECT -63.525 -291.150 -63.355 -289.695 ;
        RECT -62.545 -291.150 -62.375 -289.695 ;
        RECT -55.190 -291.150 -55.020 -289.695 ;
        RECT -54.210 -291.150 -54.040 -289.695 ;
        RECT -53.230 -291.150 -53.060 -289.695 ;
        RECT -51.005 -291.150 -50.835 -289.695 ;
        RECT -50.025 -291.150 -49.855 -289.695 ;
        RECT -49.045 -291.150 -48.875 -289.695 ;
        RECT -36.765 -290.275 -36.540 -289.670 ;
        RECT -34.655 -290.270 -34.430 -289.670 ;
        RECT -136.945 -293.020 -136.015 -292.970 ;
        RECT -136.945 -293.980 -136.705 -293.020 ;
        RECT -139.180 -294.080 -136.705 -293.980 ;
        RECT -136.345 -294.080 -136.015 -293.020 ;
        RECT -107.670 -293.655 -69.485 -292.820 ;
        RECT -36.745 -293.235 -36.575 -290.275 ;
        RECT -34.630 -293.235 -34.460 -290.270 ;
        RECT -33.680 -290.285 -33.455 -289.670 ;
        RECT -30.565 -290.245 -30.120 -289.670 ;
        RECT -33.650 -293.235 -33.480 -290.285 ;
        RECT -30.565 -290.690 -30.115 -290.245 ;
        RECT -29.125 -290.690 -27.780 -286.050 ;
        RECT -26.395 -290.690 -25.050 -286.050 ;
        RECT -22.010 -290.690 -20.665 -286.050 ;
        RECT -17.700 -290.690 -16.355 -286.050 ;
        RECT -13.185 -290.690 -11.840 -286.050 ;
        RECT -8.030 -290.690 -6.685 -286.050 ;
        RECT 93.855 -286.560 94.120 -286.000 ;
        RECT 94.835 -286.560 95.100 -285.920 ;
        RECT 93.855 -287.225 98.195 -286.560 ;
        RECT 100.505 -287.055 100.675 -285.600 ;
        RECT 101.485 -287.055 101.655 -285.600 ;
        RECT 102.465 -287.055 102.635 -285.600 ;
        RECT 104.915 -287.055 105.085 -285.600 ;
        RECT 105.895 -287.055 106.065 -285.600 ;
        RECT 106.875 -287.055 107.045 -285.600 ;
        RECT 113.630 -287.055 113.800 -285.600 ;
        RECT 114.610 -287.055 114.780 -285.600 ;
        RECT 115.590 -287.055 115.760 -285.600 ;
        RECT 118.415 -287.055 118.585 -285.600 ;
        RECT 119.395 -287.055 119.565 -285.600 ;
        RECT 120.375 -287.055 120.545 -285.600 ;
        RECT 127.130 -287.055 127.300 -285.600 ;
        RECT 128.110 -287.055 128.280 -285.600 ;
        RECT 129.090 -287.055 129.260 -285.600 ;
        RECT 100.460 -287.080 107.350 -287.055 ;
        RECT 113.585 -287.060 120.850 -287.055 ;
        RECT 112.020 -287.080 120.850 -287.060 ;
        RECT 127.085 -287.070 129.560 -287.055 ;
        RECT 130.550 -287.070 130.995 -280.365 ;
        RECT 141.615 -280.575 152.170 -280.365 ;
        RECT 157.010 -280.335 159.035 -280.015 ;
        RECT 154.195 -280.385 154.685 -280.370 ;
        RECT 157.010 -280.385 157.595 -280.335 ;
        RECT 141.615 -280.610 152.690 -280.575 ;
        RECT 153.055 -280.610 153.365 -280.470 ;
        RECT 141.615 -280.785 153.365 -280.610 ;
        RECT 143.625 -280.820 144.755 -280.785 ;
        RECT 143.810 -280.855 144.755 -280.820 ;
        RECT 148.845 -280.870 153.365 -280.785 ;
        RECT 148.845 -280.905 152.690 -280.870 ;
        RECT 141.615 -281.100 143.825 -281.025 ;
        RECT 141.615 -281.345 148.060 -281.100 ;
        RECT 141.665 -283.430 141.835 -281.345 ;
        RECT 142.645 -283.430 142.815 -281.345 ;
        RECT 143.625 -281.595 148.060 -281.345 ;
        RECT 148.875 -281.535 149.100 -280.905 ;
        RECT 149.850 -281.520 150.075 -280.905 ;
        RECT 143.625 -283.430 143.795 -281.595 ;
        RECT 144.710 -282.425 144.880 -281.595 ;
        RECT 145.690 -282.425 145.860 -281.595 ;
        RECT 146.670 -282.425 146.840 -281.595 ;
        RECT 147.650 -282.425 147.820 -281.595 ;
        RECT 148.900 -284.485 149.070 -281.535 ;
        RECT 149.880 -284.485 150.050 -281.520 ;
        RECT 151.960 -281.525 152.185 -280.905 ;
        RECT 153.055 -280.940 153.365 -280.870 ;
        RECT 154.195 -280.970 157.595 -280.385 ;
        RECT 158.845 -280.810 159.035 -280.335 ;
        RECT 159.830 -280.800 160.020 -280.015 ;
        RECT 154.195 -281.000 154.685 -280.970 ;
        RECT 151.995 -284.485 152.165 -281.525 ;
        RECT 158.860 -283.275 159.030 -280.810 ;
        RECT 159.840 -283.275 160.010 -280.800 ;
        RECT 162.790 -280.915 163.040 -280.015 ;
        RECT 163.420 -280.900 163.670 -280.015 ;
        RECT 164.575 -280.825 164.790 -280.015 ;
        RECT 165.560 -280.815 165.775 -280.015 ;
        RECT 170.395 -280.075 171.005 -280.010 ;
        RECT 184.665 -280.075 185.525 -279.125 ;
        RECT 188.860 -279.530 189.030 -277.445 ;
        RECT 189.840 -279.530 190.010 -277.445 ;
        RECT 190.820 -279.280 190.990 -277.445 ;
        RECT 191.905 -279.280 192.075 -278.450 ;
        RECT 192.885 -279.280 193.055 -278.450 ;
        RECT 193.865 -279.280 194.035 -278.450 ;
        RECT 194.845 -279.280 195.015 -278.450 ;
        RECT 228.310 -278.825 228.480 -277.495 ;
        RECT 229.290 -278.825 229.460 -277.495 ;
        RECT 230.270 -278.825 230.440 -277.495 ;
        RECT 231.250 -278.825 231.420 -277.495 ;
        RECT 228.070 -279.245 231.660 -278.825 ;
        RECT 190.820 -279.530 195.255 -279.280 ;
        RECT 207.905 -279.320 231.660 -279.245 ;
        RECT 207.905 -279.455 229.840 -279.320 ;
        RECT 188.810 -279.775 195.255 -279.530 ;
        RECT 188.810 -279.845 191.020 -279.775 ;
        RECT 201.045 -279.805 229.840 -279.455 ;
        RECT 233.175 -279.725 233.345 -277.640 ;
        RECT 234.155 -279.725 234.325 -277.640 ;
        RECT 235.135 -279.475 235.305 -277.640 ;
        RECT 236.220 -279.475 236.390 -278.645 ;
        RECT 237.200 -279.475 237.370 -278.645 ;
        RECT 238.180 -279.475 238.350 -278.645 ;
        RECT 239.160 -279.475 239.330 -278.645 ;
        RECT 274.300 -278.655 274.470 -277.325 ;
        RECT 275.280 -278.655 275.450 -277.325 ;
        RECT 276.260 -278.655 276.430 -277.325 ;
        RECT 277.240 -278.655 277.410 -277.325 ;
        RECT 274.060 -278.995 277.650 -278.655 ;
        RECT 252.160 -279.150 277.650 -278.995 ;
        RECT 235.135 -279.725 239.570 -279.475 ;
        RECT 252.160 -279.650 275.830 -279.150 ;
        RECT 279.165 -279.555 279.335 -277.470 ;
        RECT 280.145 -279.555 280.315 -277.470 ;
        RECT 281.125 -279.305 281.295 -277.470 ;
        RECT 318.070 -278.325 318.240 -276.995 ;
        RECT 319.050 -278.325 319.220 -276.995 ;
        RECT 320.030 -278.325 320.200 -276.995 ;
        RECT 321.010 -278.325 321.180 -276.995 ;
        RECT 282.210 -279.305 282.380 -278.475 ;
        RECT 283.190 -279.305 283.360 -278.475 ;
        RECT 284.170 -279.305 284.340 -278.475 ;
        RECT 285.150 -279.305 285.320 -278.475 ;
        RECT 317.830 -278.510 321.420 -278.325 ;
        RECT 298.075 -278.820 321.420 -278.510 ;
        RECT 281.125 -279.555 285.560 -279.305 ;
        RECT 298.075 -279.480 319.600 -278.820 ;
        RECT 322.935 -279.225 323.105 -277.140 ;
        RECT 323.915 -279.225 324.085 -277.140 ;
        RECT 324.895 -278.975 325.065 -277.140 ;
        RECT 325.980 -278.975 326.150 -278.145 ;
        RECT 326.960 -278.975 327.130 -278.145 ;
        RECT 327.940 -278.975 328.110 -278.145 ;
        RECT 328.920 -278.975 329.090 -278.145 ;
        RECT 363.835 -278.240 364.005 -276.910 ;
        RECT 364.815 -278.240 364.985 -276.910 ;
        RECT 365.795 -278.240 365.965 -276.910 ;
        RECT 366.775 -278.240 366.945 -276.910 ;
        RECT 363.595 -278.615 367.185 -278.240 ;
        RECT 341.810 -278.735 367.185 -278.615 ;
        RECT 324.895 -279.225 329.330 -278.975 ;
        RECT 341.810 -279.150 365.365 -278.735 ;
        RECT 368.700 -279.140 368.870 -277.055 ;
        RECT 369.680 -279.140 369.850 -277.055 ;
        RECT 370.660 -278.890 370.830 -277.055 ;
        RECT 410.655 -278.050 410.825 -276.720 ;
        RECT 411.635 -278.050 411.805 -276.720 ;
        RECT 412.615 -278.050 412.785 -276.720 ;
        RECT 413.595 -278.050 413.765 -276.720 ;
        RECT 371.745 -278.890 371.915 -278.060 ;
        RECT 372.725 -278.890 372.895 -278.060 ;
        RECT 373.705 -278.890 373.875 -278.060 ;
        RECT 374.685 -278.890 374.855 -278.060 ;
        RECT 410.415 -278.270 414.005 -278.050 ;
        RECT 387.620 -278.545 414.005 -278.270 ;
        RECT 370.660 -279.140 375.095 -278.890 ;
        RECT 387.620 -279.065 412.185 -278.545 ;
        RECT 415.520 -278.950 415.690 -276.865 ;
        RECT 416.500 -278.950 416.670 -276.865 ;
        RECT 417.480 -278.700 417.650 -276.865 ;
        RECT 418.565 -278.700 418.735 -277.870 ;
        RECT 419.545 -278.700 419.715 -277.870 ;
        RECT 420.525 -278.700 420.695 -277.870 ;
        RECT 421.505 -278.700 421.675 -277.870 ;
        RECT 417.480 -278.950 421.915 -278.700 ;
        RECT 436.495 -278.875 438.870 -259.315 ;
        RECT 188.805 -279.990 191.020 -279.845 ;
        RECT 188.805 -280.075 191.895 -279.990 ;
        RECT 199.210 -280.070 229.840 -279.805 ;
        RECT 233.125 -279.970 239.570 -279.725 ;
        RECT 233.125 -280.040 235.335 -279.970 ;
        RECT 245.360 -280.000 275.830 -279.650 ;
        RECT 279.115 -279.800 285.560 -279.555 ;
        RECT 291.350 -279.770 319.600 -279.480 ;
        RECT 322.885 -279.470 329.330 -279.225 ;
        RECT 322.885 -279.540 325.095 -279.470 ;
        RECT 335.120 -279.500 365.365 -279.150 ;
        RECT 368.650 -279.385 375.095 -279.140 ;
        RECT 368.650 -279.455 370.860 -279.385 ;
        RECT 380.885 -279.415 412.185 -279.065 ;
        RECT 415.470 -279.195 421.915 -278.950 ;
        RECT 415.470 -279.265 417.680 -279.195 ;
        RECT 427.705 -279.225 439.865 -278.875 ;
        RECT 322.880 -279.685 325.095 -279.540 ;
        RECT 333.285 -279.685 365.365 -279.500 ;
        RECT 368.645 -279.600 370.860 -279.455 ;
        RECT 379.050 -279.495 412.185 -279.415 ;
        RECT 415.465 -279.410 417.680 -279.265 ;
        RECT 415.465 -279.495 418.555 -279.410 ;
        RECT 425.870 -279.485 439.865 -279.225 ;
        RECT 425.870 -279.490 434.635 -279.485 ;
        RECT 368.645 -279.685 371.735 -279.600 ;
        RECT 379.050 -279.680 421.030 -279.495 ;
        RECT 322.880 -279.770 325.970 -279.685 ;
        RECT 333.285 -279.765 374.210 -279.685 ;
        RECT 279.115 -279.870 281.325 -279.800 ;
        RECT 291.350 -279.830 328.445 -279.770 ;
        RECT 170.395 -280.630 194.370 -280.075 ;
        RECT 199.210 -280.390 201.235 -280.070 ;
        RECT 196.395 -280.440 196.885 -280.425 ;
        RECT 199.210 -280.440 199.795 -280.390 ;
        RECT 170.395 -280.665 194.890 -280.630 ;
        RECT 195.255 -280.665 195.565 -280.525 ;
        RECT 162.815 -283.275 162.985 -280.915 ;
        RECT 163.465 -283.275 163.635 -280.900 ;
        RECT 164.605 -282.275 164.775 -280.825 ;
        RECT 165.585 -282.275 165.755 -280.815 ;
        RECT 170.395 -280.840 195.565 -280.665 ;
        RECT 125.475 -287.080 130.995 -287.070 ;
        RECT 100.460 -287.395 130.995 -287.080 ;
        RECT 112.020 -287.400 114.385 -287.395 ;
        RECT 112.970 -288.495 114.130 -287.400 ;
        RECT 125.475 -287.410 130.995 -287.395 ;
        RECT 112.680 -288.815 114.890 -288.495 ;
        RECT -30.565 -291.005 -4.440 -290.690 ;
        RECT -30.565 -291.030 -22.700 -291.005 ;
        RECT -18.210 -291.030 -9.200 -291.005 ;
        RECT -139.180 -294.150 -136.015 -294.080 ;
        RECT -136.945 -294.375 -136.015 -294.150 ;
        RECT -105.820 -294.350 -101.910 -293.655 ;
        RECT -100.030 -294.285 -97.440 -293.655 ;
        RECT -136.945 -295.160 -136.705 -294.375 ;
        RECT -139.180 -295.330 -136.705 -295.160 ;
        RECT -136.945 -295.810 -136.705 -295.330 ;
        RECT -139.180 -295.980 -136.705 -295.810 ;
        RECT -136.945 -296.990 -136.705 -295.980 ;
        RECT -139.180 -297.020 -136.705 -296.990 ;
        RECT -136.345 -297.020 -136.015 -294.375 ;
        RECT -106.120 -295.015 -101.780 -294.350 ;
        RECT -100.105 -294.630 -97.335 -294.285 ;
        RECT -95.585 -294.290 -92.820 -293.655 ;
        RECT -95.585 -294.495 -92.810 -294.290 ;
        RECT -106.120 -295.575 -105.855 -295.015 ;
        RECT -139.180 -297.160 -136.015 -297.020 ;
        RECT -136.945 -297.315 -136.015 -297.160 ;
        RECT -136.945 -298.170 -136.705 -297.315 ;
        RECT -139.180 -298.340 -136.705 -298.170 ;
        RECT -136.345 -298.320 -136.015 -297.315 ;
        RECT -106.075 -298.575 -105.905 -295.575 ;
        RECT -105.140 -295.655 -104.875 -295.015 ;
        RECT -100.080 -295.265 -99.840 -294.630 ;
        RECT -105.095 -298.575 -104.925 -295.655 ;
        RECT -100.045 -297.220 -99.875 -295.265 ;
        RECT -99.095 -295.295 -98.855 -294.630 ;
        RECT -95.580 -294.635 -92.810 -294.495 ;
        RECT -95.555 -295.270 -95.315 -294.635 ;
        RECT -99.065 -297.220 -98.895 -295.295 ;
        RECT -95.520 -297.225 -95.350 -295.270 ;
        RECT -94.570 -295.300 -94.330 -294.635 ;
        RECT -94.540 -297.225 -94.370 -295.300 ;
        RECT -69.935 -298.170 -69.490 -293.655 ;
        RECT -68.200 -298.155 -68.030 -296.700 ;
        RECT -67.220 -298.155 -67.050 -296.700 ;
        RECT -66.240 -298.155 -66.070 -296.700 ;
        RECT -59.485 -298.155 -59.315 -296.700 ;
        RECT -58.505 -298.155 -58.335 -296.700 ;
        RECT -57.525 -298.155 -57.355 -296.700 ;
        RECT -54.700 -298.155 -54.530 -296.700 ;
        RECT -53.720 -298.155 -53.550 -296.700 ;
        RECT -52.740 -298.155 -52.570 -296.700 ;
        RECT -45.985 -298.155 -45.815 -296.700 ;
        RECT -45.005 -298.155 -44.835 -296.700 ;
        RECT -44.025 -298.155 -43.855 -296.700 ;
        RECT -41.575 -298.155 -41.405 -296.700 ;
        RECT -40.595 -298.155 -40.425 -296.700 ;
        RECT -39.615 -298.155 -39.445 -296.700 ;
        RECT -68.500 -298.170 -66.025 -298.155 ;
        RECT -59.790 -298.160 -52.525 -298.155 ;
        RECT -69.935 -298.180 -64.415 -298.170 ;
        RECT -59.790 -298.180 -50.960 -298.160 ;
        RECT -46.290 -298.180 -39.400 -298.155 ;
        RECT -69.935 -298.495 -39.400 -298.180 ;
        RECT -69.935 -298.510 -64.415 -298.495 ;
        RECT -53.325 -298.500 -50.960 -298.495 ;
        RECT -88.510 -301.915 -88.340 -299.830 ;
        RECT -87.530 -301.915 -87.360 -299.830 ;
        RECT -86.550 -301.665 -86.380 -299.830 ;
        RECT -85.465 -301.665 -85.295 -300.835 ;
        RECT -84.485 -301.665 -84.315 -300.835 ;
        RECT -83.505 -301.665 -83.335 -300.835 ;
        RECT -82.525 -301.665 -82.355 -300.835 ;
        RECT -86.550 -301.915 -82.115 -301.665 ;
        RECT -81.275 -301.725 -81.105 -298.775 ;
        RECT -88.560 -302.160 -82.115 -301.915 ;
        RECT -88.560 -302.235 -86.350 -302.160 ;
        RECT -81.300 -302.355 -81.075 -301.725 ;
        RECT -80.295 -301.740 -80.125 -298.775 ;
        RECT -78.180 -301.735 -78.010 -298.775 ;
        RECT -30.565 -299.505 -30.120 -291.030 ;
        RECT -29.320 -292.485 -29.150 -291.030 ;
        RECT -28.340 -292.485 -28.170 -291.030 ;
        RECT -27.360 -292.485 -27.190 -291.030 ;
        RECT -25.135 -292.485 -24.965 -291.030 ;
        RECT -24.155 -292.485 -23.985 -291.030 ;
        RECT -23.175 -292.485 -23.005 -291.030 ;
        RECT -15.820 -292.485 -15.650 -291.030 ;
        RECT -14.840 -292.485 -14.670 -291.030 ;
        RECT -13.860 -292.485 -13.690 -291.030 ;
        RECT -11.635 -292.485 -11.465 -291.030 ;
        RECT -10.655 -292.485 -10.485 -291.030 ;
        RECT -9.675 -292.485 -9.505 -291.030 ;
        RECT 112.730 -291.400 112.900 -288.815 ;
        RECT 113.710 -291.400 113.880 -288.815 ;
        RECT 114.690 -291.400 114.860 -288.815 ;
        RECT -28.830 -299.490 -28.660 -298.035 ;
        RECT -27.850 -299.490 -27.680 -298.035 ;
        RECT -26.870 -299.490 -26.700 -298.035 ;
        RECT -20.115 -299.490 -19.945 -298.035 ;
        RECT -19.135 -299.490 -18.965 -298.035 ;
        RECT -18.155 -299.490 -17.985 -298.035 ;
        RECT -15.330 -299.490 -15.160 -298.035 ;
        RECT -14.350 -299.490 -14.180 -298.035 ;
        RECT -13.370 -299.490 -13.200 -298.035 ;
        RECT -6.615 -299.490 -6.445 -298.035 ;
        RECT -5.635 -299.490 -5.465 -298.035 ;
        RECT -4.655 -299.490 -4.485 -298.035 ;
        RECT -2.205 -299.490 -2.035 -298.035 ;
        RECT -1.225 -299.490 -1.055 -298.035 ;
        RECT -0.245 -299.260 -0.075 -298.035 ;
        RECT -0.605 -299.490 0.010 -299.260 ;
        RECT 1.465 -299.265 1.635 -297.950 ;
        RECT -29.130 -299.505 -26.655 -299.490 ;
        RECT -20.420 -299.495 -13.155 -299.490 ;
        RECT -30.565 -299.515 -25.045 -299.505 ;
        RECT -20.420 -299.515 -11.590 -299.495 ;
        RECT -6.920 -299.515 0.010 -299.490 ;
        RECT -30.565 -299.830 0.010 -299.515 ;
        RECT -30.565 -299.845 -25.045 -299.830 ;
        RECT -80.325 -302.355 -80.100 -301.740 ;
        RECT -78.215 -302.355 -77.990 -301.735 ;
        RECT -86.365 -302.440 -85.420 -302.405 ;
        RECT -86.550 -302.475 -85.420 -302.440 ;
        RECT -81.330 -302.475 -77.485 -302.355 ;
        RECT -94.730 -302.685 -77.485 -302.475 ;
        RECT -19.710 -302.590 -19.135 -299.830 ;
        RECT -13.955 -299.835 -11.590 -299.830 ;
        RECT -94.730 -303.240 -78.005 -302.685 ;
        RECT -94.730 -303.335 -86.850 -303.240 ;
        RECT -94.730 -308.310 -93.870 -303.335 ;
        RECT -87.710 -304.190 -86.850 -303.335 ;
        RECT -83.570 -303.325 -80.480 -303.240 ;
        RECT -19.735 -303.270 -19.120 -302.590 ;
        RECT -6.880 -303.310 -6.305 -299.830 ;
        RECT -0.605 -299.940 0.010 -299.830 ;
        RECT 0.865 -299.410 1.635 -299.265 ;
        RECT 2.445 -299.410 2.615 -297.950 ;
        RECT 0.865 -299.415 2.640 -299.410 ;
        RECT 5.155 -299.415 5.325 -297.950 ;
        RECT 6.135 -299.415 6.305 -297.950 ;
        RECT 7.115 -299.415 7.285 -297.950 ;
        RECT 8.095 -299.415 8.265 -297.950 ;
        RECT 10.130 -299.215 10.300 -298.385 ;
        RECT 11.110 -299.215 11.280 -298.385 ;
        RECT 12.090 -299.215 12.260 -298.385 ;
        RECT 13.070 -299.215 13.240 -298.385 ;
        RECT 14.155 -299.215 14.325 -297.380 ;
        RECT 9.890 -299.415 14.325 -299.215 ;
        RECT 15.135 -299.415 15.305 -297.380 ;
        RECT 16.115 -299.200 16.285 -297.380 ;
        RECT 15.755 -299.415 16.370 -299.200 ;
        RECT 18.155 -299.205 18.325 -298.375 ;
        RECT 19.135 -299.205 19.305 -298.375 ;
        RECT 20.115 -299.205 20.285 -298.375 ;
        RECT 21.095 -299.205 21.265 -298.375 ;
        RECT 22.180 -299.205 22.350 -297.370 ;
        RECT 0.865 -299.810 16.370 -299.415 ;
        RECT 0.865 -299.945 1.480 -299.810 ;
        RECT -83.570 -303.470 -81.355 -303.325 ;
        RECT -83.565 -303.540 -81.355 -303.470 ;
        RECT -83.565 -303.785 -77.120 -303.540 ;
        RECT -88.620 -304.685 -85.030 -304.190 ;
        RECT -88.380 -306.015 -88.210 -304.685 ;
        RECT -87.400 -306.015 -87.230 -304.685 ;
        RECT -86.420 -306.015 -86.250 -304.685 ;
        RECT -85.440 -306.015 -85.270 -304.685 ;
        RECT -83.515 -305.870 -83.345 -303.785 ;
        RECT -82.535 -305.870 -82.365 -303.785 ;
        RECT -81.555 -304.035 -77.120 -303.785 ;
        RECT -6.900 -303.990 -6.285 -303.310 ;
        RECT 5.540 -303.850 6.115 -299.810 ;
        RECT 15.755 -299.880 16.370 -299.810 ;
        RECT 17.700 -299.455 22.350 -299.205 ;
        RECT 23.160 -299.455 23.330 -297.370 ;
        RECT 24.140 -299.320 24.310 -297.370 ;
        RECT 93.875 -297.685 94.045 -295.730 ;
        RECT 94.855 -297.655 95.025 -295.730 ;
        RECT 23.840 -299.455 24.455 -299.320 ;
        RECT 26.275 -299.330 26.445 -297.995 ;
        RECT 17.700 -299.700 24.455 -299.455 ;
        RECT 17.700 -299.885 18.315 -299.700 ;
        RECT 22.150 -299.775 24.455 -299.700 ;
        RECT 23.840 -300.000 24.455 -299.775 ;
        RECT 25.845 -299.455 26.460 -299.330 ;
        RECT 27.255 -299.455 27.425 -297.995 ;
        RECT 25.845 -299.480 27.450 -299.455 ;
        RECT 29.965 -299.475 30.135 -297.995 ;
        RECT 30.945 -299.475 31.115 -297.995 ;
        RECT 31.925 -299.475 32.095 -297.995 ;
        RECT 32.905 -299.305 33.075 -297.995 ;
        RECT 38.710 -298.855 38.880 -297.940 ;
        RECT 39.690 -298.855 39.860 -297.940 ;
        RECT 38.710 -299.300 38.910 -298.855 ;
        RECT 32.625 -299.475 33.240 -299.305 ;
        RECT 29.965 -299.480 33.240 -299.475 ;
        RECT 25.845 -299.820 33.240 -299.480 ;
        RECT 25.845 -299.845 30.325 -299.820 ;
        RECT 25.845 -300.010 26.460 -299.845 ;
        RECT 32.625 -299.985 33.240 -299.820 ;
        RECT 38.705 -299.500 39.320 -299.300 ;
        RECT 39.655 -299.500 39.885 -298.855 ;
        RECT 40.670 -298.875 40.840 -297.940 ;
        RECT 41.240 -298.855 41.410 -297.940 ;
        RECT 40.645 -299.500 40.875 -298.875 ;
        RECT 41.210 -299.500 41.440 -298.855 ;
        RECT 42.220 -298.880 42.390 -297.940 ;
        RECT 42.785 -298.830 42.955 -297.940 ;
        RECT 42.190 -299.500 42.420 -298.880 ;
        RECT 42.755 -299.500 42.985 -298.830 ;
        RECT 43.765 -298.890 43.935 -297.940 ;
        RECT 93.840 -298.320 94.080 -297.685 ;
        RECT 94.825 -298.320 95.065 -297.655 ;
        RECT 98.605 -297.685 98.775 -295.730 ;
        RECT 99.585 -297.655 99.755 -295.730 ;
        RECT 98.570 -298.320 98.810 -297.685 ;
        RECT 99.555 -298.320 99.795 -297.655 ;
        RECT 101.960 -298.320 102.390 -298.280 ;
        RECT 89.725 -298.380 102.390 -298.320 ;
        RECT 103.185 -298.380 103.355 -296.900 ;
        RECT 104.165 -298.380 104.335 -296.900 ;
        RECT 105.145 -298.380 105.315 -296.900 ;
        RECT 106.125 -298.380 106.295 -296.900 ;
        RECT 107.560 -298.360 107.875 -298.290 ;
        RECT 108.835 -298.360 109.005 -296.900 ;
        RECT 109.815 -298.360 109.985 -296.900 ;
        RECT 110.965 -298.320 111.335 -298.290 ;
        RECT 112.480 -298.320 112.650 -296.865 ;
        RECT 113.460 -298.320 113.630 -296.865 ;
        RECT 114.440 -298.185 114.610 -296.865 ;
        RECT 116.880 -298.185 117.050 -294.010 ;
        RECT 117.860 -298.185 118.030 -294.010 ;
        RECT 118.880 -298.185 119.050 -294.010 ;
        RECT 119.860 -298.185 120.030 -294.010 ;
        RECT 121.880 -298.185 122.050 -294.010 ;
        RECT 122.860 -298.185 123.030 -294.010 ;
        RECT 123.880 -298.185 124.050 -294.010 ;
        RECT 124.860 -298.185 125.030 -294.010 ;
        RECT 126.880 -298.185 127.050 -294.010 ;
        RECT 127.860 -298.185 128.030 -294.010 ;
        RECT 128.880 -298.185 129.050 -294.010 ;
        RECT 129.860 -298.185 130.030 -294.010 ;
        RECT 130.550 -298.185 130.995 -287.410 ;
        RECT 154.230 -290.960 156.240 -290.630 ;
        RECT 141.755 -295.840 141.925 -294.510 ;
        RECT 142.735 -295.840 142.905 -294.510 ;
        RECT 143.715 -295.840 143.885 -294.510 ;
        RECT 144.695 -295.840 144.865 -294.510 ;
        RECT 141.515 -296.335 145.105 -295.840 ;
        RECT 142.425 -297.285 143.285 -296.335 ;
        RECT 146.620 -296.740 146.790 -294.655 ;
        RECT 147.600 -296.740 147.770 -294.655 ;
        RECT 148.580 -296.490 148.750 -294.655 ;
        RECT 149.665 -296.490 149.835 -295.660 ;
        RECT 150.645 -296.490 150.815 -295.660 ;
        RECT 151.625 -296.490 151.795 -295.660 ;
        RECT 152.605 -296.490 152.775 -295.660 ;
        RECT 148.580 -296.740 153.015 -296.490 ;
        RECT 146.570 -296.985 153.015 -296.740 ;
        RECT 146.570 -297.055 148.780 -296.985 ;
        RECT 146.565 -297.200 148.780 -297.055 ;
        RECT 146.565 -297.285 149.655 -297.200 ;
        RECT 141.575 -297.840 152.130 -297.285 ;
        RECT 154.230 -297.465 154.560 -290.960 ;
        RECT 141.575 -298.050 152.650 -297.840 ;
        RECT 154.145 -298.030 154.565 -297.465 ;
        RECT 155.910 -297.610 156.240 -290.960 ;
        RECT 170.395 -291.995 171.005 -280.840 ;
        RECT 185.825 -280.875 186.955 -280.840 ;
        RECT 186.010 -280.910 186.955 -280.875 ;
        RECT 191.045 -280.925 195.565 -280.840 ;
        RECT 191.045 -280.960 194.890 -280.925 ;
        RECT 183.815 -281.155 186.025 -281.080 ;
        RECT 183.815 -281.400 190.260 -281.155 ;
        RECT 183.865 -283.485 184.035 -281.400 ;
        RECT 184.845 -283.485 185.015 -281.400 ;
        RECT 185.825 -281.650 190.260 -281.400 ;
        RECT 191.075 -281.590 191.300 -280.960 ;
        RECT 192.050 -281.575 192.275 -280.960 ;
        RECT 185.825 -283.485 185.995 -281.650 ;
        RECT 186.910 -282.480 187.080 -281.650 ;
        RECT 187.890 -282.480 188.060 -281.650 ;
        RECT 188.870 -282.480 189.040 -281.650 ;
        RECT 189.850 -282.480 190.020 -281.650 ;
        RECT 191.100 -284.540 191.270 -281.590 ;
        RECT 192.080 -284.540 192.250 -281.575 ;
        RECT 194.160 -281.580 194.385 -280.960 ;
        RECT 195.255 -280.995 195.565 -280.925 ;
        RECT 196.395 -281.025 199.795 -280.440 ;
        RECT 201.045 -280.865 201.235 -280.390 ;
        RECT 202.030 -280.855 202.220 -280.070 ;
        RECT 196.395 -281.055 196.885 -281.025 ;
        RECT 194.195 -284.540 194.365 -281.580 ;
        RECT 201.060 -283.330 201.230 -280.865 ;
        RECT 202.040 -283.330 202.210 -280.855 ;
        RECT 204.990 -280.970 205.240 -280.070 ;
        RECT 205.620 -280.955 205.870 -280.070 ;
        RECT 206.775 -280.880 206.990 -280.070 ;
        RECT 207.760 -280.270 229.840 -280.070 ;
        RECT 233.120 -280.185 235.335 -280.040 ;
        RECT 243.525 -280.100 275.830 -280.000 ;
        RECT 279.110 -280.015 281.325 -279.870 ;
        RECT 279.110 -280.100 282.200 -280.015 ;
        RECT 289.515 -280.095 328.445 -279.830 ;
        RECT 233.120 -280.270 236.210 -280.185 ;
        RECT 243.525 -280.265 284.675 -280.100 ;
        RECT 207.760 -280.515 238.685 -280.270 ;
        RECT 207.760 -280.870 207.975 -280.515 ;
        RECT 205.015 -283.330 205.185 -280.970 ;
        RECT 205.665 -283.330 205.835 -280.955 ;
        RECT 206.805 -282.330 206.975 -280.880 ;
        RECT 207.785 -282.330 207.955 -280.870 ;
        RECT 196.430 -291.015 198.440 -290.685 ;
        RECT 170.395 -292.605 173.555 -291.995 ;
        RECT 160.095 -295.995 160.265 -294.665 ;
        RECT 161.075 -295.995 161.245 -294.665 ;
        RECT 162.055 -295.995 162.225 -294.665 ;
        RECT 163.035 -295.995 163.205 -294.665 ;
        RECT 159.855 -296.490 163.445 -295.995 ;
        RECT 160.765 -297.440 161.625 -296.490 ;
        RECT 164.960 -296.895 165.130 -294.810 ;
        RECT 165.940 -296.895 166.110 -294.810 ;
        RECT 166.920 -296.645 167.090 -294.810 ;
        RECT 168.005 -296.645 168.175 -295.815 ;
        RECT 168.985 -296.645 169.155 -295.815 ;
        RECT 169.965 -296.645 170.135 -295.815 ;
        RECT 170.945 -296.645 171.115 -295.815 ;
        RECT 166.920 -296.895 171.355 -296.645 ;
        RECT 164.910 -297.140 171.355 -296.895 ;
        RECT 164.910 -297.210 167.120 -297.140 ;
        RECT 164.905 -297.355 167.120 -297.210 ;
        RECT 164.905 -297.440 167.995 -297.355 ;
        RECT 159.915 -297.610 170.470 -297.440 ;
        RECT 172.945 -297.585 173.555 -292.605 ;
        RECT 183.955 -295.895 184.125 -294.565 ;
        RECT 184.935 -295.895 185.105 -294.565 ;
        RECT 185.915 -295.895 186.085 -294.565 ;
        RECT 186.895 -295.895 187.065 -294.565 ;
        RECT 183.715 -296.390 187.305 -295.895 ;
        RECT 184.625 -297.340 185.485 -296.390 ;
        RECT 188.820 -296.795 188.990 -294.710 ;
        RECT 189.800 -296.795 189.970 -294.710 ;
        RECT 190.780 -296.545 190.950 -294.710 ;
        RECT 191.865 -296.545 192.035 -295.715 ;
        RECT 192.845 -296.545 193.015 -295.715 ;
        RECT 193.825 -296.545 193.995 -295.715 ;
        RECT 194.805 -296.545 194.975 -295.715 ;
        RECT 190.780 -296.795 195.215 -296.545 ;
        RECT 188.770 -297.040 195.215 -296.795 ;
        RECT 188.770 -297.110 190.980 -297.040 ;
        RECT 188.765 -297.255 190.980 -297.110 ;
        RECT 188.765 -297.340 191.855 -297.255 ;
        RECT 155.910 -297.940 170.470 -297.610 ;
        RECT 171.245 -297.815 171.640 -297.660 ;
        RECT 159.915 -297.995 170.470 -297.940 ;
        RECT 170.745 -297.995 171.640 -297.815 ;
        RECT 143.585 -298.085 144.715 -298.050 ;
        RECT 143.770 -298.120 144.715 -298.085 ;
        RECT 148.805 -298.170 152.650 -298.050 ;
        RECT 114.440 -298.320 130.995 -298.185 ;
        RECT 110.965 -298.360 130.995 -298.320 ;
        RECT 107.560 -298.380 130.995 -298.360 ;
        RECT 89.725 -298.660 130.995 -298.380 ;
        RECT 141.575 -298.365 143.785 -298.290 ;
        RECT 141.575 -298.610 148.020 -298.365 ;
        RECT 89.725 -298.665 111.335 -298.660 ;
        RECT 43.740 -299.500 43.970 -298.890 ;
        RECT 38.705 -299.845 43.970 -299.500 ;
        RECT 38.705 -299.980 39.320 -299.845 ;
        RECT 89.725 -301.020 90.355 -298.665 ;
        RECT 101.960 -298.695 111.335 -298.665 ;
        RECT 101.960 -298.725 107.875 -298.695 ;
        RECT 110.965 -298.725 111.335 -298.695 ;
        RECT 114.550 -298.700 130.995 -298.660 ;
        RECT 101.960 -298.745 102.390 -298.725 ;
        RECT 107.560 -298.780 107.875 -298.725 ;
        RECT 141.625 -300.695 141.795 -298.610 ;
        RECT 142.605 -300.695 142.775 -298.610 ;
        RECT 143.585 -298.860 148.020 -298.610 ;
        RECT 148.835 -298.800 149.060 -298.170 ;
        RECT 149.810 -298.785 150.035 -298.170 ;
        RECT 143.585 -300.695 143.755 -298.860 ;
        RECT 144.670 -299.690 144.840 -298.860 ;
        RECT 145.650 -299.690 145.820 -298.860 ;
        RECT 146.630 -299.690 146.800 -298.860 ;
        RECT 147.610 -299.690 147.780 -298.860 ;
        RECT 71.380 -301.035 73.745 -301.030 ;
        RECT 84.835 -301.035 90.355 -301.020 ;
        RECT 59.820 -301.350 90.355 -301.035 ;
        RECT 59.820 -301.375 66.710 -301.350 ;
        RECT 71.380 -301.370 80.210 -301.350 ;
        RECT 84.835 -301.360 90.355 -301.350 ;
        RECT 72.945 -301.375 80.210 -301.370 ;
        RECT 86.445 -301.375 88.920 -301.360 ;
        RECT 59.865 -302.830 60.035 -301.375 ;
        RECT 60.845 -302.830 61.015 -301.375 ;
        RECT 61.825 -302.830 61.995 -301.375 ;
        RECT 64.275 -302.830 64.445 -301.375 ;
        RECT 65.255 -302.830 65.425 -301.375 ;
        RECT 66.235 -302.830 66.405 -301.375 ;
        RECT 72.990 -302.830 73.160 -301.375 ;
        RECT 73.970 -302.830 74.140 -301.375 ;
        RECT 74.950 -302.830 75.120 -301.375 ;
        RECT 77.775 -302.830 77.945 -301.375 ;
        RECT 78.755 -302.830 78.925 -301.375 ;
        RECT 79.735 -302.830 79.905 -301.375 ;
        RECT 86.490 -302.830 86.660 -301.375 ;
        RECT 87.470 -302.830 87.640 -301.375 ;
        RECT 88.450 -302.830 88.620 -301.375 ;
        RECT -81.555 -305.870 -81.385 -304.035 ;
        RECT -80.470 -304.865 -80.300 -304.035 ;
        RECT -79.490 -304.865 -79.320 -304.035 ;
        RECT -78.510 -304.865 -78.340 -304.035 ;
        RECT -77.530 -304.865 -77.360 -304.035 ;
        RECT 5.515 -304.160 7.045 -303.850 ;
        RECT 5.515 -304.165 6.130 -304.160 ;
        RECT -19.730 -307.105 -19.115 -306.425 ;
        RECT -6.895 -306.930 -6.280 -306.250 ;
        RECT 5.520 -306.930 6.135 -306.250 ;
        RECT -94.740 -308.745 -93.860 -308.310 ;
        RECT -107.760 -311.085 -107.590 -309.625 ;
        RECT -106.780 -311.005 -106.610 -309.625 ;
        RECT -104.070 -311.005 -103.900 -309.625 ;
        RECT -103.090 -311.005 -102.920 -309.625 ;
        RECT -102.110 -311.005 -101.940 -309.625 ;
        RECT -101.130 -311.005 -100.960 -309.625 ;
        RECT -26.340 -310.110 -26.170 -309.195 ;
        RECT -25.360 -310.110 -25.190 -309.195 ;
        RECT -26.340 -310.755 -26.140 -310.110 ;
        RECT -25.395 -310.755 -25.165 -310.110 ;
        RECT -24.380 -310.130 -24.210 -309.195 ;
        RECT -23.810 -310.110 -23.640 -309.195 ;
        RECT -24.405 -310.755 -24.175 -310.130 ;
        RECT -23.840 -310.755 -23.610 -310.110 ;
        RECT -22.830 -310.135 -22.660 -309.195 ;
        RECT -22.265 -310.085 -22.095 -309.195 ;
        RECT -22.860 -310.755 -22.630 -310.135 ;
        RECT -22.295 -310.755 -22.065 -310.085 ;
        RECT -21.285 -310.145 -21.115 -309.195 ;
        RECT -21.310 -310.755 -21.080 -310.145 ;
        RECT -106.870 -311.085 -93.860 -311.005 ;
        RECT -107.810 -311.420 -93.860 -311.085 ;
        RECT -26.340 -311.290 -21.080 -310.755 ;
        RECT -19.705 -311.290 -19.130 -307.105 ;
        RECT -13.840 -310.110 -13.670 -309.195 ;
        RECT -12.860 -310.110 -12.690 -309.195 ;
        RECT -13.840 -310.755 -13.640 -310.110 ;
        RECT -12.895 -310.755 -12.665 -310.110 ;
        RECT -11.880 -310.130 -11.710 -309.195 ;
        RECT -11.310 -310.110 -11.140 -309.195 ;
        RECT -11.905 -310.755 -11.675 -310.130 ;
        RECT -11.340 -310.755 -11.110 -310.110 ;
        RECT -10.330 -310.135 -10.160 -309.195 ;
        RECT -9.765 -310.085 -9.595 -309.195 ;
        RECT -10.360 -310.755 -10.130 -310.135 ;
        RECT -9.795 -310.755 -9.565 -310.085 ;
        RECT -8.785 -310.145 -8.615 -309.195 ;
        RECT -8.810 -310.755 -8.580 -310.145 ;
        RECT -13.840 -311.100 -8.580 -310.755 ;
        RECT -12.270 -311.290 -9.305 -311.100 ;
        RECT -6.865 -311.290 -6.295 -306.930 ;
        RECT -1.340 -310.110 -1.170 -309.195 ;
        RECT -0.360 -310.110 -0.190 -309.195 ;
        RECT -1.340 -310.755 -1.140 -310.110 ;
        RECT -0.395 -310.755 -0.165 -310.110 ;
        RECT 0.620 -310.130 0.790 -309.195 ;
        RECT 1.190 -310.110 1.360 -309.195 ;
        RECT 0.595 -310.755 0.825 -310.130 ;
        RECT 1.160 -310.755 1.390 -310.110 ;
        RECT 2.170 -310.135 2.340 -309.195 ;
        RECT 2.735 -310.085 2.905 -309.195 ;
        RECT 2.140 -310.755 2.370 -310.135 ;
        RECT 2.705 -310.755 2.935 -310.085 ;
        RECT 3.715 -310.145 3.885 -309.195 ;
        RECT 3.690 -310.755 3.920 -310.145 ;
        RECT -1.340 -311.100 3.920 -310.755 ;
        RECT 0.310 -311.290 3.275 -311.100 ;
        RECT 5.545 -311.290 6.120 -306.930 ;
        RECT 11.160 -310.110 11.330 -309.195 ;
        RECT 12.140 -310.110 12.310 -309.195 ;
        RECT 11.160 -310.755 11.360 -310.110 ;
        RECT 12.105 -310.755 12.335 -310.110 ;
        RECT 13.120 -310.130 13.290 -309.195 ;
        RECT 13.690 -310.110 13.860 -309.195 ;
        RECT 13.095 -310.755 13.325 -310.130 ;
        RECT 13.660 -310.755 13.890 -310.110 ;
        RECT 14.670 -310.135 14.840 -309.195 ;
        RECT 15.235 -310.085 15.405 -309.195 ;
        RECT 14.640 -310.755 14.870 -310.135 ;
        RECT 15.205 -310.755 15.435 -310.085 ;
        RECT 16.215 -310.145 16.385 -309.195 ;
        RECT 23.660 -310.110 23.830 -309.195 ;
        RECT 24.640 -310.110 24.810 -309.195 ;
        RECT 16.190 -310.755 16.420 -310.145 ;
        RECT 11.160 -311.100 16.420 -310.755 ;
        RECT 23.660 -310.755 23.860 -310.110 ;
        RECT 24.605 -310.755 24.835 -310.110 ;
        RECT 25.620 -310.130 25.790 -309.195 ;
        RECT 26.190 -310.110 26.360 -309.195 ;
        RECT 25.595 -310.755 25.825 -310.130 ;
        RECT 26.160 -310.755 26.390 -310.110 ;
        RECT 27.170 -310.135 27.340 -309.195 ;
        RECT 27.735 -310.085 27.905 -309.195 ;
        RECT 27.140 -310.755 27.370 -310.135 ;
        RECT 27.705 -310.755 27.935 -310.085 ;
        RECT 28.715 -310.145 28.885 -309.195 ;
        RECT 38.660 -310.110 38.830 -309.195 ;
        RECT 39.640 -310.110 39.810 -309.195 ;
        RECT 28.690 -310.755 28.920 -310.145 ;
        RECT 23.660 -311.100 28.920 -310.755 ;
        RECT 38.660 -310.755 38.860 -310.110 ;
        RECT 39.605 -310.755 39.835 -310.110 ;
        RECT 40.620 -310.130 40.790 -309.195 ;
        RECT 41.190 -310.110 41.360 -309.195 ;
        RECT 40.595 -310.755 40.825 -310.130 ;
        RECT 41.160 -310.755 41.390 -310.110 ;
        RECT 42.170 -310.135 42.340 -309.195 ;
        RECT 42.735 -310.085 42.905 -309.195 ;
        RECT 42.140 -310.755 42.370 -310.135 ;
        RECT 42.705 -310.755 42.935 -310.085 ;
        RECT 43.715 -310.145 43.885 -309.195 ;
        RECT 69.295 -309.835 69.465 -308.380 ;
        RECT 70.275 -309.835 70.445 -308.380 ;
        RECT 71.255 -309.835 71.425 -308.380 ;
        RECT 73.480 -309.835 73.650 -308.380 ;
        RECT 74.460 -309.835 74.630 -308.380 ;
        RECT 75.440 -309.835 75.610 -308.380 ;
        RECT 82.795 -309.835 82.965 -308.380 ;
        RECT 83.775 -309.835 83.945 -308.380 ;
        RECT 84.755 -309.835 84.925 -308.380 ;
        RECT 86.980 -309.835 87.150 -308.380 ;
        RECT 87.960 -309.835 88.130 -308.380 ;
        RECT 88.940 -309.835 89.110 -308.380 ;
        RECT 89.910 -309.835 90.355 -301.360 ;
        RECT 148.860 -301.750 149.030 -298.800 ;
        RECT 149.840 -301.750 150.010 -298.785 ;
        RECT 151.920 -298.790 152.145 -298.170 ;
        RECT 159.915 -298.205 171.640 -297.995 ;
        RECT 161.925 -298.240 163.055 -298.205 ;
        RECT 162.110 -298.275 163.055 -298.240 ;
        RECT 167.145 -298.230 171.640 -298.205 ;
        RECT 167.145 -298.325 170.990 -298.230 ;
        RECT 159.915 -298.520 162.125 -298.445 ;
        RECT 159.915 -298.765 166.360 -298.520 ;
        RECT 151.955 -301.750 152.125 -298.790 ;
        RECT 159.965 -300.850 160.135 -298.765 ;
        RECT 160.945 -300.850 161.115 -298.765 ;
        RECT 161.925 -299.015 166.360 -298.765 ;
        RECT 167.175 -298.955 167.400 -298.325 ;
        RECT 168.150 -298.940 168.375 -298.325 ;
        RECT 161.925 -300.850 162.095 -299.015 ;
        RECT 163.010 -299.845 163.180 -299.015 ;
        RECT 163.990 -299.845 164.160 -299.015 ;
        RECT 164.970 -299.845 165.140 -299.015 ;
        RECT 165.950 -299.845 166.120 -299.015 ;
        RECT 167.200 -301.905 167.370 -298.955 ;
        RECT 168.180 -301.905 168.350 -298.940 ;
        RECT 170.260 -298.945 170.485 -298.325 ;
        RECT 171.245 -298.355 171.640 -298.230 ;
        RECT 172.495 -298.280 173.555 -297.585 ;
        RECT 183.775 -297.895 194.330 -297.340 ;
        RECT 196.430 -297.520 196.760 -291.015 ;
        RECT 183.775 -298.105 194.850 -297.895 ;
        RECT 196.345 -298.085 196.765 -297.520 ;
        RECT 198.110 -297.665 198.440 -291.015 ;
        RECT 212.595 -292.050 213.205 -280.515 ;
        RECT 228.130 -280.825 238.685 -280.515 ;
        RECT 243.525 -280.585 245.550 -280.265 ;
        RECT 240.710 -280.635 241.200 -280.620 ;
        RECT 243.525 -280.635 244.110 -280.585 ;
        RECT 228.130 -280.860 239.205 -280.825 ;
        RECT 239.570 -280.860 239.880 -280.720 ;
        RECT 228.130 -281.035 239.880 -280.860 ;
        RECT 230.140 -281.070 231.270 -281.035 ;
        RECT 230.325 -281.105 231.270 -281.070 ;
        RECT 235.360 -281.120 239.880 -281.035 ;
        RECT 235.360 -281.155 239.205 -281.120 ;
        RECT 228.130 -281.350 230.340 -281.275 ;
        RECT 228.130 -281.595 234.575 -281.350 ;
        RECT 228.180 -283.680 228.350 -281.595 ;
        RECT 229.160 -283.680 229.330 -281.595 ;
        RECT 230.140 -281.845 234.575 -281.595 ;
        RECT 235.390 -281.785 235.615 -281.155 ;
        RECT 236.365 -281.770 236.590 -281.155 ;
        RECT 230.140 -283.680 230.310 -281.845 ;
        RECT 231.225 -282.675 231.395 -281.845 ;
        RECT 232.205 -282.675 232.375 -281.845 ;
        RECT 233.185 -282.675 233.355 -281.845 ;
        RECT 234.165 -282.675 234.335 -281.845 ;
        RECT 235.415 -284.735 235.585 -281.785 ;
        RECT 236.395 -284.735 236.565 -281.770 ;
        RECT 238.475 -281.775 238.700 -281.155 ;
        RECT 239.570 -281.190 239.880 -281.120 ;
        RECT 240.710 -281.220 244.110 -280.635 ;
        RECT 245.360 -281.060 245.550 -280.585 ;
        RECT 246.345 -281.050 246.535 -280.265 ;
        RECT 240.710 -281.250 241.200 -281.220 ;
        RECT 238.510 -284.735 238.680 -281.775 ;
        RECT 245.375 -283.525 245.545 -281.060 ;
        RECT 246.355 -283.525 246.525 -281.050 ;
        RECT 249.305 -281.165 249.555 -280.265 ;
        RECT 249.935 -281.150 250.185 -280.265 ;
        RECT 251.090 -281.075 251.305 -280.265 ;
        RECT 252.075 -280.565 284.675 -280.265 ;
        RECT 289.515 -280.415 291.540 -280.095 ;
        RECT 286.700 -280.465 287.190 -280.450 ;
        RECT 289.515 -280.465 290.100 -280.415 ;
        RECT 252.075 -281.065 252.290 -280.565 ;
        RECT 249.330 -283.525 249.500 -281.165 ;
        RECT 249.980 -283.525 250.150 -281.150 ;
        RECT 251.120 -282.525 251.290 -281.075 ;
        RECT 252.100 -282.525 252.270 -281.065 ;
        RECT 240.745 -291.210 242.755 -290.880 ;
        RECT 212.595 -292.660 215.755 -292.050 ;
        RECT 202.295 -296.050 202.465 -294.720 ;
        RECT 203.275 -296.050 203.445 -294.720 ;
        RECT 204.255 -296.050 204.425 -294.720 ;
        RECT 205.235 -296.050 205.405 -294.720 ;
        RECT 202.055 -296.545 205.645 -296.050 ;
        RECT 202.965 -297.495 203.825 -296.545 ;
        RECT 207.160 -296.950 207.330 -294.865 ;
        RECT 208.140 -296.950 208.310 -294.865 ;
        RECT 209.120 -296.700 209.290 -294.865 ;
        RECT 210.205 -296.700 210.375 -295.870 ;
        RECT 211.185 -296.700 211.355 -295.870 ;
        RECT 212.165 -296.700 212.335 -295.870 ;
        RECT 213.145 -296.700 213.315 -295.870 ;
        RECT 209.120 -296.950 213.555 -296.700 ;
        RECT 207.110 -297.195 213.555 -296.950 ;
        RECT 207.110 -297.265 209.320 -297.195 ;
        RECT 207.105 -297.410 209.320 -297.265 ;
        RECT 207.105 -297.495 210.195 -297.410 ;
        RECT 202.115 -297.665 212.670 -297.495 ;
        RECT 215.145 -297.640 215.755 -292.660 ;
        RECT 228.270 -296.090 228.440 -294.760 ;
        RECT 229.250 -296.090 229.420 -294.760 ;
        RECT 230.230 -296.090 230.400 -294.760 ;
        RECT 231.210 -296.090 231.380 -294.760 ;
        RECT 228.030 -296.585 231.620 -296.090 ;
        RECT 228.940 -297.535 229.800 -296.585 ;
        RECT 233.135 -296.990 233.305 -294.905 ;
        RECT 234.115 -296.990 234.285 -294.905 ;
        RECT 235.095 -296.740 235.265 -294.905 ;
        RECT 236.180 -296.740 236.350 -295.910 ;
        RECT 237.160 -296.740 237.330 -295.910 ;
        RECT 238.140 -296.740 238.310 -295.910 ;
        RECT 239.120 -296.740 239.290 -295.910 ;
        RECT 235.095 -296.990 239.530 -296.740 ;
        RECT 233.085 -297.235 239.530 -296.990 ;
        RECT 233.085 -297.305 235.295 -297.235 ;
        RECT 233.080 -297.450 235.295 -297.305 ;
        RECT 233.080 -297.535 236.170 -297.450 ;
        RECT 198.110 -297.995 212.670 -297.665 ;
        RECT 213.445 -297.870 213.840 -297.715 ;
        RECT 202.115 -298.050 212.670 -297.995 ;
        RECT 212.945 -298.050 213.840 -297.870 ;
        RECT 185.785 -298.140 186.915 -298.105 ;
        RECT 185.970 -298.175 186.915 -298.140 ;
        RECT 191.005 -298.225 194.850 -298.105 ;
        RECT 172.495 -298.420 173.190 -298.280 ;
        RECT 183.775 -298.420 185.985 -298.345 ;
        RECT 183.775 -298.665 190.220 -298.420 ;
        RECT 170.295 -301.905 170.465 -298.945 ;
        RECT 183.825 -300.750 183.995 -298.665 ;
        RECT 184.805 -300.750 184.975 -298.665 ;
        RECT 185.785 -298.915 190.220 -298.665 ;
        RECT 191.035 -298.855 191.260 -298.225 ;
        RECT 192.010 -298.840 192.235 -298.225 ;
        RECT 185.785 -300.750 185.955 -298.915 ;
        RECT 186.870 -299.745 187.040 -298.915 ;
        RECT 187.850 -299.745 188.020 -298.915 ;
        RECT 188.830 -299.745 189.000 -298.915 ;
        RECT 189.810 -299.745 189.980 -298.915 ;
        RECT 191.060 -301.805 191.230 -298.855 ;
        RECT 192.040 -301.805 192.210 -298.840 ;
        RECT 194.120 -298.845 194.345 -298.225 ;
        RECT 202.115 -298.260 213.840 -298.050 ;
        RECT 204.125 -298.295 205.255 -298.260 ;
        RECT 204.310 -298.330 205.255 -298.295 ;
        RECT 209.345 -298.285 213.840 -298.260 ;
        RECT 209.345 -298.380 213.190 -298.285 ;
        RECT 202.115 -298.575 204.325 -298.500 ;
        RECT 202.115 -298.820 208.560 -298.575 ;
        RECT 194.155 -301.805 194.325 -298.845 ;
        RECT 202.165 -300.905 202.335 -298.820 ;
        RECT 203.145 -300.905 203.315 -298.820 ;
        RECT 204.125 -299.070 208.560 -298.820 ;
        RECT 209.375 -299.010 209.600 -298.380 ;
        RECT 210.350 -298.995 210.575 -298.380 ;
        RECT 204.125 -300.905 204.295 -299.070 ;
        RECT 205.210 -299.900 205.380 -299.070 ;
        RECT 206.190 -299.900 206.360 -299.070 ;
        RECT 207.170 -299.900 207.340 -299.070 ;
        RECT 208.150 -299.900 208.320 -299.070 ;
        RECT 209.400 -301.960 209.570 -299.010 ;
        RECT 210.380 -301.960 210.550 -298.995 ;
        RECT 212.460 -299.000 212.685 -298.380 ;
        RECT 213.445 -298.410 213.840 -298.285 ;
        RECT 214.695 -298.335 215.755 -297.640 ;
        RECT 228.090 -298.090 238.645 -297.535 ;
        RECT 240.745 -297.715 241.075 -291.210 ;
        RECT 228.090 -298.300 239.165 -298.090 ;
        RECT 240.660 -298.280 241.080 -297.715 ;
        RECT 242.425 -297.860 242.755 -291.210 ;
        RECT 256.910 -292.245 257.520 -280.565 ;
        RECT 274.120 -280.655 284.675 -280.565 ;
        RECT 274.120 -280.690 285.195 -280.655 ;
        RECT 285.560 -280.690 285.870 -280.550 ;
        RECT 274.120 -280.865 285.870 -280.690 ;
        RECT 276.130 -280.900 277.260 -280.865 ;
        RECT 276.315 -280.935 277.260 -280.900 ;
        RECT 281.350 -280.950 285.870 -280.865 ;
        RECT 281.350 -280.985 285.195 -280.950 ;
        RECT 274.120 -281.180 276.330 -281.105 ;
        RECT 274.120 -281.425 280.565 -281.180 ;
        RECT 274.170 -283.510 274.340 -281.425 ;
        RECT 275.150 -283.510 275.320 -281.425 ;
        RECT 276.130 -281.675 280.565 -281.425 ;
        RECT 281.380 -281.615 281.605 -280.985 ;
        RECT 282.355 -281.600 282.580 -280.985 ;
        RECT 276.130 -283.510 276.300 -281.675 ;
        RECT 277.215 -282.505 277.385 -281.675 ;
        RECT 278.195 -282.505 278.365 -281.675 ;
        RECT 279.175 -282.505 279.345 -281.675 ;
        RECT 280.155 -282.505 280.325 -281.675 ;
        RECT 281.405 -284.565 281.575 -281.615 ;
        RECT 282.385 -284.565 282.555 -281.600 ;
        RECT 284.465 -281.605 284.690 -280.985 ;
        RECT 285.560 -281.020 285.870 -280.950 ;
        RECT 286.700 -281.050 290.100 -280.465 ;
        RECT 291.350 -280.890 291.540 -280.415 ;
        RECT 292.335 -280.880 292.525 -280.095 ;
        RECT 286.700 -281.080 287.190 -281.050 ;
        RECT 284.500 -284.565 284.670 -281.605 ;
        RECT 291.365 -283.355 291.535 -280.890 ;
        RECT 292.345 -283.355 292.515 -280.880 ;
        RECT 295.295 -280.995 295.545 -280.095 ;
        RECT 295.925 -280.980 296.175 -280.095 ;
        RECT 297.080 -280.905 297.295 -280.095 ;
        RECT 298.065 -280.325 328.445 -280.095 ;
        RECT 333.285 -280.085 335.310 -279.765 ;
        RECT 330.470 -280.135 330.960 -280.120 ;
        RECT 333.285 -280.135 333.870 -280.085 ;
        RECT 298.065 -280.360 328.965 -280.325 ;
        RECT 329.330 -280.360 329.640 -280.220 ;
        RECT 298.065 -280.405 329.640 -280.360 ;
        RECT 298.065 -280.895 298.280 -280.405 ;
        RECT 295.320 -283.355 295.490 -280.995 ;
        RECT 295.970 -283.355 296.140 -280.980 ;
        RECT 297.110 -282.355 297.280 -280.905 ;
        RECT 298.090 -282.355 298.260 -280.895 ;
        RECT 286.735 -291.040 288.745 -290.710 ;
        RECT 256.910 -292.855 260.070 -292.245 ;
        RECT 246.610 -296.245 246.780 -294.915 ;
        RECT 247.590 -296.245 247.760 -294.915 ;
        RECT 248.570 -296.245 248.740 -294.915 ;
        RECT 249.550 -296.245 249.720 -294.915 ;
        RECT 246.370 -296.740 249.960 -296.245 ;
        RECT 247.280 -297.690 248.140 -296.740 ;
        RECT 251.475 -297.145 251.645 -295.060 ;
        RECT 252.455 -297.145 252.625 -295.060 ;
        RECT 253.435 -296.895 253.605 -295.060 ;
        RECT 254.520 -296.895 254.690 -296.065 ;
        RECT 255.500 -296.895 255.670 -296.065 ;
        RECT 256.480 -296.895 256.650 -296.065 ;
        RECT 257.460 -296.895 257.630 -296.065 ;
        RECT 253.435 -297.145 257.870 -296.895 ;
        RECT 251.425 -297.390 257.870 -297.145 ;
        RECT 251.425 -297.460 253.635 -297.390 ;
        RECT 251.420 -297.605 253.635 -297.460 ;
        RECT 251.420 -297.690 254.510 -297.605 ;
        RECT 246.430 -297.860 256.985 -297.690 ;
        RECT 259.460 -297.835 260.070 -292.855 ;
        RECT 274.260 -295.920 274.430 -294.590 ;
        RECT 275.240 -295.920 275.410 -294.590 ;
        RECT 276.220 -295.920 276.390 -294.590 ;
        RECT 277.200 -295.920 277.370 -294.590 ;
        RECT 274.020 -296.415 277.610 -295.920 ;
        RECT 274.930 -297.365 275.790 -296.415 ;
        RECT 279.125 -296.820 279.295 -294.735 ;
        RECT 280.105 -296.820 280.275 -294.735 ;
        RECT 281.085 -296.570 281.255 -294.735 ;
        RECT 282.170 -296.570 282.340 -295.740 ;
        RECT 283.150 -296.570 283.320 -295.740 ;
        RECT 284.130 -296.570 284.300 -295.740 ;
        RECT 285.110 -296.570 285.280 -295.740 ;
        RECT 281.085 -296.820 285.520 -296.570 ;
        RECT 279.075 -297.065 285.520 -296.820 ;
        RECT 279.075 -297.135 281.285 -297.065 ;
        RECT 279.070 -297.280 281.285 -297.135 ;
        RECT 279.070 -297.365 282.160 -297.280 ;
        RECT 242.425 -298.190 256.985 -297.860 ;
        RECT 257.760 -298.065 258.155 -297.910 ;
        RECT 246.430 -298.245 256.985 -298.190 ;
        RECT 257.260 -298.245 258.155 -298.065 ;
        RECT 230.100 -298.335 231.230 -298.300 ;
        RECT 214.695 -298.475 215.390 -298.335 ;
        RECT 230.285 -298.370 231.230 -298.335 ;
        RECT 235.320 -298.420 239.165 -298.300 ;
        RECT 228.090 -298.615 230.300 -298.540 ;
        RECT 228.090 -298.860 234.535 -298.615 ;
        RECT 212.495 -301.960 212.665 -299.000 ;
        RECT 228.140 -300.945 228.310 -298.860 ;
        RECT 229.120 -300.945 229.290 -298.860 ;
        RECT 230.100 -299.110 234.535 -298.860 ;
        RECT 235.350 -299.050 235.575 -298.420 ;
        RECT 236.325 -299.035 236.550 -298.420 ;
        RECT 230.100 -300.945 230.270 -299.110 ;
        RECT 231.185 -299.940 231.355 -299.110 ;
        RECT 232.165 -299.940 232.335 -299.110 ;
        RECT 233.145 -299.940 233.315 -299.110 ;
        RECT 234.125 -299.940 234.295 -299.110 ;
        RECT 235.375 -302.000 235.545 -299.050 ;
        RECT 236.355 -302.000 236.525 -299.035 ;
        RECT 238.435 -299.040 238.660 -298.420 ;
        RECT 246.430 -298.455 258.155 -298.245 ;
        RECT 248.440 -298.490 249.570 -298.455 ;
        RECT 248.625 -298.525 249.570 -298.490 ;
        RECT 253.660 -298.480 258.155 -298.455 ;
        RECT 253.660 -298.575 257.505 -298.480 ;
        RECT 246.430 -298.770 248.640 -298.695 ;
        RECT 246.430 -299.015 252.875 -298.770 ;
        RECT 238.470 -302.000 238.640 -299.040 ;
        RECT 246.480 -301.100 246.650 -299.015 ;
        RECT 247.460 -301.100 247.630 -299.015 ;
        RECT 248.440 -299.265 252.875 -299.015 ;
        RECT 253.690 -299.205 253.915 -298.575 ;
        RECT 254.665 -299.190 254.890 -298.575 ;
        RECT 248.440 -301.100 248.610 -299.265 ;
        RECT 249.525 -300.095 249.695 -299.265 ;
        RECT 250.505 -300.095 250.675 -299.265 ;
        RECT 251.485 -300.095 251.655 -299.265 ;
        RECT 252.465 -300.095 252.635 -299.265 ;
        RECT 253.715 -302.155 253.885 -299.205 ;
        RECT 254.695 -302.155 254.865 -299.190 ;
        RECT 256.775 -299.195 257.000 -298.575 ;
        RECT 257.760 -298.605 258.155 -298.480 ;
        RECT 259.010 -298.530 260.070 -297.835 ;
        RECT 274.080 -297.920 284.635 -297.365 ;
        RECT 286.735 -297.545 287.065 -291.040 ;
        RECT 274.080 -298.130 285.155 -297.920 ;
        RECT 286.650 -298.110 287.070 -297.545 ;
        RECT 288.415 -297.690 288.745 -291.040 ;
        RECT 302.900 -292.075 303.510 -280.405 ;
        RECT 317.890 -280.535 329.640 -280.405 ;
        RECT 319.900 -280.570 321.030 -280.535 ;
        RECT 320.085 -280.605 321.030 -280.570 ;
        RECT 325.120 -280.620 329.640 -280.535 ;
        RECT 325.120 -280.655 328.965 -280.620 ;
        RECT 317.890 -280.850 320.100 -280.775 ;
        RECT 317.890 -281.095 324.335 -280.850 ;
        RECT 317.940 -283.180 318.110 -281.095 ;
        RECT 318.920 -283.180 319.090 -281.095 ;
        RECT 319.900 -281.345 324.335 -281.095 ;
        RECT 325.150 -281.285 325.375 -280.655 ;
        RECT 326.125 -281.270 326.350 -280.655 ;
        RECT 319.900 -283.180 320.070 -281.345 ;
        RECT 320.985 -282.175 321.155 -281.345 ;
        RECT 321.965 -282.175 322.135 -281.345 ;
        RECT 322.945 -282.175 323.115 -281.345 ;
        RECT 323.925 -282.175 324.095 -281.345 ;
        RECT 325.175 -284.235 325.345 -281.285 ;
        RECT 326.155 -284.235 326.325 -281.270 ;
        RECT 328.235 -281.275 328.460 -280.655 ;
        RECT 329.330 -280.690 329.640 -280.620 ;
        RECT 330.470 -280.720 333.870 -280.135 ;
        RECT 335.120 -280.560 335.310 -280.085 ;
        RECT 336.105 -280.550 336.295 -279.765 ;
        RECT 330.470 -280.750 330.960 -280.720 ;
        RECT 328.270 -284.235 328.440 -281.275 ;
        RECT 335.135 -283.025 335.305 -280.560 ;
        RECT 336.115 -283.025 336.285 -280.550 ;
        RECT 339.065 -280.665 339.315 -279.765 ;
        RECT 339.695 -280.650 339.945 -279.765 ;
        RECT 340.850 -280.575 341.065 -279.765 ;
        RECT 341.810 -279.935 374.210 -279.765 ;
        RECT 341.835 -280.565 342.050 -279.935 ;
        RECT 339.090 -283.025 339.260 -280.665 ;
        RECT 339.740 -283.025 339.910 -280.650 ;
        RECT 340.880 -282.025 341.050 -280.575 ;
        RECT 341.860 -282.025 342.030 -280.565 ;
        RECT 330.505 -290.710 332.515 -290.380 ;
        RECT 302.900 -292.685 306.060 -292.075 ;
        RECT 292.600 -296.075 292.770 -294.745 ;
        RECT 293.580 -296.075 293.750 -294.745 ;
        RECT 294.560 -296.075 294.730 -294.745 ;
        RECT 295.540 -296.075 295.710 -294.745 ;
        RECT 292.360 -296.570 295.950 -296.075 ;
        RECT 293.270 -297.520 294.130 -296.570 ;
        RECT 297.465 -296.975 297.635 -294.890 ;
        RECT 298.445 -296.975 298.615 -294.890 ;
        RECT 299.425 -296.725 299.595 -294.890 ;
        RECT 300.510 -296.725 300.680 -295.895 ;
        RECT 301.490 -296.725 301.660 -295.895 ;
        RECT 302.470 -296.725 302.640 -295.895 ;
        RECT 303.450 -296.725 303.620 -295.895 ;
        RECT 299.425 -296.975 303.860 -296.725 ;
        RECT 297.415 -297.220 303.860 -296.975 ;
        RECT 297.415 -297.290 299.625 -297.220 ;
        RECT 297.410 -297.435 299.625 -297.290 ;
        RECT 297.410 -297.520 300.500 -297.435 ;
        RECT 292.420 -297.690 302.975 -297.520 ;
        RECT 305.450 -297.665 306.060 -292.685 ;
        RECT 318.030 -295.590 318.200 -294.260 ;
        RECT 319.010 -295.590 319.180 -294.260 ;
        RECT 319.990 -295.590 320.160 -294.260 ;
        RECT 320.970 -295.590 321.140 -294.260 ;
        RECT 317.790 -296.085 321.380 -295.590 ;
        RECT 318.700 -297.035 319.560 -296.085 ;
        RECT 322.895 -296.490 323.065 -294.405 ;
        RECT 323.875 -296.490 324.045 -294.405 ;
        RECT 324.855 -296.240 325.025 -294.405 ;
        RECT 325.940 -296.240 326.110 -295.410 ;
        RECT 326.920 -296.240 327.090 -295.410 ;
        RECT 327.900 -296.240 328.070 -295.410 ;
        RECT 328.880 -296.240 329.050 -295.410 ;
        RECT 324.855 -296.490 329.290 -296.240 ;
        RECT 322.845 -296.735 329.290 -296.490 ;
        RECT 322.845 -296.805 325.055 -296.735 ;
        RECT 322.840 -296.950 325.055 -296.805 ;
        RECT 322.840 -297.035 325.930 -296.950 ;
        RECT 288.415 -298.020 302.975 -297.690 ;
        RECT 303.750 -297.895 304.145 -297.740 ;
        RECT 292.420 -298.075 302.975 -298.020 ;
        RECT 303.250 -298.075 304.145 -297.895 ;
        RECT 276.090 -298.165 277.220 -298.130 ;
        RECT 276.275 -298.200 277.220 -298.165 ;
        RECT 281.310 -298.250 285.155 -298.130 ;
        RECT 274.080 -298.445 276.290 -298.370 ;
        RECT 259.010 -298.670 259.705 -298.530 ;
        RECT 274.080 -298.690 280.525 -298.445 ;
        RECT 256.810 -302.155 256.980 -299.195 ;
        RECT 274.130 -300.775 274.300 -298.690 ;
        RECT 275.110 -300.775 275.280 -298.690 ;
        RECT 276.090 -298.940 280.525 -298.690 ;
        RECT 281.340 -298.880 281.565 -298.250 ;
        RECT 282.315 -298.865 282.540 -298.250 ;
        RECT 276.090 -300.775 276.260 -298.940 ;
        RECT 277.175 -299.770 277.345 -298.940 ;
        RECT 278.155 -299.770 278.325 -298.940 ;
        RECT 279.135 -299.770 279.305 -298.940 ;
        RECT 280.115 -299.770 280.285 -298.940 ;
        RECT 281.365 -301.830 281.535 -298.880 ;
        RECT 282.345 -301.830 282.515 -298.865 ;
        RECT 284.425 -298.870 284.650 -298.250 ;
        RECT 292.420 -298.285 304.145 -298.075 ;
        RECT 294.430 -298.320 295.560 -298.285 ;
        RECT 294.615 -298.355 295.560 -298.320 ;
        RECT 299.650 -298.310 304.145 -298.285 ;
        RECT 299.650 -298.405 303.495 -298.310 ;
        RECT 292.420 -298.600 294.630 -298.525 ;
        RECT 292.420 -298.845 298.865 -298.600 ;
        RECT 284.460 -301.830 284.630 -298.870 ;
        RECT 292.470 -300.930 292.640 -298.845 ;
        RECT 293.450 -300.930 293.620 -298.845 ;
        RECT 294.430 -299.095 298.865 -298.845 ;
        RECT 299.680 -299.035 299.905 -298.405 ;
        RECT 300.655 -299.020 300.880 -298.405 ;
        RECT 294.430 -300.930 294.600 -299.095 ;
        RECT 295.515 -299.925 295.685 -299.095 ;
        RECT 296.495 -299.925 296.665 -299.095 ;
        RECT 297.475 -299.925 297.645 -299.095 ;
        RECT 298.455 -299.925 298.625 -299.095 ;
        RECT 299.705 -301.985 299.875 -299.035 ;
        RECT 300.685 -301.985 300.855 -299.020 ;
        RECT 302.765 -299.025 302.990 -298.405 ;
        RECT 303.750 -298.435 304.145 -298.310 ;
        RECT 305.000 -298.360 306.060 -297.665 ;
        RECT 317.850 -297.590 328.405 -297.035 ;
        RECT 330.505 -297.215 330.835 -290.710 ;
        RECT 317.850 -297.800 328.925 -297.590 ;
        RECT 330.420 -297.780 330.840 -297.215 ;
        RECT 332.185 -297.360 332.515 -290.710 ;
        RECT 346.670 -291.745 347.280 -279.935 ;
        RECT 363.655 -280.240 374.210 -279.935 ;
        RECT 379.050 -280.000 381.075 -279.680 ;
        RECT 376.235 -280.050 376.725 -280.035 ;
        RECT 379.050 -280.050 379.635 -280.000 ;
        RECT 363.655 -280.275 374.730 -280.240 ;
        RECT 375.095 -280.275 375.405 -280.135 ;
        RECT 363.655 -280.450 375.405 -280.275 ;
        RECT 365.665 -280.485 366.795 -280.450 ;
        RECT 365.850 -280.520 366.795 -280.485 ;
        RECT 370.885 -280.535 375.405 -280.450 ;
        RECT 370.885 -280.570 374.730 -280.535 ;
        RECT 363.655 -280.765 365.865 -280.690 ;
        RECT 363.655 -281.010 370.100 -280.765 ;
        RECT 363.705 -283.095 363.875 -281.010 ;
        RECT 364.685 -283.095 364.855 -281.010 ;
        RECT 365.665 -281.260 370.100 -281.010 ;
        RECT 370.915 -281.200 371.140 -280.570 ;
        RECT 371.890 -281.185 372.115 -280.570 ;
        RECT 365.665 -283.095 365.835 -281.260 ;
        RECT 366.750 -282.090 366.920 -281.260 ;
        RECT 367.730 -282.090 367.900 -281.260 ;
        RECT 368.710 -282.090 368.880 -281.260 ;
        RECT 369.690 -282.090 369.860 -281.260 ;
        RECT 370.940 -284.150 371.110 -281.200 ;
        RECT 371.920 -284.150 372.090 -281.185 ;
        RECT 374.000 -281.190 374.225 -280.570 ;
        RECT 375.095 -280.605 375.405 -280.535 ;
        RECT 376.235 -280.635 379.635 -280.050 ;
        RECT 380.885 -280.475 381.075 -280.000 ;
        RECT 381.870 -280.465 382.060 -279.680 ;
        RECT 376.235 -280.665 376.725 -280.635 ;
        RECT 374.035 -284.150 374.205 -281.190 ;
        RECT 380.900 -282.940 381.070 -280.475 ;
        RECT 381.880 -282.940 382.050 -280.465 ;
        RECT 384.830 -280.580 385.080 -279.680 ;
        RECT 385.460 -280.565 385.710 -279.680 ;
        RECT 386.615 -280.490 386.830 -279.680 ;
        RECT 387.600 -279.980 421.030 -279.680 ;
        RECT 425.870 -279.810 427.895 -279.490 ;
        RECT 423.055 -279.860 423.545 -279.845 ;
        RECT 425.870 -279.860 426.455 -279.810 ;
        RECT 387.600 -280.480 387.815 -279.980 ;
        RECT 384.855 -282.940 385.025 -280.580 ;
        RECT 385.505 -282.940 385.675 -280.565 ;
        RECT 386.645 -281.940 386.815 -280.490 ;
        RECT 387.625 -281.940 387.795 -280.480 ;
        RECT 376.270 -290.625 378.280 -290.295 ;
        RECT 346.670 -292.355 349.830 -291.745 ;
        RECT 336.370 -295.745 336.540 -294.415 ;
        RECT 337.350 -295.745 337.520 -294.415 ;
        RECT 338.330 -295.745 338.500 -294.415 ;
        RECT 339.310 -295.745 339.480 -294.415 ;
        RECT 336.130 -296.240 339.720 -295.745 ;
        RECT 337.040 -297.190 337.900 -296.240 ;
        RECT 341.235 -296.645 341.405 -294.560 ;
        RECT 342.215 -296.645 342.385 -294.560 ;
        RECT 343.195 -296.395 343.365 -294.560 ;
        RECT 344.280 -296.395 344.450 -295.565 ;
        RECT 345.260 -296.395 345.430 -295.565 ;
        RECT 346.240 -296.395 346.410 -295.565 ;
        RECT 347.220 -296.395 347.390 -295.565 ;
        RECT 343.195 -296.645 347.630 -296.395 ;
        RECT 341.185 -296.890 347.630 -296.645 ;
        RECT 341.185 -296.960 343.395 -296.890 ;
        RECT 341.180 -297.105 343.395 -296.960 ;
        RECT 341.180 -297.190 344.270 -297.105 ;
        RECT 336.190 -297.360 346.745 -297.190 ;
        RECT 349.220 -297.335 349.830 -292.355 ;
        RECT 363.795 -295.505 363.965 -294.175 ;
        RECT 364.775 -295.505 364.945 -294.175 ;
        RECT 365.755 -295.505 365.925 -294.175 ;
        RECT 366.735 -295.505 366.905 -294.175 ;
        RECT 363.555 -296.000 367.145 -295.505 ;
        RECT 364.465 -296.950 365.325 -296.000 ;
        RECT 368.660 -296.405 368.830 -294.320 ;
        RECT 369.640 -296.405 369.810 -294.320 ;
        RECT 370.620 -296.155 370.790 -294.320 ;
        RECT 371.705 -296.155 371.875 -295.325 ;
        RECT 372.685 -296.155 372.855 -295.325 ;
        RECT 373.665 -296.155 373.835 -295.325 ;
        RECT 374.645 -296.155 374.815 -295.325 ;
        RECT 370.620 -296.405 375.055 -296.155 ;
        RECT 368.610 -296.650 375.055 -296.405 ;
        RECT 368.610 -296.720 370.820 -296.650 ;
        RECT 368.605 -296.865 370.820 -296.720 ;
        RECT 368.605 -296.950 371.695 -296.865 ;
        RECT 332.185 -297.690 346.745 -297.360 ;
        RECT 347.520 -297.565 347.915 -297.410 ;
        RECT 336.190 -297.745 346.745 -297.690 ;
        RECT 347.020 -297.745 347.915 -297.565 ;
        RECT 319.860 -297.835 320.990 -297.800 ;
        RECT 320.045 -297.870 320.990 -297.835 ;
        RECT 325.080 -297.920 328.925 -297.800 ;
        RECT 317.850 -298.115 320.060 -298.040 ;
        RECT 317.850 -298.360 324.295 -298.115 ;
        RECT 305.000 -298.500 305.695 -298.360 ;
        RECT 302.800 -301.985 302.970 -299.025 ;
        RECT 317.900 -300.445 318.070 -298.360 ;
        RECT 318.880 -300.445 319.050 -298.360 ;
        RECT 319.860 -298.610 324.295 -298.360 ;
        RECT 325.110 -298.550 325.335 -297.920 ;
        RECT 326.085 -298.535 326.310 -297.920 ;
        RECT 319.860 -300.445 320.030 -298.610 ;
        RECT 320.945 -299.440 321.115 -298.610 ;
        RECT 321.925 -299.440 322.095 -298.610 ;
        RECT 322.905 -299.440 323.075 -298.610 ;
        RECT 323.885 -299.440 324.055 -298.610 ;
        RECT 325.135 -301.500 325.305 -298.550 ;
        RECT 326.115 -301.500 326.285 -298.535 ;
        RECT 328.195 -298.540 328.420 -297.920 ;
        RECT 336.190 -297.955 347.915 -297.745 ;
        RECT 338.200 -297.990 339.330 -297.955 ;
        RECT 338.385 -298.025 339.330 -297.990 ;
        RECT 343.420 -297.980 347.915 -297.955 ;
        RECT 343.420 -298.075 347.265 -297.980 ;
        RECT 336.190 -298.270 338.400 -298.195 ;
        RECT 336.190 -298.515 342.635 -298.270 ;
        RECT 328.230 -301.500 328.400 -298.540 ;
        RECT 336.240 -300.600 336.410 -298.515 ;
        RECT 337.220 -300.600 337.390 -298.515 ;
        RECT 338.200 -298.765 342.635 -298.515 ;
        RECT 343.450 -298.705 343.675 -298.075 ;
        RECT 344.425 -298.690 344.650 -298.075 ;
        RECT 338.200 -300.600 338.370 -298.765 ;
        RECT 339.285 -299.595 339.455 -298.765 ;
        RECT 340.265 -299.595 340.435 -298.765 ;
        RECT 341.245 -299.595 341.415 -298.765 ;
        RECT 342.225 -299.595 342.395 -298.765 ;
        RECT 343.475 -301.655 343.645 -298.705 ;
        RECT 344.455 -301.655 344.625 -298.690 ;
        RECT 346.535 -298.695 346.760 -298.075 ;
        RECT 347.520 -298.105 347.915 -297.980 ;
        RECT 348.770 -298.030 349.830 -297.335 ;
        RECT 363.615 -297.505 374.170 -296.950 ;
        RECT 376.270 -297.130 376.600 -290.625 ;
        RECT 363.615 -297.715 374.690 -297.505 ;
        RECT 376.185 -297.695 376.605 -297.130 ;
        RECT 377.950 -297.275 378.280 -290.625 ;
        RECT 392.435 -291.660 393.045 -279.980 ;
        RECT 410.475 -280.050 421.030 -279.980 ;
        RECT 410.475 -280.085 421.550 -280.050 ;
        RECT 421.915 -280.085 422.225 -279.945 ;
        RECT 410.475 -280.260 422.225 -280.085 ;
        RECT 412.485 -280.295 413.615 -280.260 ;
        RECT 412.670 -280.330 413.615 -280.295 ;
        RECT 417.705 -280.345 422.225 -280.260 ;
        RECT 417.705 -280.380 421.550 -280.345 ;
        RECT 410.475 -280.575 412.685 -280.500 ;
        RECT 410.475 -280.820 416.920 -280.575 ;
        RECT 410.525 -282.905 410.695 -280.820 ;
        RECT 411.505 -282.905 411.675 -280.820 ;
        RECT 412.485 -281.070 416.920 -280.820 ;
        RECT 417.735 -281.010 417.960 -280.380 ;
        RECT 418.710 -280.995 418.935 -280.380 ;
        RECT 412.485 -282.905 412.655 -281.070 ;
        RECT 413.570 -281.900 413.740 -281.070 ;
        RECT 414.550 -281.900 414.720 -281.070 ;
        RECT 415.530 -281.900 415.700 -281.070 ;
        RECT 416.510 -281.900 416.680 -281.070 ;
        RECT 417.760 -283.960 417.930 -281.010 ;
        RECT 418.740 -283.960 418.910 -280.995 ;
        RECT 420.820 -281.000 421.045 -280.380 ;
        RECT 421.915 -280.415 422.225 -280.345 ;
        RECT 423.055 -280.445 426.455 -279.860 ;
        RECT 427.705 -280.285 427.895 -279.810 ;
        RECT 428.690 -280.275 428.880 -279.490 ;
        RECT 423.055 -280.475 423.545 -280.445 ;
        RECT 420.855 -283.960 421.025 -281.000 ;
        RECT 427.720 -282.750 427.890 -280.285 ;
        RECT 428.700 -282.750 428.870 -280.275 ;
        RECT 431.650 -280.390 431.900 -279.490 ;
        RECT 432.280 -280.375 432.530 -279.490 ;
        RECT 433.435 -280.300 433.650 -279.490 ;
        RECT 434.420 -280.290 434.635 -279.490 ;
        RECT 431.675 -282.750 431.845 -280.390 ;
        RECT 432.325 -282.750 432.495 -280.375 ;
        RECT 433.465 -281.750 433.635 -280.300 ;
        RECT 434.445 -281.750 434.615 -280.290 ;
        RECT 423.090 -290.435 425.100 -290.105 ;
        RECT 392.435 -292.270 395.595 -291.660 ;
        RECT 382.135 -295.660 382.305 -294.330 ;
        RECT 383.115 -295.660 383.285 -294.330 ;
        RECT 384.095 -295.660 384.265 -294.330 ;
        RECT 385.075 -295.660 385.245 -294.330 ;
        RECT 381.895 -296.155 385.485 -295.660 ;
        RECT 382.805 -297.105 383.665 -296.155 ;
        RECT 387.000 -296.560 387.170 -294.475 ;
        RECT 387.980 -296.560 388.150 -294.475 ;
        RECT 388.960 -296.310 389.130 -294.475 ;
        RECT 390.045 -296.310 390.215 -295.480 ;
        RECT 391.025 -296.310 391.195 -295.480 ;
        RECT 392.005 -296.310 392.175 -295.480 ;
        RECT 392.985 -296.310 393.155 -295.480 ;
        RECT 388.960 -296.560 393.395 -296.310 ;
        RECT 386.950 -296.805 393.395 -296.560 ;
        RECT 386.950 -296.875 389.160 -296.805 ;
        RECT 386.945 -297.020 389.160 -296.875 ;
        RECT 386.945 -297.105 390.035 -297.020 ;
        RECT 381.955 -297.275 392.510 -297.105 ;
        RECT 394.985 -297.250 395.595 -292.270 ;
        RECT 410.615 -295.315 410.785 -293.985 ;
        RECT 411.595 -295.315 411.765 -293.985 ;
        RECT 412.575 -295.315 412.745 -293.985 ;
        RECT 413.555 -295.315 413.725 -293.985 ;
        RECT 410.375 -295.810 413.965 -295.315 ;
        RECT 411.285 -296.760 412.145 -295.810 ;
        RECT 415.480 -296.215 415.650 -294.130 ;
        RECT 416.460 -296.215 416.630 -294.130 ;
        RECT 417.440 -295.965 417.610 -294.130 ;
        RECT 418.525 -295.965 418.695 -295.135 ;
        RECT 419.505 -295.965 419.675 -295.135 ;
        RECT 420.485 -295.965 420.655 -295.135 ;
        RECT 421.465 -295.965 421.635 -295.135 ;
        RECT 417.440 -296.215 421.875 -295.965 ;
        RECT 415.430 -296.460 421.875 -296.215 ;
        RECT 415.430 -296.530 417.640 -296.460 ;
        RECT 415.425 -296.675 417.640 -296.530 ;
        RECT 415.425 -296.760 418.515 -296.675 ;
        RECT 377.950 -297.605 392.510 -297.275 ;
        RECT 393.285 -297.480 393.680 -297.325 ;
        RECT 381.955 -297.660 392.510 -297.605 ;
        RECT 392.785 -297.660 393.680 -297.480 ;
        RECT 365.625 -297.750 366.755 -297.715 ;
        RECT 365.810 -297.785 366.755 -297.750 ;
        RECT 370.845 -297.835 374.690 -297.715 ;
        RECT 363.615 -298.030 365.825 -297.955 ;
        RECT 348.770 -298.170 349.465 -298.030 ;
        RECT 363.615 -298.275 370.060 -298.030 ;
        RECT 346.570 -301.655 346.740 -298.695 ;
        RECT 363.665 -300.360 363.835 -298.275 ;
        RECT 364.645 -300.360 364.815 -298.275 ;
        RECT 365.625 -298.525 370.060 -298.275 ;
        RECT 370.875 -298.465 371.100 -297.835 ;
        RECT 371.850 -298.450 372.075 -297.835 ;
        RECT 365.625 -300.360 365.795 -298.525 ;
        RECT 366.710 -299.355 366.880 -298.525 ;
        RECT 367.690 -299.355 367.860 -298.525 ;
        RECT 368.670 -299.355 368.840 -298.525 ;
        RECT 369.650 -299.355 369.820 -298.525 ;
        RECT 370.900 -301.415 371.070 -298.465 ;
        RECT 371.880 -301.415 372.050 -298.450 ;
        RECT 373.960 -298.455 374.185 -297.835 ;
        RECT 381.955 -297.870 393.680 -297.660 ;
        RECT 383.965 -297.905 385.095 -297.870 ;
        RECT 384.150 -297.940 385.095 -297.905 ;
        RECT 389.185 -297.895 393.680 -297.870 ;
        RECT 389.185 -297.990 393.030 -297.895 ;
        RECT 381.955 -298.185 384.165 -298.110 ;
        RECT 381.955 -298.430 388.400 -298.185 ;
        RECT 373.995 -301.415 374.165 -298.455 ;
        RECT 382.005 -300.515 382.175 -298.430 ;
        RECT 382.985 -300.515 383.155 -298.430 ;
        RECT 383.965 -298.680 388.400 -298.430 ;
        RECT 389.215 -298.620 389.440 -297.990 ;
        RECT 390.190 -298.605 390.415 -297.990 ;
        RECT 383.965 -300.515 384.135 -298.680 ;
        RECT 385.050 -299.510 385.220 -298.680 ;
        RECT 386.030 -299.510 386.200 -298.680 ;
        RECT 387.010 -299.510 387.180 -298.680 ;
        RECT 387.990 -299.510 388.160 -298.680 ;
        RECT 389.240 -301.570 389.410 -298.620 ;
        RECT 390.220 -301.570 390.390 -298.605 ;
        RECT 392.300 -298.610 392.525 -297.990 ;
        RECT 393.285 -298.020 393.680 -297.895 ;
        RECT 394.535 -297.945 395.595 -297.250 ;
        RECT 410.435 -297.315 420.990 -296.760 ;
        RECT 423.090 -296.940 423.420 -290.435 ;
        RECT 410.435 -297.525 421.510 -297.315 ;
        RECT 423.005 -297.505 423.425 -296.940 ;
        RECT 424.770 -297.085 425.100 -290.435 ;
        RECT 439.255 -291.470 439.865 -279.485 ;
        RECT 439.255 -292.080 442.415 -291.470 ;
        RECT 428.955 -295.470 429.125 -294.140 ;
        RECT 429.935 -295.470 430.105 -294.140 ;
        RECT 430.915 -295.470 431.085 -294.140 ;
        RECT 431.895 -295.470 432.065 -294.140 ;
        RECT 428.715 -295.965 432.305 -295.470 ;
        RECT 429.625 -296.915 430.485 -295.965 ;
        RECT 433.820 -296.370 433.990 -294.285 ;
        RECT 434.800 -296.370 434.970 -294.285 ;
        RECT 435.780 -296.120 435.950 -294.285 ;
        RECT 436.865 -296.120 437.035 -295.290 ;
        RECT 437.845 -296.120 438.015 -295.290 ;
        RECT 438.825 -296.120 438.995 -295.290 ;
        RECT 439.805 -296.120 439.975 -295.290 ;
        RECT 435.780 -296.370 440.215 -296.120 ;
        RECT 433.770 -296.615 440.215 -296.370 ;
        RECT 433.770 -296.685 435.980 -296.615 ;
        RECT 433.765 -296.830 435.980 -296.685 ;
        RECT 433.765 -296.915 436.855 -296.830 ;
        RECT 428.775 -297.085 439.330 -296.915 ;
        RECT 441.805 -297.060 442.415 -292.080 ;
        RECT 424.770 -297.415 439.330 -297.085 ;
        RECT 440.105 -297.290 440.500 -297.135 ;
        RECT 428.775 -297.470 439.330 -297.415 ;
        RECT 439.605 -297.470 440.500 -297.290 ;
        RECT 412.445 -297.560 413.575 -297.525 ;
        RECT 412.630 -297.595 413.575 -297.560 ;
        RECT 417.665 -297.645 421.510 -297.525 ;
        RECT 410.435 -297.840 412.645 -297.765 ;
        RECT 394.535 -298.085 395.230 -297.945 ;
        RECT 410.435 -298.085 416.880 -297.840 ;
        RECT 392.335 -301.570 392.505 -298.610 ;
        RECT 410.485 -300.170 410.655 -298.085 ;
        RECT 411.465 -300.170 411.635 -298.085 ;
        RECT 412.445 -298.335 416.880 -298.085 ;
        RECT 417.695 -298.275 417.920 -297.645 ;
        RECT 418.670 -298.260 418.895 -297.645 ;
        RECT 412.445 -300.170 412.615 -298.335 ;
        RECT 413.530 -299.165 413.700 -298.335 ;
        RECT 414.510 -299.165 414.680 -298.335 ;
        RECT 415.490 -299.165 415.660 -298.335 ;
        RECT 416.470 -299.165 416.640 -298.335 ;
        RECT 417.720 -301.225 417.890 -298.275 ;
        RECT 418.700 -301.225 418.870 -298.260 ;
        RECT 420.780 -298.265 421.005 -297.645 ;
        RECT 428.775 -297.680 440.500 -297.470 ;
        RECT 430.785 -297.715 431.915 -297.680 ;
        RECT 430.970 -297.750 431.915 -297.715 ;
        RECT 436.005 -297.705 440.500 -297.680 ;
        RECT 436.005 -297.800 439.850 -297.705 ;
        RECT 428.775 -297.995 430.985 -297.920 ;
        RECT 428.775 -298.240 435.220 -297.995 ;
        RECT 420.815 -301.225 420.985 -298.265 ;
        RECT 428.825 -300.325 428.995 -298.240 ;
        RECT 429.805 -300.325 429.975 -298.240 ;
        RECT 430.785 -298.490 435.220 -298.240 ;
        RECT 436.035 -298.430 436.260 -297.800 ;
        RECT 437.010 -298.415 437.235 -297.800 ;
        RECT 430.785 -300.325 430.955 -298.490 ;
        RECT 431.870 -299.320 432.040 -298.490 ;
        RECT 432.850 -299.320 433.020 -298.490 ;
        RECT 433.830 -299.320 434.000 -298.490 ;
        RECT 434.810 -299.320 434.980 -298.490 ;
        RECT 436.060 -301.380 436.230 -298.430 ;
        RECT 437.040 -301.380 437.210 -298.415 ;
        RECT 439.120 -298.420 439.345 -297.800 ;
        RECT 440.105 -297.830 440.500 -297.705 ;
        RECT 441.355 -297.755 442.415 -297.060 ;
        RECT 441.355 -297.895 442.050 -297.755 ;
        RECT 439.155 -301.380 439.325 -298.420 ;
        RECT 68.990 -309.860 78.000 -309.835 ;
        RECT 82.490 -309.860 90.355 -309.835 ;
        RECT 43.690 -310.755 43.920 -310.145 ;
        RECT 64.230 -310.175 90.355 -309.860 ;
        RECT 12.980 -311.290 15.945 -311.100 ;
        RECT 25.045 -311.290 28.010 -311.100 ;
        RECT 38.660 -311.290 43.920 -310.755 ;
        RECT -106.870 -311.465 -93.860 -311.420 ;
        RECT -30.665 -312.255 44.145 -311.290 ;
      LAYER met1 ;
        RECT -56.790 600.885 -55.835 601.640 ;
        RECT -56.665 600.090 -55.970 600.885 ;
        RECT -56.725 599.635 -55.910 600.090 ;
        RECT -54.645 599.335 -54.145 599.565 ;
        RECT -60.195 598.685 -57.195 598.915 ;
        RECT -54.645 598.355 -54.145 598.585 ;
        RECT -54.645 597.375 -54.145 597.605 ;
        RECT -60.195 596.570 -57.195 596.800 ;
        RECT -54.645 596.395 -54.145 596.625 ;
        RECT -60.195 595.590 -57.195 595.820 ;
        RECT -54.640 595.310 -53.140 595.540 ;
        RECT -58.135 594.340 -57.635 594.570 ;
        RECT -54.640 594.330 -53.140 594.560 ;
        RECT -40.565 593.975 -39.065 594.205 ;
        RECT -58.135 593.360 -57.635 593.590 ;
        RECT -54.640 593.350 -53.140 593.580 ;
        RECT -40.565 592.995 -39.065 593.225 ;
        RECT -58.135 592.380 -57.635 592.610 ;
        RECT -41.565 591.855 -39.065 592.085 ;
        RECT -58.135 591.400 -57.635 591.630 ;
        RECT -53.995 591.425 -52.995 591.655 ;
        RECT -41.565 591.205 -39.065 591.435 ;
        RECT -59.140 590.315 -57.640 590.545 ;
        RECT -53.995 590.445 -52.995 590.675 ;
        RECT -59.140 589.335 -57.640 589.565 ;
        RECT -53.995 589.465 -52.995 589.695 ;
        RECT -59.140 588.355 -57.640 588.585 ;
        RECT -53.995 588.485 -52.995 588.715 ;
        RECT -41.565 588.230 -39.065 588.460 ;
        RECT -41.565 587.250 -39.065 587.480 ;
        RECT -56.400 582.535 -55.715 583.015 ;
        RECT -39.370 582.585 -38.620 583.135 ;
        RECT -60.040 580.345 -57.040 580.575 ;
        RECT -60.040 578.230 -57.040 578.460 ;
        RECT -60.040 577.250 -57.040 577.480 ;
        RECT -56.270 576.935 -55.860 582.535 ;
        RECT -39.280 581.815 -38.800 582.585 ;
        RECT -39.310 581.445 -38.720 581.815 ;
        RECT -54.490 580.995 -53.990 581.225 ;
        RECT -37.225 581.035 -36.725 581.265 ;
        RECT -42.775 580.385 -39.775 580.615 ;
        RECT -54.490 580.015 -53.990 580.245 ;
        RECT -37.225 580.055 -36.725 580.285 ;
        RECT -54.490 579.035 -53.990 579.265 ;
        RECT -37.225 579.075 -36.725 579.305 ;
        RECT -54.490 578.055 -53.990 578.285 ;
        RECT -42.775 578.270 -39.775 578.500 ;
        RECT -37.225 578.095 -36.725 578.325 ;
        RECT -42.775 577.290 -39.775 577.520 ;
        RECT -54.485 576.970 -52.985 577.200 ;
        RECT -37.220 577.010 -35.720 577.240 ;
        RECT -57.980 576.000 -57.480 576.230 ;
        RECT -56.305 576.020 -55.655 576.935 ;
        RECT -54.485 575.990 -52.985 576.220 ;
        RECT -40.715 576.040 -40.215 576.270 ;
        RECT -37.220 576.030 -35.720 576.260 ;
        RECT -57.980 575.020 -57.480 575.250 ;
        RECT -54.485 575.010 -52.985 575.240 ;
        RECT -40.715 575.060 -40.215 575.290 ;
        RECT -37.220 575.050 -35.720 575.280 ;
        RECT -57.980 574.040 -57.480 574.270 ;
        RECT -40.715 574.080 -40.215 574.310 ;
        RECT -57.980 573.060 -57.480 573.290 ;
        RECT -53.840 573.085 -52.840 573.315 ;
        RECT -40.715 573.100 -40.215 573.330 ;
        RECT -36.575 573.125 -35.575 573.355 ;
        RECT -58.985 571.975 -57.485 572.205 ;
        RECT -53.840 572.105 -52.840 572.335 ;
        RECT -41.720 572.015 -40.220 572.245 ;
        RECT -36.575 572.145 -35.575 572.375 ;
        RECT -58.985 570.995 -57.485 571.225 ;
        RECT -53.840 571.125 -52.840 571.355 ;
        RECT -41.720 571.035 -40.220 571.265 ;
        RECT -36.575 571.165 -35.575 571.395 ;
        RECT -58.985 570.015 -57.485 570.245 ;
        RECT -53.840 570.145 -52.840 570.375 ;
        RECT -41.720 570.055 -40.220 570.285 ;
        RECT -36.575 570.185 -35.575 570.415 ;
        RECT -56.980 554.065 -56.025 554.820 ;
        RECT -56.855 553.270 -56.160 554.065 ;
        RECT -56.915 552.815 -56.100 553.270 ;
        RECT -54.835 552.515 -54.335 552.745 ;
        RECT -60.385 551.865 -57.385 552.095 ;
        RECT -54.835 551.535 -54.335 551.765 ;
        RECT -54.835 550.555 -54.335 550.785 ;
        RECT -60.385 549.750 -57.385 549.980 ;
        RECT -54.835 549.575 -54.335 549.805 ;
        RECT -60.385 548.770 -57.385 549.000 ;
        RECT -54.830 548.490 -53.330 548.720 ;
        RECT -58.325 547.520 -57.825 547.750 ;
        RECT -54.830 547.510 -53.330 547.740 ;
        RECT -40.755 547.155 -39.255 547.385 ;
        RECT -58.325 546.540 -57.825 546.770 ;
        RECT -54.830 546.530 -53.330 546.760 ;
        RECT -40.755 546.175 -39.255 546.405 ;
        RECT -58.325 545.560 -57.825 545.790 ;
        RECT -41.755 545.035 -39.255 545.265 ;
        RECT -58.325 544.580 -57.825 544.810 ;
        RECT -54.185 544.605 -53.185 544.835 ;
        RECT -41.755 544.385 -39.255 544.615 ;
        RECT -59.330 543.495 -57.830 543.725 ;
        RECT -54.185 543.625 -53.185 543.855 ;
        RECT -59.330 542.515 -57.830 542.745 ;
        RECT -54.185 542.645 -53.185 542.875 ;
        RECT -59.330 541.535 -57.830 541.765 ;
        RECT -54.185 541.665 -53.185 541.895 ;
        RECT -41.755 541.410 -39.255 541.640 ;
        RECT -41.755 540.430 -39.255 540.660 ;
        RECT -56.590 535.715 -55.905 536.195 ;
        RECT -39.560 535.765 -38.810 536.315 ;
        RECT -60.230 533.525 -57.230 533.755 ;
        RECT -60.230 531.410 -57.230 531.640 ;
        RECT -60.230 530.430 -57.230 530.660 ;
        RECT -56.460 530.115 -56.050 535.715 ;
        RECT -39.470 534.995 -38.990 535.765 ;
        RECT -39.500 534.625 -38.910 534.995 ;
        RECT -54.680 534.175 -54.180 534.405 ;
        RECT -37.415 534.215 -36.915 534.445 ;
        RECT -42.965 533.565 -39.965 533.795 ;
        RECT -54.680 533.195 -54.180 533.425 ;
        RECT -37.415 533.235 -36.915 533.465 ;
        RECT -54.680 532.215 -54.180 532.445 ;
        RECT -37.415 532.255 -36.915 532.485 ;
        RECT -54.680 531.235 -54.180 531.465 ;
        RECT -42.965 531.450 -39.965 531.680 ;
        RECT -37.415 531.275 -36.915 531.505 ;
        RECT -42.965 530.470 -39.965 530.700 ;
        RECT -54.675 530.150 -53.175 530.380 ;
        RECT -37.410 530.190 -35.910 530.420 ;
        RECT -58.170 529.180 -57.670 529.410 ;
        RECT -56.495 529.200 -55.845 530.115 ;
        RECT -54.675 529.170 -53.175 529.400 ;
        RECT -40.905 529.220 -40.405 529.450 ;
        RECT -37.410 529.210 -35.910 529.440 ;
        RECT -58.170 528.200 -57.670 528.430 ;
        RECT -54.675 528.190 -53.175 528.420 ;
        RECT -40.905 528.240 -40.405 528.470 ;
        RECT -37.410 528.230 -35.910 528.460 ;
        RECT -58.170 527.220 -57.670 527.450 ;
        RECT -40.905 527.260 -40.405 527.490 ;
        RECT -58.170 526.240 -57.670 526.470 ;
        RECT -54.030 526.265 -53.030 526.495 ;
        RECT -40.905 526.280 -40.405 526.510 ;
        RECT -36.765 526.305 -35.765 526.535 ;
        RECT -59.175 525.155 -57.675 525.385 ;
        RECT -54.030 525.285 -53.030 525.515 ;
        RECT -41.910 525.195 -40.410 525.425 ;
        RECT -36.765 525.325 -35.765 525.555 ;
        RECT -59.175 524.175 -57.675 524.405 ;
        RECT -54.030 524.305 -53.030 524.535 ;
        RECT -41.910 524.215 -40.410 524.445 ;
        RECT -36.765 524.345 -35.765 524.575 ;
        RECT -59.175 523.195 -57.675 523.425 ;
        RECT -54.030 523.325 -53.030 523.555 ;
        RECT -41.910 523.235 -40.410 523.465 ;
        RECT -36.765 523.365 -35.765 523.595 ;
        RECT -57.065 508.300 -56.110 509.055 ;
        RECT -56.940 507.505 -56.245 508.300 ;
        RECT -57.000 507.050 -56.185 507.505 ;
        RECT -54.920 506.750 -54.420 506.980 ;
        RECT -60.470 506.100 -57.470 506.330 ;
        RECT -54.920 505.770 -54.420 506.000 ;
        RECT -54.920 504.790 -54.420 505.020 ;
        RECT -60.470 503.985 -57.470 504.215 ;
        RECT -54.920 503.810 -54.420 504.040 ;
        RECT -60.470 503.005 -57.470 503.235 ;
        RECT -54.915 502.725 -53.415 502.955 ;
        RECT -58.410 501.755 -57.910 501.985 ;
        RECT -54.915 501.745 -53.415 501.975 ;
        RECT -40.840 501.390 -39.340 501.620 ;
        RECT -58.410 500.775 -57.910 501.005 ;
        RECT -54.915 500.765 -53.415 500.995 ;
        RECT -40.840 500.410 -39.340 500.640 ;
        RECT -58.410 499.795 -57.910 500.025 ;
        RECT -41.840 499.270 -39.340 499.500 ;
        RECT -58.410 498.815 -57.910 499.045 ;
        RECT -54.270 498.840 -53.270 499.070 ;
        RECT -41.840 498.620 -39.340 498.850 ;
        RECT -59.415 497.730 -57.915 497.960 ;
        RECT -54.270 497.860 -53.270 498.090 ;
        RECT -59.415 496.750 -57.915 496.980 ;
        RECT -54.270 496.880 -53.270 497.110 ;
        RECT -59.415 495.770 -57.915 496.000 ;
        RECT -54.270 495.900 -53.270 496.130 ;
        RECT -41.840 495.645 -39.340 495.875 ;
        RECT -41.840 494.665 -39.340 494.895 ;
        RECT -56.675 489.950 -55.990 490.430 ;
        RECT -39.645 490.000 -38.895 490.550 ;
        RECT -60.315 487.760 -57.315 487.990 ;
        RECT -60.315 485.645 -57.315 485.875 ;
        RECT -60.315 484.665 -57.315 484.895 ;
        RECT -56.545 484.350 -56.135 489.950 ;
        RECT -39.555 489.230 -39.075 490.000 ;
        RECT -39.585 488.860 -38.995 489.230 ;
        RECT -54.765 488.410 -54.265 488.640 ;
        RECT -37.500 488.450 -37.000 488.680 ;
        RECT -43.050 487.800 -40.050 488.030 ;
        RECT -54.765 487.430 -54.265 487.660 ;
        RECT -37.500 487.470 -37.000 487.700 ;
        RECT -54.765 486.450 -54.265 486.680 ;
        RECT -37.500 486.490 -37.000 486.720 ;
        RECT -54.765 485.470 -54.265 485.700 ;
        RECT -43.050 485.685 -40.050 485.915 ;
        RECT -37.500 485.510 -37.000 485.740 ;
        RECT -43.050 484.705 -40.050 484.935 ;
        RECT -54.760 484.385 -53.260 484.615 ;
        RECT -37.495 484.425 -35.995 484.655 ;
        RECT -58.255 483.415 -57.755 483.645 ;
        RECT -56.580 483.435 -55.930 484.350 ;
        RECT -54.760 483.405 -53.260 483.635 ;
        RECT -40.990 483.455 -40.490 483.685 ;
        RECT -37.495 483.445 -35.995 483.675 ;
        RECT -58.255 482.435 -57.755 482.665 ;
        RECT -54.760 482.425 -53.260 482.655 ;
        RECT -40.990 482.475 -40.490 482.705 ;
        RECT -37.495 482.465 -35.995 482.695 ;
        RECT -58.255 481.455 -57.755 481.685 ;
        RECT -40.990 481.495 -40.490 481.725 ;
        RECT -58.255 480.475 -57.755 480.705 ;
        RECT -54.115 480.500 -53.115 480.730 ;
        RECT -40.990 480.515 -40.490 480.745 ;
        RECT -36.850 480.540 -35.850 480.770 ;
        RECT -59.260 479.390 -57.760 479.620 ;
        RECT -54.115 479.520 -53.115 479.750 ;
        RECT -41.995 479.430 -40.495 479.660 ;
        RECT -36.850 479.560 -35.850 479.790 ;
        RECT -59.260 478.410 -57.760 478.640 ;
        RECT -54.115 478.540 -53.115 478.770 ;
        RECT -41.995 478.450 -40.495 478.680 ;
        RECT -36.850 478.580 -35.850 478.810 ;
        RECT -59.260 477.430 -57.760 477.660 ;
        RECT -54.115 477.560 -53.115 477.790 ;
        RECT -41.995 477.470 -40.495 477.700 ;
        RECT -36.850 477.600 -35.850 477.830 ;
        RECT -57.395 464.530 -56.440 465.285 ;
        RECT -57.270 463.735 -56.575 464.530 ;
        RECT -57.330 463.280 -56.515 463.735 ;
        RECT -55.250 462.980 -54.750 463.210 ;
        RECT -60.800 462.330 -57.800 462.560 ;
        RECT -55.250 462.000 -54.750 462.230 ;
        RECT -55.250 461.020 -54.750 461.250 ;
        RECT -60.800 460.215 -57.800 460.445 ;
        RECT -55.250 460.040 -54.750 460.270 ;
        RECT -60.800 459.235 -57.800 459.465 ;
        RECT -55.245 458.955 -53.745 459.185 ;
        RECT -58.740 457.985 -58.240 458.215 ;
        RECT -55.245 457.975 -53.745 458.205 ;
        RECT -41.170 457.620 -39.670 457.850 ;
        RECT -58.740 457.005 -58.240 457.235 ;
        RECT -55.245 456.995 -53.745 457.225 ;
        RECT -41.170 456.640 -39.670 456.870 ;
        RECT -58.740 456.025 -58.240 456.255 ;
        RECT -42.170 455.500 -39.670 455.730 ;
        RECT -58.740 455.045 -58.240 455.275 ;
        RECT -54.600 455.070 -53.600 455.300 ;
        RECT -42.170 454.850 -39.670 455.080 ;
        RECT -59.745 453.960 -58.245 454.190 ;
        RECT -54.600 454.090 -53.600 454.320 ;
        RECT -59.745 452.980 -58.245 453.210 ;
        RECT -54.600 453.110 -53.600 453.340 ;
        RECT -59.745 452.000 -58.245 452.230 ;
        RECT -54.600 452.130 -53.600 452.360 ;
        RECT -42.170 451.875 -39.670 452.105 ;
        RECT -42.170 450.895 -39.670 451.125 ;
        RECT -57.005 446.180 -56.320 446.660 ;
        RECT -39.975 446.230 -39.225 446.780 ;
        RECT -60.645 443.990 -57.645 444.220 ;
        RECT -60.645 441.875 -57.645 442.105 ;
        RECT -60.645 440.895 -57.645 441.125 ;
        RECT -56.875 440.580 -56.465 446.180 ;
        RECT -39.885 445.460 -39.405 446.230 ;
        RECT -39.915 445.090 -39.325 445.460 ;
        RECT -55.095 444.640 -54.595 444.870 ;
        RECT -37.830 444.680 -37.330 444.910 ;
        RECT -43.380 444.030 -40.380 444.260 ;
        RECT -55.095 443.660 -54.595 443.890 ;
        RECT -37.830 443.700 -37.330 443.930 ;
        RECT -55.095 442.680 -54.595 442.910 ;
        RECT -37.830 442.720 -37.330 442.950 ;
        RECT -55.095 441.700 -54.595 441.930 ;
        RECT -43.380 441.915 -40.380 442.145 ;
        RECT -37.830 441.740 -37.330 441.970 ;
        RECT -43.380 440.935 -40.380 441.165 ;
        RECT -55.090 440.615 -53.590 440.845 ;
        RECT -37.825 440.655 -36.325 440.885 ;
        RECT -58.585 439.645 -58.085 439.875 ;
        RECT -56.910 439.665 -56.260 440.580 ;
        RECT -55.090 439.635 -53.590 439.865 ;
        RECT -41.320 439.685 -40.820 439.915 ;
        RECT -37.825 439.675 -36.325 439.905 ;
        RECT -58.585 438.665 -58.085 438.895 ;
        RECT -55.090 438.655 -53.590 438.885 ;
        RECT -41.320 438.705 -40.820 438.935 ;
        RECT -37.825 438.695 -36.325 438.925 ;
        RECT -58.585 437.685 -58.085 437.915 ;
        RECT -41.320 437.725 -40.820 437.955 ;
        RECT -58.585 436.705 -58.085 436.935 ;
        RECT -54.445 436.730 -53.445 436.960 ;
        RECT -41.320 436.745 -40.820 436.975 ;
        RECT -37.180 436.770 -36.180 437.000 ;
        RECT -59.590 435.620 -58.090 435.850 ;
        RECT -54.445 435.750 -53.445 435.980 ;
        RECT -42.325 435.660 -40.825 435.890 ;
        RECT -37.180 435.790 -36.180 436.020 ;
        RECT -59.590 434.640 -58.090 434.870 ;
        RECT -54.445 434.770 -53.445 435.000 ;
        RECT -42.325 434.680 -40.825 434.910 ;
        RECT -37.180 434.810 -36.180 435.040 ;
        RECT -59.590 433.660 -58.090 433.890 ;
        RECT -54.445 433.790 -53.445 434.020 ;
        RECT -42.325 433.700 -40.825 433.930 ;
        RECT -37.180 433.830 -36.180 434.060 ;
        RECT -57.565 418.540 -56.610 419.295 ;
        RECT -57.440 417.745 -56.745 418.540 ;
        RECT -57.500 417.290 -56.685 417.745 ;
        RECT -55.420 416.990 -54.920 417.220 ;
        RECT -60.970 416.340 -57.970 416.570 ;
        RECT -55.420 416.010 -54.920 416.240 ;
        RECT -55.420 415.030 -54.920 415.260 ;
        RECT -60.970 414.225 -57.970 414.455 ;
        RECT -55.420 414.050 -54.920 414.280 ;
        RECT -60.970 413.245 -57.970 413.475 ;
        RECT -55.415 412.965 -53.915 413.195 ;
        RECT -58.910 411.995 -58.410 412.225 ;
        RECT -55.415 411.985 -53.915 412.215 ;
        RECT -41.340 411.630 -39.840 411.860 ;
        RECT -58.910 411.015 -58.410 411.245 ;
        RECT -55.415 411.005 -53.915 411.235 ;
        RECT -41.340 410.650 -39.840 410.880 ;
        RECT -58.910 410.035 -58.410 410.265 ;
        RECT -42.340 409.510 -39.840 409.740 ;
        RECT -58.910 409.055 -58.410 409.285 ;
        RECT -54.770 409.080 -53.770 409.310 ;
        RECT -42.340 408.860 -39.840 409.090 ;
        RECT -59.915 407.970 -58.415 408.200 ;
        RECT -54.770 408.100 -53.770 408.330 ;
        RECT -59.915 406.990 -58.415 407.220 ;
        RECT -54.770 407.120 -53.770 407.350 ;
        RECT -59.915 406.010 -58.415 406.240 ;
        RECT -54.770 406.140 -53.770 406.370 ;
        RECT -42.340 405.885 -39.840 406.115 ;
        RECT -42.340 404.905 -39.840 405.135 ;
        RECT -57.175 400.190 -56.490 400.670 ;
        RECT -40.145 400.240 -39.395 400.790 ;
        RECT -60.815 398.000 -57.815 398.230 ;
        RECT -60.815 395.885 -57.815 396.115 ;
        RECT -60.815 394.905 -57.815 395.135 ;
        RECT -57.045 394.590 -56.635 400.190 ;
        RECT -40.055 399.470 -39.575 400.240 ;
        RECT -40.085 399.100 -39.495 399.470 ;
        RECT -55.265 398.650 -54.765 398.880 ;
        RECT -38.000 398.690 -37.500 398.920 ;
        RECT -43.550 398.040 -40.550 398.270 ;
        RECT -55.265 397.670 -54.765 397.900 ;
        RECT -38.000 397.710 -37.500 397.940 ;
        RECT -55.265 396.690 -54.765 396.920 ;
        RECT -38.000 396.730 -37.500 396.960 ;
        RECT -55.265 395.710 -54.765 395.940 ;
        RECT -43.550 395.925 -40.550 396.155 ;
        RECT -38.000 395.750 -37.500 395.980 ;
        RECT -43.550 394.945 -40.550 395.175 ;
        RECT -55.260 394.625 -53.760 394.855 ;
        RECT -37.995 394.665 -36.495 394.895 ;
        RECT -58.755 393.655 -58.255 393.885 ;
        RECT -57.080 393.675 -56.430 394.590 ;
        RECT -55.260 393.645 -53.760 393.875 ;
        RECT -41.490 393.695 -40.990 393.925 ;
        RECT -37.995 393.685 -36.495 393.915 ;
        RECT -58.755 392.675 -58.255 392.905 ;
        RECT -55.260 392.665 -53.760 392.895 ;
        RECT -41.490 392.715 -40.990 392.945 ;
        RECT -37.995 392.705 -36.495 392.935 ;
        RECT -58.755 391.695 -58.255 391.925 ;
        RECT -41.490 391.735 -40.990 391.965 ;
        RECT -58.755 390.715 -58.255 390.945 ;
        RECT -54.615 390.740 -53.615 390.970 ;
        RECT -41.490 390.755 -40.990 390.985 ;
        RECT -37.350 390.780 -36.350 391.010 ;
        RECT -59.760 389.630 -58.260 389.860 ;
        RECT -54.615 389.760 -53.615 389.990 ;
        RECT -42.495 389.670 -40.995 389.900 ;
        RECT -37.350 389.800 -36.350 390.030 ;
        RECT -59.760 388.650 -58.260 388.880 ;
        RECT -54.615 388.780 -53.615 389.010 ;
        RECT -42.495 388.690 -40.995 388.920 ;
        RECT -37.350 388.820 -36.350 389.050 ;
        RECT -59.760 387.670 -58.260 387.900 ;
        RECT -54.615 387.800 -53.615 388.030 ;
        RECT -42.495 387.710 -40.995 387.940 ;
        RECT -37.350 387.840 -36.350 388.070 ;
        RECT -57.370 374.225 -56.415 374.980 ;
        RECT -57.245 373.430 -56.550 374.225 ;
        RECT -57.305 372.975 -56.490 373.430 ;
        RECT -55.225 372.675 -54.725 372.905 ;
        RECT -60.775 372.025 -57.775 372.255 ;
        RECT -55.225 371.695 -54.725 371.925 ;
        RECT -55.225 370.715 -54.725 370.945 ;
        RECT -60.775 369.910 -57.775 370.140 ;
        RECT -55.225 369.735 -54.725 369.965 ;
        RECT -60.775 368.930 -57.775 369.160 ;
        RECT -55.220 368.650 -53.720 368.880 ;
        RECT -58.715 367.680 -58.215 367.910 ;
        RECT -55.220 367.670 -53.720 367.900 ;
        RECT -41.145 367.315 -39.645 367.545 ;
        RECT -58.715 366.700 -58.215 366.930 ;
        RECT -55.220 366.690 -53.720 366.920 ;
        RECT -41.145 366.335 -39.645 366.565 ;
        RECT -58.715 365.720 -58.215 365.950 ;
        RECT -42.145 365.195 -39.645 365.425 ;
        RECT -58.715 364.740 -58.215 364.970 ;
        RECT -54.575 364.765 -53.575 364.995 ;
        RECT -42.145 364.545 -39.645 364.775 ;
        RECT -59.720 363.655 -58.220 363.885 ;
        RECT -54.575 363.785 -53.575 364.015 ;
        RECT -59.720 362.675 -58.220 362.905 ;
        RECT -54.575 362.805 -53.575 363.035 ;
        RECT -59.720 361.695 -58.220 361.925 ;
        RECT -54.575 361.825 -53.575 362.055 ;
        RECT -42.145 361.570 -39.645 361.800 ;
        RECT -42.145 360.590 -39.645 360.820 ;
        RECT -56.980 355.875 -56.295 356.355 ;
        RECT -39.950 355.925 -39.200 356.475 ;
        RECT -60.620 353.685 -57.620 353.915 ;
        RECT -60.620 351.570 -57.620 351.800 ;
        RECT -60.620 350.590 -57.620 350.820 ;
        RECT -56.850 350.275 -56.440 355.875 ;
        RECT -39.860 355.155 -39.380 355.925 ;
        RECT -39.890 354.785 -39.300 355.155 ;
        RECT -55.070 354.335 -54.570 354.565 ;
        RECT -37.805 354.375 -37.305 354.605 ;
        RECT -43.355 353.725 -40.355 353.955 ;
        RECT -55.070 353.355 -54.570 353.585 ;
        RECT -37.805 353.395 -37.305 353.625 ;
        RECT -55.070 352.375 -54.570 352.605 ;
        RECT -37.805 352.415 -37.305 352.645 ;
        RECT -55.070 351.395 -54.570 351.625 ;
        RECT -43.355 351.610 -40.355 351.840 ;
        RECT -37.805 351.435 -37.305 351.665 ;
        RECT -43.355 350.630 -40.355 350.860 ;
        RECT -55.065 350.310 -53.565 350.540 ;
        RECT -37.800 350.350 -36.300 350.580 ;
        RECT -58.560 349.340 -58.060 349.570 ;
        RECT -56.885 349.360 -56.235 350.275 ;
        RECT -55.065 349.330 -53.565 349.560 ;
        RECT -41.295 349.380 -40.795 349.610 ;
        RECT -37.800 349.370 -36.300 349.600 ;
        RECT -58.560 348.360 -58.060 348.590 ;
        RECT -55.065 348.350 -53.565 348.580 ;
        RECT -41.295 348.400 -40.795 348.630 ;
        RECT -37.800 348.390 -36.300 348.620 ;
        RECT -58.560 347.380 -58.060 347.610 ;
        RECT -41.295 347.420 -40.795 347.650 ;
        RECT -58.560 346.400 -58.060 346.630 ;
        RECT -54.420 346.425 -53.420 346.655 ;
        RECT -41.295 346.440 -40.795 346.670 ;
        RECT -37.155 346.465 -36.155 346.695 ;
        RECT -59.565 345.315 -58.065 345.545 ;
        RECT -54.420 345.445 -53.420 345.675 ;
        RECT -42.300 345.355 -40.800 345.585 ;
        RECT -37.155 345.485 -36.155 345.715 ;
        RECT -59.565 344.335 -58.065 344.565 ;
        RECT -54.420 344.465 -53.420 344.695 ;
        RECT -42.300 344.375 -40.800 344.605 ;
        RECT -37.155 344.505 -36.155 344.735 ;
        RECT -59.565 343.355 -58.065 343.585 ;
        RECT -54.420 343.485 -53.420 343.715 ;
        RECT -42.300 343.395 -40.800 343.625 ;
        RECT -37.155 343.525 -36.155 343.755 ;
        RECT -57.315 332.025 -56.360 332.780 ;
        RECT -57.190 331.230 -56.495 332.025 ;
        RECT -57.250 330.775 -56.435 331.230 ;
        RECT -55.170 330.475 -54.670 330.705 ;
        RECT -60.720 329.825 -57.720 330.055 ;
        RECT -55.170 329.495 -54.670 329.725 ;
        RECT -55.170 328.515 -54.670 328.745 ;
        RECT -60.720 327.710 -57.720 327.940 ;
        RECT -55.170 327.535 -54.670 327.765 ;
        RECT -60.720 326.730 -57.720 326.960 ;
        RECT -55.165 326.450 -53.665 326.680 ;
        RECT -58.660 325.480 -58.160 325.710 ;
        RECT -55.165 325.470 -53.665 325.700 ;
        RECT -41.090 325.115 -39.590 325.345 ;
        RECT -58.660 324.500 -58.160 324.730 ;
        RECT -55.165 324.490 -53.665 324.720 ;
        RECT -41.090 324.135 -39.590 324.365 ;
        RECT -58.660 323.520 -58.160 323.750 ;
        RECT -42.090 322.995 -39.590 323.225 ;
        RECT -58.660 322.540 -58.160 322.770 ;
        RECT -54.520 322.565 -53.520 322.795 ;
        RECT -42.090 322.345 -39.590 322.575 ;
        RECT -59.665 321.455 -58.165 321.685 ;
        RECT -54.520 321.585 -53.520 321.815 ;
        RECT -59.665 320.475 -58.165 320.705 ;
        RECT -54.520 320.605 -53.520 320.835 ;
        RECT -59.665 319.495 -58.165 319.725 ;
        RECT -54.520 319.625 -53.520 319.855 ;
        RECT -42.090 319.370 -39.590 319.600 ;
        RECT -42.090 318.390 -39.590 318.620 ;
        RECT -56.925 313.675 -56.240 314.155 ;
        RECT -39.895 313.725 -39.145 314.275 ;
        RECT -60.565 311.485 -57.565 311.715 ;
        RECT -60.565 309.370 -57.565 309.600 ;
        RECT -60.565 308.390 -57.565 308.620 ;
        RECT -56.795 308.075 -56.385 313.675 ;
        RECT -39.805 312.955 -39.325 313.725 ;
        RECT -39.835 312.585 -39.245 312.955 ;
        RECT -55.015 312.135 -54.515 312.365 ;
        RECT -37.750 312.175 -37.250 312.405 ;
        RECT -43.300 311.525 -40.300 311.755 ;
        RECT -55.015 311.155 -54.515 311.385 ;
        RECT -37.750 311.195 -37.250 311.425 ;
        RECT -55.015 310.175 -54.515 310.405 ;
        RECT -37.750 310.215 -37.250 310.445 ;
        RECT -55.015 309.195 -54.515 309.425 ;
        RECT -43.300 309.410 -40.300 309.640 ;
        RECT -37.750 309.235 -37.250 309.465 ;
        RECT -43.300 308.430 -40.300 308.660 ;
        RECT -55.010 308.110 -53.510 308.340 ;
        RECT -37.745 308.150 -36.245 308.380 ;
        RECT -58.505 307.140 -58.005 307.370 ;
        RECT -56.830 307.160 -56.180 308.075 ;
        RECT -55.010 307.130 -53.510 307.360 ;
        RECT -41.240 307.180 -40.740 307.410 ;
        RECT -37.745 307.170 -36.245 307.400 ;
        RECT -58.505 306.160 -58.005 306.390 ;
        RECT -55.010 306.150 -53.510 306.380 ;
        RECT -41.240 306.200 -40.740 306.430 ;
        RECT -37.745 306.190 -36.245 306.420 ;
        RECT -58.505 305.180 -58.005 305.410 ;
        RECT -41.240 305.220 -40.740 305.450 ;
        RECT -58.505 304.200 -58.005 304.430 ;
        RECT -54.365 304.225 -53.365 304.455 ;
        RECT -41.240 304.240 -40.740 304.470 ;
        RECT -37.100 304.265 -36.100 304.495 ;
        RECT -59.510 303.115 -58.010 303.345 ;
        RECT -54.365 303.245 -53.365 303.475 ;
        RECT -42.245 303.155 -40.745 303.385 ;
        RECT -37.100 303.285 -36.100 303.515 ;
        RECT -59.510 302.135 -58.010 302.365 ;
        RECT -54.365 302.265 -53.365 302.495 ;
        RECT -42.245 302.175 -40.745 302.405 ;
        RECT -37.100 302.305 -36.100 302.535 ;
        RECT -59.510 301.155 -58.010 301.385 ;
        RECT -54.365 301.285 -53.365 301.515 ;
        RECT -42.245 301.195 -40.745 301.425 ;
        RECT -37.100 301.325 -36.100 301.555 ;
        RECT -56.365 289.390 -52.865 289.620 ;
        RECT -38.865 289.110 -37.865 289.340 ;
        RECT -56.365 288.410 -52.865 288.640 ;
        RECT -45.455 288.620 -44.455 288.850 ;
        RECT -38.865 288.130 -37.865 288.360 ;
        RECT -45.455 287.640 -44.455 287.870 ;
        RECT -56.365 287.390 -52.865 287.620 ;
        RECT -38.865 287.150 -37.865 287.380 ;
        RECT -45.455 286.660 -44.455 286.890 ;
        RECT -56.365 286.410 -52.865 286.640 ;
        RECT -38.865 284.925 -37.865 285.155 ;
        RECT -56.365 284.390 -52.865 284.620 ;
        RECT -38.865 283.945 -37.865 284.175 ;
        RECT -56.365 283.410 -52.865 283.640 ;
        RECT -38.865 282.965 -37.865 283.195 ;
        RECT -56.365 282.390 -52.865 282.620 ;
        RECT -56.365 281.410 -52.865 281.640 ;
        RECT -45.455 279.905 -44.455 280.135 ;
        RECT -56.365 279.390 -52.865 279.620 ;
        RECT -45.455 278.925 -44.455 279.155 ;
        RECT -56.365 278.410 -52.865 278.640 ;
        RECT -45.455 277.945 -44.455 278.175 ;
        RECT -56.365 277.390 -52.865 277.620 ;
        RECT -56.365 276.410 -52.865 276.640 ;
        RECT -38.865 275.610 -37.865 275.840 ;
        RECT -45.455 275.120 -44.455 275.350 ;
        RECT -38.865 274.630 -37.865 274.860 ;
        RECT -50.215 274.220 -48.215 274.450 ;
        RECT -56.720 273.970 -55.720 274.200 ;
        RECT -45.455 274.140 -44.455 274.370 ;
        RECT -38.865 273.650 -37.865 273.880 ;
        RECT -50.215 273.240 -48.215 273.470 ;
        RECT -56.720 272.990 -55.720 273.220 ;
        RECT -45.455 273.160 -44.455 273.390 ;
        RECT -50.215 272.260 -48.215 272.490 ;
        RECT -56.720 272.010 -55.720 272.240 ;
        RECT -38.865 271.425 -37.865 271.655 ;
        RECT -38.865 270.445 -37.865 270.675 ;
        RECT -56.755 269.345 -55.755 269.575 ;
        RECT -38.865 269.465 -37.865 269.695 ;
        RECT -56.755 268.365 -55.755 268.595 ;
        RECT -45.455 266.405 -44.455 266.635 ;
        RECT -56.755 265.655 -55.755 265.885 ;
        RECT -45.455 265.425 -44.455 265.655 ;
        RECT -56.755 264.675 -55.755 264.905 ;
        RECT -45.455 264.445 -44.455 264.675 ;
        RECT -56.755 263.695 -55.755 263.925 ;
        RECT -56.755 262.715 -55.755 262.945 ;
        RECT -45.455 261.995 -44.455 262.225 ;
        RECT -45.455 261.015 -44.455 261.245 ;
        RECT -45.455 260.035 -44.455 260.265 ;
        RECT -56.585 259.115 -54.585 259.345 ;
        RECT -56.585 258.135 -54.585 258.365 ;
        RECT -56.585 254.385 -54.585 254.615 ;
        RECT -44.855 254.410 -41.855 254.640 ;
        RECT -56.585 253.405 -54.585 253.635 ;
        RECT -44.855 253.430 -41.855 253.660 ;
        RECT -68.235 248.470 -67.235 248.700 ;
        RECT -61.645 247.980 -60.645 248.210 ;
        RECT -68.235 247.490 -67.235 247.720 ;
        RECT -61.645 247.000 -60.645 247.230 ;
        RECT -68.235 246.510 -67.235 246.740 ;
        RECT -61.645 246.020 -60.645 246.250 ;
        RECT -68.235 244.285 -67.235 244.515 ;
        RECT -68.235 243.305 -67.235 243.535 ;
        RECT -68.235 242.325 -67.235 242.555 ;
        RECT -61.645 239.265 -60.645 239.495 ;
        RECT -61.645 238.285 -60.645 238.515 ;
        RECT -61.645 237.305 -60.645 237.535 ;
        RECT -68.235 234.970 -67.235 235.200 ;
        RECT -61.645 234.480 -60.645 234.710 ;
        RECT -68.235 233.990 -67.235 234.220 ;
        RECT -61.645 233.500 -60.645 233.730 ;
        RECT -68.235 233.010 -67.235 233.240 ;
        RECT -61.645 232.520 -60.645 232.750 ;
        RECT -68.235 230.785 -67.235 231.015 ;
        RECT -68.235 229.805 -67.235 230.035 ;
        RECT -68.235 228.825 -67.235 229.055 ;
        RECT -61.645 225.765 -60.645 225.995 ;
        RECT -61.645 224.785 -60.645 225.015 ;
        RECT -61.645 223.805 -60.645 224.035 ;
        RECT -61.645 221.355 -60.645 221.585 ;
        RECT -61.645 220.375 -60.645 220.605 ;
        RECT -61.645 219.395 -60.645 219.625 ;
        RECT -69.050 203.245 -68.050 203.475 ;
        RECT -57.795 203.295 -56.795 203.525 ;
        RECT -37.615 203.295 -36.615 203.525 ;
        RECT -26.360 203.245 -25.360 203.475 ;
        RECT -69.050 202.265 -68.050 202.495 ;
        RECT -57.795 202.315 -56.795 202.545 ;
        RECT -37.615 202.315 -36.615 202.545 ;
        RECT -26.360 202.265 -25.360 202.495 ;
        RECT -69.050 201.700 -68.050 201.930 ;
        RECT -57.795 201.750 -56.795 201.980 ;
        RECT -37.615 201.750 -36.615 201.980 ;
        RECT -26.360 201.700 -25.360 201.930 ;
        RECT -18.710 201.180 -12.635 202.855 ;
        RECT -69.050 200.720 -68.050 200.950 ;
        RECT -57.795 200.770 -56.795 201.000 ;
        RECT -37.615 200.770 -36.615 201.000 ;
        RECT -26.360 200.720 -25.360 200.950 ;
        RECT -69.050 200.150 -68.050 200.380 ;
        RECT -57.795 200.200 -56.795 200.430 ;
        RECT -37.615 200.200 -36.615 200.430 ;
        RECT -26.360 200.150 -25.360 200.380 ;
        RECT -69.050 199.170 -68.050 199.400 ;
        RECT -57.795 199.220 -56.795 199.450 ;
        RECT -37.615 199.220 -36.615 199.450 ;
        RECT -26.360 199.170 -25.360 199.400 ;
        RECT -69.050 198.190 -68.050 198.420 ;
        RECT -58.815 198.265 -58.135 198.880 ;
        RECT -58.755 192.800 -58.230 198.265 ;
        RECT -57.795 198.240 -56.795 198.470 ;
        RECT -37.615 198.240 -36.615 198.470 ;
        RECT -36.275 198.265 -35.595 198.880 ;
        RECT -36.180 192.800 -35.655 198.265 ;
        RECT -26.360 198.190 -25.360 198.420 ;
        RECT -18.710 196.780 -11.835 201.180 ;
        RECT -58.820 192.185 -58.140 192.800 ;
        RECT -57.850 192.435 -56.850 192.665 ;
        RECT -37.560 192.435 -36.560 192.665 ;
        RECT -36.270 192.185 -35.590 192.800 ;
        RECT -57.850 191.455 -56.850 191.685 ;
        RECT -37.560 191.455 -36.560 191.685 ;
        RECT -57.850 190.475 -56.850 190.705 ;
        RECT -37.560 190.475 -36.560 190.705 ;
        RECT -57.850 189.495 -56.850 189.725 ;
        RECT -37.560 189.495 -36.560 189.725 ;
        RECT -69.050 188.245 -68.050 188.475 ;
        RECT -26.360 188.245 -25.360 188.475 ;
        RECT -69.050 187.265 -68.050 187.495 ;
        RECT -26.360 187.265 -25.360 187.495 ;
        RECT -69.050 186.700 -68.050 186.930 ;
        RECT -57.850 186.785 -56.850 187.015 ;
        RECT -37.560 186.785 -36.560 187.015 ;
        RECT -26.360 186.700 -25.360 186.930 ;
        RECT -69.050 185.720 -68.050 185.950 ;
        RECT -58.845 185.405 -58.165 186.020 ;
        RECT -57.850 185.805 -56.850 186.035 ;
        RECT -37.560 185.805 -36.560 186.035 ;
        RECT -36.245 185.405 -35.565 186.020 ;
        RECT -26.360 185.720 -25.360 185.950 ;
        RECT -69.050 185.150 -68.050 185.380 ;
        RECT -69.050 184.170 -68.050 184.400 ;
        RECT -58.790 184.015 -58.255 185.405 ;
        RECT -36.155 184.015 -35.620 185.405 ;
        RECT -26.360 185.150 -25.360 185.380 ;
        RECT -26.360 184.170 -25.360 184.400 ;
        RECT -69.050 183.190 -68.050 183.420 ;
        RECT -58.835 183.400 -58.155 184.015 ;
        RECT -57.725 183.670 -56.225 183.900 ;
        RECT -38.185 183.670 -36.685 183.900 ;
        RECT -36.255 183.400 -35.575 184.015 ;
        RECT -26.360 183.190 -25.360 183.420 ;
        RECT -57.725 182.690 -56.225 182.920 ;
        RECT -38.185 182.690 -36.685 182.920 ;
        RECT -57.725 181.710 -56.225 181.940 ;
        RECT -38.185 181.710 -36.685 181.940 ;
        RECT -57.730 180.625 -57.230 180.855 ;
        RECT -37.180 180.625 -36.680 180.855 ;
        RECT -57.730 179.645 -57.230 179.875 ;
        RECT -37.180 179.645 -36.680 179.875 ;
        RECT -57.730 178.665 -57.230 178.895 ;
        RECT -37.180 178.665 -36.680 178.895 ;
        RECT -58.720 177.260 -58.040 177.875 ;
        RECT -57.730 177.685 -57.230 177.915 ;
        RECT -37.180 177.685 -36.680 177.915 ;
        RECT -36.370 177.260 -35.690 177.875 ;
        RECT -69.050 175.745 -68.050 175.975 ;
        RECT -58.640 175.930 -58.105 177.260 ;
        RECT -36.305 175.930 -35.770 177.260 ;
        RECT -58.715 175.315 -58.035 175.930 ;
        RECT -57.735 175.645 -56.235 175.875 ;
        RECT -38.175 175.645 -36.675 175.875 ;
        RECT -36.375 175.315 -35.695 175.930 ;
        RECT -26.360 175.745 -25.360 175.975 ;
        RECT -69.050 174.765 -68.050 174.995 ;
        RECT -57.735 174.665 -56.235 174.895 ;
        RECT -38.175 174.665 -36.675 174.895 ;
        RECT -26.360 174.765 -25.360 174.995 ;
        RECT -69.050 174.200 -68.050 174.430 ;
        RECT -26.360 174.200 -25.360 174.430 ;
        RECT -57.735 173.685 -56.235 173.915 ;
        RECT -38.175 173.685 -36.675 173.915 ;
        RECT -69.050 173.220 -68.050 173.450 ;
        RECT -26.360 173.220 -25.360 173.450 ;
        RECT -69.050 172.650 -68.050 172.880 ;
        RECT -57.740 172.600 -57.240 172.830 ;
        RECT -37.170 172.600 -36.670 172.830 ;
        RECT -26.360 172.650 -25.360 172.880 ;
        RECT -69.050 171.670 -68.050 171.900 ;
        RECT -57.740 171.620 -57.240 171.850 ;
        RECT -37.170 171.620 -36.670 171.850 ;
        RECT -26.360 171.670 -25.360 171.900 ;
        RECT -69.050 170.690 -68.050 170.920 ;
        RECT -57.740 170.640 -57.240 170.870 ;
        RECT -37.170 170.640 -36.670 170.870 ;
        RECT -26.360 170.690 -25.360 170.920 ;
        RECT -57.740 169.660 -57.240 169.890 ;
        RECT -37.170 169.660 -36.670 169.890 ;
        RECT -57.805 167.625 -56.805 167.855 ;
        RECT -37.605 167.625 -36.605 167.855 ;
        RECT -57.805 166.645 -56.805 166.875 ;
        RECT -37.605 166.645 -36.605 166.875 ;
        RECT -65.765 165.670 -65.085 165.695 ;
        RECT -62.995 165.690 -62.685 166.605 ;
        RECT -63.000 165.670 -62.685 165.690 ;
        RECT -65.765 165.100 -62.685 165.670 ;
        RECT -57.805 165.665 -56.805 165.895 ;
        RECT -37.605 165.665 -36.605 165.895 ;
        RECT -31.725 165.690 -31.415 166.605 ;
        RECT -31.725 165.670 -31.410 165.690 ;
        RECT -29.325 165.670 -28.645 165.695 ;
        RECT -65.765 165.080 -65.085 165.100 ;
        RECT -63.000 165.075 -62.685 165.100 ;
        RECT -31.725 165.100 -28.645 165.670 ;
        RECT -31.725 165.075 -31.410 165.100 ;
        RECT -29.325 165.080 -28.645 165.100 ;
        RECT -57.805 164.685 -56.805 164.915 ;
        RECT -37.605 164.685 -36.605 164.915 ;
        RECT -69.050 163.245 -68.050 163.475 ;
        RECT -26.360 163.245 -25.360 163.475 ;
        RECT -69.050 162.265 -68.050 162.495 ;
        RECT -26.360 162.265 -25.360 162.495 ;
        RECT -57.805 161.975 -56.805 162.205 ;
        RECT -37.605 161.975 -36.605 162.205 ;
        RECT -69.050 161.700 -68.050 161.930 ;
        RECT -26.360 161.700 -25.360 161.930 ;
        RECT -69.050 160.720 -68.050 160.950 ;
        RECT -58.780 160.425 -58.100 161.040 ;
        RECT -57.805 160.995 -56.805 161.225 ;
        RECT -37.605 160.995 -36.605 161.225 ;
        RECT -36.310 160.425 -35.630 161.040 ;
        RECT -26.360 160.720 -25.360 160.950 ;
        RECT -69.050 160.150 -68.050 160.380 ;
        RECT -58.715 159.570 -58.140 160.425 ;
        RECT -36.270 159.570 -35.695 160.425 ;
        RECT -26.360 160.150 -25.360 160.380 ;
        RECT -69.050 159.170 -68.050 159.400 ;
        RECT -58.775 158.955 -58.095 159.570 ;
        RECT -57.890 159.285 -56.890 159.515 ;
        RECT -37.520 159.285 -36.520 159.515 ;
        RECT -36.315 158.955 -35.635 159.570 ;
        RECT -26.360 159.170 -25.360 159.400 ;
        RECT -69.050 158.190 -68.050 158.420 ;
        RECT -57.890 158.305 -56.890 158.535 ;
        RECT -37.520 158.305 -36.520 158.535 ;
        RECT -26.360 158.190 -25.360 158.420 ;
        RECT -57.890 157.325 -56.890 157.555 ;
        RECT -37.520 157.325 -36.520 157.555 ;
        RECT -57.890 154.875 -56.890 155.105 ;
        RECT -37.520 154.875 -36.520 155.105 ;
        RECT -57.890 153.895 -56.890 154.125 ;
        RECT -37.520 153.895 -36.520 154.125 ;
        RECT -65.765 153.255 -65.085 153.280 ;
        RECT -62.825 153.255 -62.145 153.275 ;
        RECT -65.765 152.685 -62.145 153.255 ;
        RECT -32.265 153.255 -31.585 153.275 ;
        RECT -29.325 153.255 -28.645 153.280 ;
        RECT -57.890 152.915 -56.890 153.145 ;
        RECT -37.520 152.915 -36.520 153.145 ;
        RECT -65.765 152.665 -65.085 152.685 ;
        RECT -62.825 152.660 -62.145 152.685 ;
        RECT -32.265 152.685 -28.645 153.255 ;
        RECT -32.265 152.660 -31.585 152.685 ;
        RECT -29.325 152.665 -28.645 152.685 ;
        RECT -69.050 150.745 -68.050 150.975 ;
        RECT -26.360 150.745 -25.360 150.975 ;
        RECT -69.050 149.765 -68.050 149.995 ;
        RECT -51.300 149.855 -50.300 150.085 ;
        RECT -44.110 149.855 -43.110 150.085 ;
        RECT -26.360 149.765 -25.360 149.995 ;
        RECT -69.050 149.200 -68.050 149.430 ;
        RECT -26.360 149.200 -25.360 149.430 ;
        RECT -51.300 148.875 -50.300 149.105 ;
        RECT -44.110 148.875 -43.110 149.105 ;
        RECT -69.050 148.220 -68.050 148.450 ;
        RECT -26.360 148.220 -25.360 148.450 ;
        RECT -51.300 147.895 -50.300 148.125 ;
        RECT -44.110 147.895 -43.110 148.125 ;
        RECT -69.050 147.650 -68.050 147.880 ;
        RECT -26.360 147.650 -25.360 147.880 ;
        RECT -69.050 146.670 -68.050 146.900 ;
        RECT -26.360 146.670 -25.360 146.900 ;
        RECT -57.890 146.160 -56.890 146.390 ;
        RECT -37.520 146.160 -36.520 146.390 ;
        RECT -69.050 145.690 -68.050 145.920 ;
        RECT -51.300 145.670 -50.300 145.900 ;
        RECT -44.110 145.670 -43.110 145.900 ;
        RECT -26.360 145.690 -25.360 145.920 ;
        RECT -57.890 145.180 -56.890 145.410 ;
        RECT -37.520 145.180 -36.520 145.410 ;
        RECT -51.300 144.690 -50.300 144.920 ;
        RECT -44.110 144.690 -43.110 144.920 ;
        RECT -57.890 144.200 -56.890 144.430 ;
        RECT -37.520 144.200 -36.520 144.430 ;
        RECT -51.300 143.710 -50.300 143.940 ;
        RECT -44.110 143.710 -43.110 143.940 ;
        RECT -57.890 141.375 -56.890 141.605 ;
        RECT -37.520 141.375 -36.520 141.605 ;
        RECT -65.940 140.420 -65.260 140.445 ;
        RECT -62.105 140.420 -61.425 140.440 ;
        RECT -65.940 139.850 -61.425 140.420 ;
        RECT -57.890 140.395 -56.890 140.625 ;
        RECT -37.520 140.395 -36.520 140.625 ;
        RECT -32.985 140.420 -32.305 140.440 ;
        RECT -29.150 140.420 -28.470 140.445 ;
        RECT -65.940 139.830 -65.260 139.850 ;
        RECT -62.105 139.825 -61.425 139.850 ;
        RECT -32.985 139.850 -28.470 140.420 ;
        RECT -32.985 139.825 -32.305 139.850 ;
        RECT -29.150 139.830 -28.470 139.850 ;
        RECT -57.890 139.415 -56.890 139.645 ;
        RECT -37.520 139.415 -36.520 139.645 ;
        RECT -69.050 138.245 -68.050 138.475 ;
        RECT -26.360 138.245 -25.360 138.475 ;
        RECT -69.050 137.265 -68.050 137.495 ;
        RECT -26.360 137.265 -25.360 137.495 ;
        RECT -69.050 136.700 -68.050 136.930 ;
        RECT -26.360 136.700 -25.360 136.930 ;
        RECT -51.300 136.355 -50.300 136.585 ;
        RECT -44.110 136.355 -43.110 136.585 ;
        RECT -69.050 135.720 -68.050 135.950 ;
        RECT -26.360 135.720 -25.360 135.950 ;
        RECT -69.050 135.150 -68.050 135.380 ;
        RECT -51.300 135.375 -50.300 135.605 ;
        RECT -44.110 135.375 -43.110 135.605 ;
        RECT -26.360 135.150 -25.360 135.380 ;
        RECT -69.050 134.170 -68.050 134.400 ;
        RECT -51.300 134.395 -50.300 134.625 ;
        RECT -44.110 134.395 -43.110 134.625 ;
        RECT -26.360 134.170 -25.360 134.400 ;
        RECT -33.005 133.455 -32.005 133.685 ;
        RECT -69.050 133.190 -68.050 133.420 ;
        RECT -26.360 133.190 -25.360 133.420 ;
        RECT -57.890 132.660 -56.890 132.890 ;
        RECT -37.520 132.660 -36.520 132.890 ;
        RECT -33.005 132.475 -32.005 132.705 ;
        RECT -51.300 132.170 -50.300 132.400 ;
        RECT -44.110 132.170 -43.110 132.400 ;
        RECT -57.890 131.680 -56.890 131.910 ;
        RECT -37.520 131.680 -36.520 131.910 ;
        RECT -33.005 131.495 -32.005 131.725 ;
        RECT -51.300 131.190 -50.300 131.420 ;
        RECT -44.110 131.190 -43.110 131.420 ;
        RECT -57.890 130.700 -56.890 130.930 ;
        RECT -37.520 130.700 -36.520 130.930 ;
        RECT -51.300 130.210 -50.300 130.440 ;
        RECT -44.110 130.210 -43.110 130.440 ;
        RECT -52.050 125.880 -49.050 126.110 ;
        RECT -27.380 125.745 -24.380 125.975 ;
        RECT -52.050 124.900 -49.050 125.130 ;
        RECT -27.380 124.765 -24.380 124.995 ;
        RECT -52.050 122.785 -49.050 123.015 ;
        RECT -27.380 122.650 -24.380 122.880 ;
        RECT -56.555 119.915 -55.555 120.145 ;
        RECT -31.920 119.915 -30.920 120.145 ;
        RECT -56.555 118.935 -55.555 119.165 ;
        RECT -31.920 118.935 -30.920 119.165 ;
        RECT -56.555 117.955 -55.555 118.185 ;
        RECT -31.920 117.955 -30.920 118.185 ;
        RECT -56.555 115.505 -55.555 115.735 ;
        RECT -31.920 115.505 -30.920 115.735 ;
        RECT -56.555 114.525 -55.555 114.755 ;
        RECT -31.920 114.525 -30.920 114.755 ;
        RECT -56.555 113.545 -55.555 113.775 ;
        RECT -31.920 113.545 -30.920 113.775 ;
        RECT -49.965 110.485 -48.965 110.715 ;
        RECT -25.330 110.485 -24.330 110.715 ;
        RECT -49.965 109.505 -48.965 109.735 ;
        RECT -25.330 109.505 -24.330 109.735 ;
        RECT -49.965 108.525 -48.965 108.755 ;
        RECT -25.330 108.525 -24.330 108.755 ;
        RECT -56.555 106.790 -55.555 107.020 ;
        RECT -43.560 106.945 -43.060 107.175 ;
        RECT -31.920 106.790 -30.920 107.020 ;
        RECT -49.965 106.300 -48.965 106.530 ;
        RECT -40.510 106.295 -37.510 106.525 ;
        RECT -25.330 106.300 -24.330 106.530 ;
        RECT -56.555 105.810 -55.555 106.040 ;
        RECT -43.560 105.965 -43.060 106.195 ;
        RECT -31.920 105.810 -30.920 106.040 ;
        RECT -49.965 105.320 -48.965 105.550 ;
        RECT -25.330 105.320 -24.330 105.550 ;
        RECT -56.555 104.830 -55.555 105.060 ;
        RECT -43.560 104.985 -43.060 105.215 ;
        RECT -31.920 104.830 -30.920 105.060 ;
        RECT -49.965 104.340 -48.965 104.570 ;
        RECT -43.560 104.005 -43.060 104.235 ;
        RECT -40.510 104.180 -37.510 104.410 ;
        RECT -25.330 104.340 -24.330 104.570 ;
        RECT -40.510 103.200 -37.510 103.430 ;
        RECT -44.565 102.920 -43.065 103.150 ;
        RECT -56.555 102.005 -55.555 102.235 ;
        RECT -44.565 101.940 -43.065 102.170 ;
        RECT -40.070 101.950 -39.570 102.180 ;
        RECT -31.920 102.005 -30.920 102.235 ;
        RECT -56.555 101.025 -55.555 101.255 ;
        RECT -44.565 100.960 -43.065 101.190 ;
        RECT -40.070 100.970 -39.570 101.200 ;
        RECT -31.920 101.025 -30.920 101.255 ;
        RECT -56.555 100.045 -55.555 100.275 ;
        RECT -40.070 99.990 -39.570 100.220 ;
        RECT -31.920 100.045 -30.920 100.275 ;
        RECT -44.710 99.035 -43.710 99.265 ;
        RECT -40.070 99.010 -39.570 99.240 ;
        RECT -44.710 98.055 -43.710 98.285 ;
        RECT -40.065 97.925 -38.565 98.155 ;
        RECT -49.965 96.985 -48.965 97.215 ;
        RECT -44.710 97.075 -43.710 97.305 ;
        RECT -40.065 96.945 -38.565 97.175 ;
        RECT -25.330 96.985 -24.330 97.215 ;
        RECT -49.965 96.005 -48.965 96.235 ;
        RECT -44.710 96.095 -43.710 96.325 ;
        RECT -40.065 95.965 -38.565 96.195 ;
        RECT -25.330 96.005 -24.330 96.235 ;
        RECT -49.965 95.025 -48.965 95.255 ;
        RECT -25.330 95.025 -24.330 95.255 ;
        RECT -56.555 93.290 -55.555 93.520 ;
        RECT -31.920 93.290 -30.920 93.520 ;
        RECT -49.965 92.800 -48.965 93.030 ;
        RECT -25.330 92.800 -24.330 93.030 ;
        RECT -56.555 92.310 -55.555 92.540 ;
        RECT -31.920 92.310 -30.920 92.540 ;
        RECT -49.965 91.820 -48.965 92.050 ;
        RECT -25.330 91.820 -24.330 92.050 ;
        RECT -56.555 91.330 -55.555 91.560 ;
        RECT -31.920 91.330 -30.920 91.560 ;
        RECT -49.965 90.840 -48.965 91.070 ;
        RECT -25.330 90.840 -24.330 91.070 ;
        RECT -63.680 82.000 -63.180 82.230 ;
        RECT -38.680 82.000 -38.180 82.230 ;
        RECT -60.630 81.350 -57.630 81.580 ;
        RECT -35.630 81.350 -32.630 81.580 ;
        RECT -63.680 81.020 -63.180 81.250 ;
        RECT -38.680 81.020 -38.180 81.250 ;
        RECT -63.680 80.040 -63.180 80.270 ;
        RECT -38.680 80.040 -38.180 80.270 ;
        RECT -63.680 79.060 -63.180 79.290 ;
        RECT -60.630 79.235 -57.630 79.465 ;
        RECT -38.680 79.060 -38.180 79.290 ;
        RECT -35.630 79.235 -32.630 79.465 ;
        RECT -60.630 78.255 -57.630 78.485 ;
        RECT -35.630 78.255 -32.630 78.485 ;
        RECT -64.685 77.975 -63.185 78.205 ;
        RECT -39.685 77.975 -38.185 78.205 ;
        RECT -64.685 76.995 -63.185 77.225 ;
        RECT -60.190 77.005 -59.690 77.235 ;
        RECT -39.685 76.995 -38.185 77.225 ;
        RECT -35.190 77.005 -34.690 77.235 ;
        RECT -64.685 76.015 -63.185 76.245 ;
        RECT -60.190 76.025 -59.690 76.255 ;
        RECT -39.685 76.015 -38.185 76.245 ;
        RECT -35.190 76.025 -34.690 76.255 ;
        RECT -60.190 75.045 -59.690 75.275 ;
        RECT -35.190 75.045 -34.690 75.275 ;
        RECT -64.830 74.090 -63.830 74.320 ;
        RECT -60.190 74.065 -59.690 74.295 ;
        RECT -39.830 74.090 -38.830 74.320 ;
        RECT -35.190 74.065 -34.690 74.295 ;
        RECT -64.830 73.110 -63.830 73.340 ;
        RECT -60.185 72.980 -58.685 73.210 ;
        RECT -39.830 73.110 -38.830 73.340 ;
        RECT -35.185 72.980 -33.685 73.210 ;
        RECT -64.830 72.130 -63.830 72.360 ;
        RECT -60.185 72.000 -58.685 72.230 ;
        RECT -39.830 72.130 -38.830 72.360 ;
        RECT -35.185 72.000 -33.685 72.230 ;
        RECT -64.830 71.150 -63.830 71.380 ;
        RECT -60.185 71.020 -58.685 71.250 ;
        RECT -39.830 71.150 -38.830 71.380 ;
        RECT -35.185 71.020 -33.685 71.250 ;
        RECT -62.170 69.480 -61.310 69.805 ;
        RECT -52.490 69.480 -51.655 69.610 ;
        RECT -62.170 68.850 -51.655 69.480 ;
        RECT -62.170 68.845 -61.310 68.850 ;
        RECT -52.490 68.715 -51.655 68.850 ;
        RECT -38.945 68.625 -37.945 68.855 ;
        RECT -29.370 68.825 -28.870 69.055 ;
        RECT -38.945 67.645 -37.945 67.875 ;
        RECT -29.370 67.845 -28.870 68.075 ;
        RECT -29.370 66.865 -28.870 67.095 ;
        RECT -29.370 65.885 -28.870 66.115 ;
        RECT -70.300 64.820 -67.145 65.700 ;
        RECT -56.040 64.990 -54.040 65.220 ;
        RECT -38.945 64.935 -37.945 65.165 ;
        RECT -30.375 64.800 -28.875 65.030 ;
        RECT -56.040 64.010 -54.040 64.240 ;
        RECT -38.945 63.955 -37.945 64.185 ;
        RECT -30.375 63.820 -28.875 64.050 ;
        RECT -38.945 62.975 -37.945 63.205 ;
        RECT -30.375 62.840 -28.875 63.070 ;
        RECT -38.945 61.995 -37.945 62.225 ;
        RECT -56.035 60.465 -54.035 60.695 ;
        RECT -56.035 59.485 -54.035 59.715 ;
        RECT -29.265 59.475 -28.265 59.705 ;
        RECT -38.915 59.115 -38.415 59.345 ;
        RECT -69.480 58.400 -68.480 58.630 ;
        RECT -29.265 58.495 -28.265 58.725 ;
        RECT -38.915 58.135 -38.415 58.365 ;
        RECT -69.480 57.420 -68.480 57.650 ;
        RECT -38.915 57.155 -38.415 57.385 ;
        RECT -69.480 56.440 -68.480 56.670 ;
        RECT -38.915 56.175 -38.415 56.405 ;
        RECT -29.265 55.785 -28.265 56.015 ;
        RECT -69.480 55.460 -68.480 55.690 ;
        RECT -39.920 55.090 -38.420 55.320 ;
        RECT -29.265 54.805 -28.265 55.035 ;
        RECT -57.390 54.435 -54.390 54.665 ;
        RECT -39.920 54.110 -38.420 54.340 ;
        RECT -29.265 53.825 -28.265 54.055 ;
        RECT -57.390 53.455 -54.390 53.685 ;
        RECT -39.920 53.130 -38.420 53.360 ;
        RECT -69.480 52.750 -68.480 52.980 ;
        RECT -29.265 52.845 -28.265 53.075 ;
        RECT -69.480 51.770 -68.480 52.000 ;
        RECT -64.875 17.830 -57.020 34.715 ;
        RECT -17.910 27.770 -11.835 196.780 ;
        RECT 77.940 50.635 78.940 50.865 ;
        RECT 73.925 49.345 74.925 49.575 ;
        RECT 77.940 48.055 78.940 48.285 ;
        RECT 73.925 46.765 74.925 46.995 ;
        RECT 77.940 45.475 78.940 45.705 ;
        RECT 78.630 44.830 79.430 45.060 ;
        RECT 16.875 37.825 20.515 41.000 ;
        RECT -65.610 16.645 -44.765 17.830 ;
        RECT -65.055 11.805 -63.315 16.645 ;
        RECT -59.545 11.805 -57.805 16.645 ;
        RECT -55.075 11.805 -53.335 16.645 ;
        RECT -51.195 11.805 -49.455 16.645 ;
        RECT -48.165 11.805 -46.425 16.645 ;
        RECT -66.975 10.620 -46.130 11.805 ;
        RECT -66.485 7.875 -66.255 9.875 ;
        RECT -65.305 7.875 -65.075 9.875 ;
        RECT -64.125 7.875 -63.895 9.875 ;
        RECT -62.945 7.875 -62.715 9.875 ;
        RECT -61.765 7.875 -61.535 9.875 ;
        RECT -60.585 7.875 -60.355 9.875 ;
        RECT -59.405 7.875 -59.175 9.875 ;
        RECT -58.225 7.875 -57.995 9.875 ;
        RECT -57.045 7.875 -56.815 9.875 ;
        RECT -55.865 7.875 -55.635 9.875 ;
        RECT -54.685 7.875 -54.455 9.875 ;
        RECT -53.505 7.875 -53.275 9.875 ;
        RECT -52.325 7.875 -52.095 9.875 ;
        RECT -51.145 7.875 -50.915 9.875 ;
        RECT -49.965 7.875 -49.735 9.875 ;
        RECT -48.785 7.875 -48.555 9.875 ;
        RECT -47.545 7.875 -47.315 9.875 ;
        RECT -46.365 7.875 -46.135 9.875 ;
        RECT -45.185 7.875 -44.955 9.875 ;
        RECT -44.005 7.875 -43.775 9.875 ;
        RECT -42.825 7.875 -42.595 9.875 ;
        RECT -41.645 7.875 -41.415 9.875 ;
        RECT -40.465 7.875 -40.235 9.875 ;
        RECT -39.285 7.875 -39.055 9.875 ;
        RECT -38.105 7.875 -37.875 9.875 ;
        RECT -37.455 7.875 -37.225 9.875 ;
        RECT -36.275 7.875 -36.045 9.875 ;
        RECT -35.095 7.875 -34.865 9.875 ;
        RECT -33.915 7.875 -33.685 9.875 ;
        RECT -32.735 7.875 -32.505 9.875 ;
        RECT -32.085 7.875 -31.855 9.875 ;
        RECT -30.905 7.875 -30.675 9.875 ;
        RECT -29.725 7.875 -29.495 9.875 ;
        RECT -17.950 9.185 -17.720 10.185 ;
        RECT -16.970 9.185 -16.740 10.185 ;
        RECT -15.990 9.185 -15.760 10.185 ;
        RECT -13.700 9.185 -13.470 10.185 ;
        RECT -12.720 9.185 -12.490 10.185 ;
        RECT -11.740 9.185 -11.510 10.185 ;
        RECT 3.535 8.265 3.765 9.105 ;
        RECT 5.215 8.495 5.445 9.095 ;
        RECT 6.095 8.495 6.325 9.095 ;
        RECT 6.975 8.495 7.205 9.095 ;
        RECT 8.420 8.195 8.650 9.095 ;
        RECT 9.150 8.195 9.380 9.095 ;
        RECT 12.470 8.265 12.700 9.105 ;
        RECT 14.015 8.265 14.245 9.105 ;
        RECT 17.500 6.395 19.375 37.825 ;
        RECT 40.690 33.480 40.920 37.480 ;
        RECT 49.270 33.480 49.500 37.480 ;
        RECT 57.850 33.480 58.080 37.480 ;
        RECT 58.500 33.480 58.730 37.480 ;
        RECT 63.080 33.480 63.310 37.480 ;
        RECT 208.360 20.925 223.200 24.220 ;
        RECT 79.070 18.610 81.655 20.855 ;
        RECT 22.545 10.065 22.775 11.065 ;
        RECT 23.525 10.065 23.755 11.065 ;
        RECT 24.505 10.065 24.735 11.065 ;
        RECT 26.795 10.065 27.025 11.065 ;
        RECT 27.775 10.065 28.005 11.065 ;
        RECT 28.755 10.065 28.985 11.065 ;
        RECT 38.060 9.285 38.290 11.285 ;
        RECT 39.240 9.285 39.470 11.285 ;
        RECT 40.420 9.285 40.650 11.285 ;
        RECT 41.070 9.285 41.300 11.285 ;
        RECT 42.250 9.285 42.480 11.285 ;
        RECT 43.430 9.285 43.660 11.285 ;
        RECT 44.610 9.285 44.840 11.285 ;
        RECT 45.790 9.285 46.020 11.285 ;
        RECT 46.440 9.285 46.670 11.285 ;
        RECT 47.620 9.285 47.850 11.285 ;
        RECT 48.800 9.285 49.030 11.285 ;
        RECT 49.980 9.285 50.210 11.285 ;
        RECT 51.160 9.285 51.390 11.285 ;
        RECT 52.340 9.285 52.570 11.285 ;
        RECT 53.520 9.285 53.750 11.285 ;
        RECT 54.700 9.285 54.930 11.285 ;
        RECT 55.880 9.285 56.110 11.285 ;
        RECT 57.120 9.285 57.350 11.285 ;
        RECT 58.300 9.285 58.530 11.285 ;
        RECT 59.480 9.285 59.710 11.285 ;
        RECT 60.660 9.285 60.890 11.285 ;
        RECT 61.840 9.285 62.070 11.285 ;
        RECT 63.020 9.285 63.250 11.285 ;
        RECT 64.200 9.285 64.430 11.285 ;
        RECT 65.380 9.285 65.610 11.285 ;
        RECT 66.560 9.285 66.790 11.285 ;
        RECT 67.740 9.285 67.970 11.285 ;
        RECT 68.920 9.285 69.150 11.285 ;
        RECT 70.100 9.285 70.330 11.285 ;
        RECT 71.280 9.285 71.510 11.285 ;
        RECT 72.460 9.285 72.690 11.285 ;
        RECT 73.640 9.285 73.870 11.285 ;
        RECT 74.820 9.285 75.050 11.285 ;
        RECT 3.535 5.205 3.765 6.045 ;
        RECT 5.215 5.215 5.445 5.815 ;
        RECT 6.095 5.215 6.325 5.815 ;
        RECT 6.975 5.215 7.205 5.815 ;
        RECT 8.420 5.215 8.650 6.115 ;
        RECT 9.150 5.215 9.380 6.115 ;
        RECT 12.470 5.205 12.700 6.045 ;
        RECT 14.015 5.205 14.245 6.045 ;
        RECT -13.700 3.810 -13.470 4.810 ;
        RECT -12.720 3.810 -12.490 4.810 ;
        RECT -11.740 3.810 -11.510 4.810 ;
        RECT 26.795 4.690 27.025 5.690 ;
        RECT 27.775 4.690 28.005 5.690 ;
        RECT 28.755 4.690 28.985 5.690 ;
        RECT 28.650 3.430 31.040 3.875 ;
        RECT 29.715 1.115 30.675 3.430 ;
        RECT 29.455 -0.610 31.180 1.115 ;
        RECT 79.070 -1.275 81.645 18.610 ;
        RECT 98.940 15.890 99.170 16.890 ;
        RECT 99.920 15.890 100.150 16.890 ;
        RECT 100.900 15.890 101.130 16.890 ;
        RECT 103.190 15.890 103.420 16.890 ;
        RECT 104.170 15.890 104.400 16.890 ;
        RECT 105.150 15.890 105.380 16.890 ;
        RECT 209.325 16.165 210.975 20.925 ;
        RECT 212.770 16.165 214.420 20.925 ;
        RECT 216.215 16.165 217.865 20.925 ;
        RECT 218.760 16.165 220.410 20.925 ;
        RECT 209.135 15.645 220.980 16.165 ;
        RECT 133.440 13.265 134.815 14.380 ;
        RECT 195.900 13.675 196.130 14.675 ;
        RECT 196.880 13.675 197.110 14.675 ;
        RECT 197.860 13.675 198.090 14.675 ;
        RECT 200.310 13.675 200.540 14.675 ;
        RECT 201.290 13.675 201.520 14.675 ;
        RECT 202.270 13.675 202.500 14.675 ;
        RECT 209.025 13.675 209.255 14.675 ;
        RECT 210.005 13.675 210.235 14.675 ;
        RECT 210.985 13.675 211.215 14.675 ;
        RECT 213.810 13.675 214.040 14.675 ;
        RECT 214.790 13.675 215.020 14.675 ;
        RECT 215.770 13.675 216.000 14.675 ;
        RECT 222.525 13.675 222.755 14.675 ;
        RECT 223.505 13.675 223.735 14.675 ;
        RECT 224.485 13.675 224.715 14.675 ;
        RECT 103.190 10.515 103.420 11.515 ;
        RECT 104.170 10.515 104.400 11.515 ;
        RECT 105.150 10.515 105.380 11.515 ;
        RECT 133.810 3.230 134.450 13.265 ;
        RECT 254.450 13.170 254.680 15.170 ;
        RECT 255.630 13.170 255.860 15.170 ;
        RECT 256.810 13.170 257.040 15.170 ;
        RECT 257.460 13.170 257.690 15.170 ;
        RECT 258.640 13.170 258.870 15.170 ;
        RECT 259.820 13.170 260.050 15.170 ;
        RECT 261.000 13.170 261.230 15.170 ;
        RECT 262.180 13.170 262.410 15.170 ;
        RECT 262.830 13.170 263.060 15.170 ;
        RECT 264.010 13.170 264.240 15.170 ;
        RECT 265.190 13.170 265.420 15.170 ;
        RECT 266.370 13.170 266.600 15.170 ;
        RECT 267.550 13.170 267.780 15.170 ;
        RECT 268.730 13.170 268.960 15.170 ;
        RECT 269.910 13.170 270.140 15.170 ;
        RECT 271.090 13.170 271.320 15.170 ;
        RECT 272.270 13.170 272.500 15.170 ;
        RECT 273.510 13.170 273.740 15.170 ;
        RECT 274.690 13.170 274.920 15.170 ;
        RECT 275.870 13.170 276.100 15.170 ;
        RECT 277.050 13.170 277.280 15.170 ;
        RECT 278.230 13.170 278.460 15.170 ;
        RECT 279.410 13.170 279.640 15.170 ;
        RECT 280.590 13.170 280.820 15.170 ;
        RECT 281.770 13.170 282.000 15.170 ;
        RECT 282.950 13.170 283.180 15.170 ;
        RECT 284.130 13.170 284.360 15.170 ;
        RECT 285.310 13.170 285.540 15.170 ;
        RECT 286.490 13.170 286.720 15.170 ;
        RECT 287.670 13.170 287.900 15.170 ;
        RECT 288.850 13.170 289.080 15.170 ;
        RECT 290.030 13.170 290.260 15.170 ;
        RECT 291.210 13.170 291.440 15.170 ;
        RECT 138.575 8.955 138.805 9.955 ;
        RECT 139.365 8.955 139.595 9.955 ;
        RECT 138.575 7.340 138.805 8.340 ;
        RECT 139.365 7.340 139.595 8.340 ;
        RECT 141.305 7.340 141.535 10.285 ;
        RECT 142.885 7.340 143.115 10.285 ;
        RECT 145.115 7.340 145.345 10.310 ;
        RECT 146.535 9.000 146.765 10.310 ;
        RECT 147.325 9.000 147.555 10.310 ;
        RECT 146.430 8.815 147.730 9.000 ;
        RECT 146.430 8.770 150.645 8.815 ;
        RECT 146.555 7.335 146.785 8.770 ;
        RECT 147.345 8.585 150.645 8.770 ;
        RECT 147.345 7.335 147.575 8.585 ;
        RECT 150.415 7.055 150.645 8.585 ;
        RECT 151.620 7.055 151.850 9.200 ;
        RECT 153.200 7.200 153.430 9.200 ;
        RECT 154.780 7.200 155.010 9.200 ;
        RECT 156.360 7.200 156.590 9.200 ;
        RECT 150.415 6.825 151.850 7.055 ;
        RECT 157.940 7.085 158.170 9.200 ;
        RECT 162.850 8.920 163.080 9.920 ;
        RECT 163.640 8.920 163.870 9.920 ;
        RECT 162.850 7.085 163.080 8.305 ;
        RECT 163.640 7.305 163.870 8.305 ;
        RECT 165.580 7.305 165.810 10.250 ;
        RECT 167.160 7.305 167.390 10.250 ;
        RECT 169.390 7.305 169.620 10.275 ;
        RECT 170.810 8.965 171.040 10.275 ;
        RECT 171.600 8.965 171.830 10.275 ;
        RECT 172.750 8.965 172.980 9.205 ;
        RECT 170.705 8.735 172.980 8.965 ;
        RECT 170.830 7.300 171.060 8.735 ;
        RECT 171.620 7.300 171.850 8.735 ;
        RECT 157.940 6.855 163.080 7.085 ;
        RECT 172.750 4.850 172.980 8.735 ;
        RECT 175.295 7.310 175.525 9.310 ;
        RECT 176.875 7.310 177.105 9.310 ;
        RECT 178.455 7.310 178.685 9.310 ;
        RECT 180.035 7.310 180.265 9.310 ;
        RECT 181.615 7.310 181.845 9.310 ;
        RECT 183.900 7.095 184.130 9.095 ;
        RECT 185.480 7.095 185.710 9.095 ;
        RECT 187.060 7.095 187.290 9.095 ;
        RECT 188.640 7.095 188.870 9.095 ;
        RECT 190.220 7.095 190.450 9.095 ;
        RECT 205.330 7.085 205.560 8.085 ;
        RECT 206.310 7.085 206.540 8.085 ;
        RECT 207.290 7.085 207.520 8.085 ;
        RECT 209.515 7.085 209.745 8.085 ;
        RECT 210.495 7.085 210.725 8.085 ;
        RECT 211.475 7.085 211.705 8.085 ;
        RECT 218.830 7.085 219.060 8.085 ;
        RECT 219.810 7.085 220.040 8.085 ;
        RECT 220.790 7.085 221.020 8.085 ;
        RECT 223.015 7.085 223.245 8.085 ;
        RECT 223.995 7.085 224.225 8.085 ;
        RECT 224.975 7.085 225.205 8.085 ;
        RECT 227.865 7.535 228.095 8.535 ;
        RECT 228.845 7.535 229.075 8.535 ;
        RECT 229.825 7.535 230.055 8.535 ;
        RECT 172.750 4.620 175.525 4.850 ;
        RECT 133.810 2.590 135.900 3.230 ;
        RECT 99.800 -0.860 100.030 0.140 ;
        RECT 100.780 -0.860 101.010 0.140 ;
        RECT 101.760 -0.860 101.990 0.140 ;
        RECT 104.050 -0.860 104.280 0.140 ;
        RECT 105.030 -0.860 105.260 0.140 ;
        RECT 106.010 -0.860 106.240 0.140 ;
        RECT 135.260 -0.190 135.900 2.590 ;
        RECT 151.620 2.200 151.850 4.200 ;
        RECT 153.200 2.200 153.430 4.200 ;
        RECT 154.780 2.200 155.010 4.200 ;
        RECT 156.360 2.200 156.590 4.200 ;
        RECT 157.940 2.200 158.170 4.200 ;
        RECT 175.295 2.315 175.525 4.620 ;
        RECT 176.875 2.315 177.105 4.315 ;
        RECT 178.455 2.315 178.685 4.315 ;
        RECT 180.035 2.315 180.265 4.315 ;
        RECT 181.615 2.315 181.845 4.315 ;
        RECT 183.900 2.530 184.130 4.530 ;
        RECT 185.480 2.530 185.710 4.530 ;
        RECT 187.060 2.530 187.290 4.530 ;
        RECT 188.640 2.530 188.870 4.530 ;
        RECT 190.220 2.530 190.450 4.530 ;
        RECT 134.940 -0.345 136.520 -0.190 ;
        RECT 134.940 -0.745 138.835 -0.345 ;
        RECT 134.940 -0.830 136.520 -0.745 ;
        RECT 136.950 -1.530 137.350 -0.745 ;
        RECT 159.330 -0.760 163.115 -0.360 ;
        RECT 159.330 -1.530 159.730 -0.760 ;
        RECT 253.435 -1.385 253.665 0.615 ;
        RECT 254.615 -1.385 254.845 0.615 ;
        RECT 255.795 -1.385 256.025 0.615 ;
        RECT 256.445 -1.385 256.675 0.615 ;
        RECT 257.625 -1.385 257.855 0.615 ;
        RECT 258.805 -1.385 259.035 0.615 ;
        RECT 259.985 -1.385 260.215 0.615 ;
        RECT 261.165 -1.385 261.395 0.615 ;
        RECT 261.815 -1.385 262.045 0.615 ;
        RECT 262.995 -1.385 263.225 0.615 ;
        RECT 264.175 -1.385 264.405 0.615 ;
        RECT 265.355 -1.385 265.585 0.615 ;
        RECT 266.535 -1.385 266.765 0.615 ;
        RECT 267.715 -1.385 267.945 0.615 ;
        RECT 268.895 -1.385 269.125 0.615 ;
        RECT 270.075 -1.385 270.305 0.615 ;
        RECT 271.255 -1.385 271.485 0.615 ;
        RECT 272.495 -1.385 272.725 0.615 ;
        RECT 273.675 -1.385 273.905 0.615 ;
        RECT 274.855 -1.385 275.085 0.615 ;
        RECT 276.035 -1.385 276.265 0.615 ;
        RECT 277.215 -1.385 277.445 0.615 ;
        RECT 278.395 -1.385 278.625 0.615 ;
        RECT 279.575 -1.385 279.805 0.615 ;
        RECT 280.755 -1.385 280.985 0.615 ;
        RECT 281.935 -1.385 282.165 0.615 ;
        RECT 283.115 -1.385 283.345 0.615 ;
        RECT 284.295 -1.385 284.525 0.615 ;
        RECT 285.475 -1.385 285.705 0.615 ;
        RECT 286.655 -1.385 286.885 0.615 ;
        RECT 287.835 -1.385 288.065 0.615 ;
        RECT 289.015 -1.385 289.245 0.615 ;
        RECT 290.195 -1.385 290.425 0.615 ;
        RECT -25.290 -2.675 -25.060 -1.675 ;
        RECT -24.310 -2.675 -24.080 -1.675 ;
        RECT -23.330 -2.675 -23.100 -1.675 ;
        RECT -21.040 -2.675 -20.810 -1.675 ;
        RECT -20.060 -2.675 -19.830 -1.675 ;
        RECT -19.080 -2.675 -18.850 -1.675 ;
        RECT 136.950 -1.930 159.730 -1.530 ;
        RECT 22.620 -3.385 22.850 -2.385 ;
        RECT 23.600 -3.385 23.830 -2.385 ;
        RECT 24.580 -3.385 24.810 -2.385 ;
        RECT 26.870 -3.385 27.100 -2.385 ;
        RECT 27.850 -3.385 28.080 -2.385 ;
        RECT 28.830 -3.385 29.060 -2.385 ;
        RECT 37.855 -4.495 38.085 -2.495 ;
        RECT 39.035 -4.495 39.265 -2.495 ;
        RECT 40.215 -4.495 40.445 -2.495 ;
        RECT 40.865 -4.495 41.095 -2.495 ;
        RECT 42.045 -4.495 42.275 -2.495 ;
        RECT 43.225 -4.495 43.455 -2.495 ;
        RECT 44.405 -4.495 44.635 -2.495 ;
        RECT 45.585 -4.495 45.815 -2.495 ;
        RECT 46.235 -4.495 46.465 -2.495 ;
        RECT 47.415 -4.495 47.645 -2.495 ;
        RECT 48.595 -4.495 48.825 -2.495 ;
        RECT 49.775 -4.495 50.005 -2.495 ;
        RECT 50.955 -4.495 51.185 -2.495 ;
        RECT 52.135 -4.495 52.365 -2.495 ;
        RECT 53.315 -4.495 53.545 -2.495 ;
        RECT 54.495 -4.495 54.725 -2.495 ;
        RECT 55.675 -4.495 55.905 -2.495 ;
        RECT 56.915 -4.495 57.145 -2.495 ;
        RECT 58.095 -4.495 58.325 -2.495 ;
        RECT 59.275 -4.495 59.505 -2.495 ;
        RECT 60.455 -4.495 60.685 -2.495 ;
        RECT 61.635 -4.495 61.865 -2.495 ;
        RECT 62.815 -4.495 63.045 -2.495 ;
        RECT 63.995 -4.495 64.225 -2.495 ;
        RECT 65.175 -4.495 65.405 -2.495 ;
        RECT 66.355 -4.495 66.585 -2.495 ;
        RECT 67.535 -4.495 67.765 -2.495 ;
        RECT 68.715 -4.495 68.945 -2.495 ;
        RECT 69.895 -4.495 70.125 -2.495 ;
        RECT 71.075 -4.495 71.305 -2.495 ;
        RECT 72.255 -4.495 72.485 -2.495 ;
        RECT 73.435 -4.495 73.665 -2.495 ;
        RECT 74.615 -4.495 74.845 -2.495 ;
        RECT 104.050 -6.235 104.280 -5.235 ;
        RECT 105.030 -6.235 105.260 -5.235 ;
        RECT 106.010 -6.235 106.240 -5.235 ;
        RECT -21.040 -8.050 -20.810 -7.050 ;
        RECT -20.060 -8.050 -19.830 -7.050 ;
        RECT -19.080 -8.050 -18.850 -7.050 ;
        RECT 26.870 -8.760 27.100 -7.760 ;
        RECT 27.850 -8.760 28.080 -7.760 ;
        RECT 28.830 -8.760 29.060 -7.760 ;
        RECT 253.435 -16.620 253.665 -14.620 ;
        RECT 254.615 -16.620 254.845 -14.620 ;
        RECT 255.795 -16.620 256.025 -14.620 ;
        RECT 256.445 -16.620 256.675 -14.620 ;
        RECT 257.625 -16.620 257.855 -14.620 ;
        RECT 258.805 -16.620 259.035 -14.620 ;
        RECT 259.985 -16.620 260.215 -14.620 ;
        RECT 261.165 -16.620 261.395 -14.620 ;
        RECT 261.815 -16.620 262.045 -14.620 ;
        RECT 262.995 -16.620 263.225 -14.620 ;
        RECT 264.175 -16.620 264.405 -14.620 ;
        RECT 265.355 -16.620 265.585 -14.620 ;
        RECT 266.535 -16.620 266.765 -14.620 ;
        RECT 267.715 -16.620 267.945 -14.620 ;
        RECT 268.895 -16.620 269.125 -14.620 ;
        RECT 270.075 -16.620 270.305 -14.620 ;
        RECT 271.255 -16.620 271.485 -14.620 ;
        RECT 272.495 -16.620 272.725 -14.620 ;
        RECT 273.675 -16.620 273.905 -14.620 ;
        RECT 274.855 -16.620 275.085 -14.620 ;
        RECT 276.035 -16.620 276.265 -14.620 ;
        RECT 277.215 -16.620 277.445 -14.620 ;
        RECT 278.395 -16.620 278.625 -14.620 ;
        RECT 279.575 -16.620 279.805 -14.620 ;
        RECT 280.755 -16.620 280.985 -14.620 ;
        RECT 281.935 -16.620 282.165 -14.620 ;
        RECT 283.115 -16.620 283.345 -14.620 ;
        RECT 284.295 -16.620 284.525 -14.620 ;
        RECT 285.475 -16.620 285.705 -14.620 ;
        RECT 286.655 -16.620 286.885 -14.620 ;
        RECT 287.835 -16.620 288.065 -14.620 ;
        RECT 289.015 -16.620 289.245 -14.620 ;
        RECT 290.195 -16.620 290.425 -14.620 ;
        RECT 311.935 -15.190 312.165 -14.190 ;
        RECT 312.915 -15.190 313.145 -14.190 ;
        RECT 313.895 -15.190 314.125 -14.190 ;
        RECT 316.185 -15.190 316.415 -14.190 ;
        RECT 317.165 -15.190 317.395 -14.190 ;
        RECT 318.145 -15.190 318.375 -14.190 ;
        RECT 316.185 -20.565 316.415 -19.565 ;
        RECT 317.165 -20.565 317.395 -19.565 ;
        RECT 318.145 -20.565 318.375 -19.565 ;
        RECT -74.685 -82.680 -74.455 -80.680 ;
        RECT -73.505 -82.680 -73.275 -80.680 ;
        RECT -72.325 -82.680 -72.095 -80.680 ;
        RECT -71.145 -82.680 -70.915 -80.680 ;
        RECT -69.965 -82.680 -69.735 -80.680 ;
        RECT -68.785 -82.680 -68.555 -80.680 ;
        RECT -67.605 -82.680 -67.375 -80.680 ;
        RECT -66.425 -82.680 -66.195 -80.680 ;
        RECT -65.245 -82.680 -65.015 -80.680 ;
        RECT -64.065 -82.680 -63.835 -80.680 ;
        RECT -62.885 -82.680 -62.655 -80.680 ;
        RECT -61.705 -82.680 -61.475 -80.680 ;
        RECT -60.525 -82.680 -60.295 -80.680 ;
        RECT -59.345 -82.680 -59.115 -80.680 ;
        RECT -58.165 -82.680 -57.935 -80.680 ;
        RECT -56.985 -82.680 -56.755 -80.680 ;
        RECT -55.745 -82.680 -55.515 -80.680 ;
        RECT -54.565 -82.680 -54.335 -80.680 ;
        RECT -53.385 -82.680 -53.155 -80.680 ;
        RECT -52.205 -82.680 -51.975 -80.680 ;
        RECT -51.025 -82.680 -50.795 -80.680 ;
        RECT -49.845 -82.680 -49.615 -80.680 ;
        RECT -48.665 -82.680 -48.435 -80.680 ;
        RECT -47.485 -82.680 -47.255 -80.680 ;
        RECT -46.305 -82.680 -46.075 -80.680 ;
        RECT -45.655 -82.680 -45.425 -80.680 ;
        RECT -44.475 -82.680 -44.245 -80.680 ;
        RECT -43.295 -82.680 -43.065 -80.680 ;
        RECT -42.115 -82.680 -41.885 -80.680 ;
        RECT -40.935 -82.680 -40.705 -80.680 ;
        RECT -40.285 -82.680 -40.055 -80.680 ;
        RECT -39.105 -82.680 -38.875 -80.680 ;
        RECT -37.925 -82.680 -37.695 -80.680 ;
        RECT -75.725 -92.985 -75.495 -91.985 ;
        RECT -74.745 -92.985 -74.515 -91.985 ;
        RECT -73.765 -92.985 -73.535 -91.985 ;
        RECT -71.540 -92.985 -71.310 -91.985 ;
        RECT -70.560 -92.985 -70.330 -91.985 ;
        RECT -69.580 -92.985 -69.350 -91.985 ;
        RECT -62.225 -92.985 -61.995 -91.985 ;
        RECT -61.245 -92.985 -61.015 -91.985 ;
        RECT -60.265 -92.985 -60.035 -91.985 ;
        RECT -58.040 -92.985 -57.810 -91.985 ;
        RECT -57.060 -92.985 -56.830 -91.985 ;
        RECT -56.080 -92.985 -55.850 -91.985 ;
        RECT -43.915 -95.035 -43.685 -92.035 ;
        RECT -41.800 -95.035 -41.570 -92.035 ;
        RECT -40.820 -95.035 -40.590 -92.035 ;
        RECT -33.375 -94.015 -33.145 -93.015 ;
        RECT -32.395 -94.015 -32.165 -93.015 ;
        RECT -31.415 -94.015 -31.185 -93.015 ;
        RECT -30.845 -94.015 -30.615 -93.015 ;
        RECT -29.865 -94.015 -29.635 -93.015 ;
        RECT -29.300 -94.015 -29.070 -93.015 ;
        RECT -28.320 -94.015 -28.090 -93.015 ;
        RECT -20.875 -94.015 -20.645 -93.015 ;
        RECT -19.895 -94.015 -19.665 -93.015 ;
        RECT -18.915 -94.015 -18.685 -93.015 ;
        RECT -18.345 -94.015 -18.115 -93.015 ;
        RECT -17.365 -94.015 -17.135 -93.015 ;
        RECT -16.800 -94.015 -16.570 -93.015 ;
        RECT -15.820 -94.015 -15.590 -93.015 ;
        RECT -8.375 -94.015 -8.145 -93.015 ;
        RECT -7.395 -94.015 -7.165 -93.015 ;
        RECT -6.415 -94.015 -6.185 -93.015 ;
        RECT -5.845 -94.015 -5.615 -93.015 ;
        RECT -4.865 -94.015 -4.635 -93.015 ;
        RECT -4.300 -94.015 -4.070 -93.015 ;
        RECT -3.320 -94.015 -3.090 -93.015 ;
        RECT 4.125 -94.015 4.355 -93.015 ;
        RECT 5.105 -94.015 5.335 -93.015 ;
        RECT 6.085 -94.015 6.315 -93.015 ;
        RECT 6.655 -94.015 6.885 -93.015 ;
        RECT 7.635 -94.015 7.865 -93.015 ;
        RECT 8.200 -94.015 8.430 -93.015 ;
        RECT 9.180 -94.015 9.410 -93.015 ;
        RECT 16.625 -94.015 16.855 -93.015 ;
        RECT 17.605 -94.015 17.835 -93.015 ;
        RECT 18.585 -94.015 18.815 -93.015 ;
        RECT 19.155 -94.015 19.385 -93.015 ;
        RECT 20.135 -94.015 20.365 -93.015 ;
        RECT 20.700 -94.015 20.930 -93.015 ;
        RECT 21.680 -94.015 21.910 -93.015 ;
        RECT 31.625 -94.015 31.855 -93.015 ;
        RECT 32.605 -94.015 32.835 -93.015 ;
        RECT 33.585 -94.015 33.815 -93.015 ;
        RECT 34.155 -94.015 34.385 -93.015 ;
        RECT 35.135 -94.015 35.365 -93.015 ;
        RECT 35.700 -94.015 35.930 -93.015 ;
        RECT 36.680 -94.015 36.910 -93.015 ;
        RECT -113.720 -96.920 -113.490 -95.920 ;
        RECT -112.740 -96.920 -112.510 -95.920 ;
        RECT -111.760 -96.920 -111.530 -95.920 ;
        RECT -110.780 -96.920 -110.550 -95.920 ;
        RECT -108.070 -96.920 -107.840 -95.920 ;
        RECT -107.090 -96.920 -106.860 -95.920 ;
        RECT -103.725 -98.030 -103.495 -96.530 ;
        RECT -102.745 -98.030 -102.515 -96.530 ;
        RECT -101.765 -98.030 -101.535 -96.530 ;
        RECT -100.680 -97.025 -100.450 -96.525 ;
        RECT -99.700 -97.025 -99.470 -96.525 ;
        RECT -98.720 -97.025 -98.490 -96.525 ;
        RECT -97.740 -97.025 -97.510 -96.525 ;
        RECT -26.735 -96.805 -26.120 -96.125 ;
        RECT -75.235 -99.575 -75.005 -98.575 ;
        RECT -74.255 -99.575 -74.025 -98.575 ;
        RECT -73.275 -99.575 -73.045 -98.575 ;
        RECT -66.520 -99.575 -66.290 -98.575 ;
        RECT -65.540 -99.575 -65.310 -98.575 ;
        RECT -64.560 -99.575 -64.330 -98.575 ;
        RECT -61.735 -99.575 -61.505 -98.575 ;
        RECT -60.755 -99.575 -60.525 -98.575 ;
        RECT -59.775 -99.575 -59.545 -98.575 ;
        RECT -53.020 -99.575 -52.790 -98.575 ;
        RECT -52.040 -99.575 -51.810 -98.575 ;
        RECT -51.060 -99.575 -50.830 -98.575 ;
        RECT -48.610 -99.575 -48.380 -98.575 ;
        RECT -47.630 -99.575 -47.400 -98.575 ;
        RECT -46.650 -99.575 -46.420 -98.575 ;
        RECT -95.545 -102.840 -95.315 -101.340 ;
        RECT -94.565 -102.840 -94.335 -101.340 ;
        RECT -93.585 -102.840 -93.355 -101.340 ;
        RECT -92.500 -102.845 -92.270 -102.345 ;
        RECT -91.520 -102.845 -91.290 -102.345 ;
        RECT -90.540 -102.845 -90.310 -102.345 ;
        RECT -89.560 -102.845 -89.330 -102.345 ;
        RECT -88.310 -103.285 -88.080 -100.285 ;
        RECT -87.330 -103.285 -87.100 -100.285 ;
        RECT -85.215 -103.285 -84.985 -100.285 ;
        RECT -35.070 -100.660 -34.840 -99.660 ;
        RECT -34.090 -100.660 -33.860 -99.660 ;
        RECT -33.110 -100.660 -32.880 -99.660 ;
        RECT -26.715 -99.960 -26.145 -96.805 ;
        RECT -13.900 -96.980 -13.285 -96.300 ;
        RECT -1.485 -96.980 -0.870 -96.300 ;
        RECT -13.880 -99.240 -13.310 -96.980 ;
        RECT -1.465 -99.065 -0.895 -96.980 ;
        RECT -1.490 -99.070 -0.875 -99.065 ;
        RECT -13.905 -99.920 -13.290 -99.240 ;
        RECT -1.490 -99.380 0.040 -99.070 ;
        RECT -26.740 -100.640 -26.125 -99.960 ;
        RECT 16.835 -103.275 17.450 -103.230 ;
        RECT 18.840 -103.275 19.455 -103.220 ;
        RECT -7.610 -103.350 -6.995 -103.290 ;
        RECT -6.140 -103.350 -5.525 -103.285 ;
        RECT -7.610 -103.925 -5.525 -103.350 ;
        RECT -7.610 -103.970 -6.995 -103.925 ;
        RECT -6.140 -103.965 -5.525 -103.925 ;
        RECT 8.750 -103.425 9.365 -103.350 ;
        RECT 10.695 -103.425 11.310 -103.345 ;
        RECT 8.750 -103.960 11.310 -103.425 ;
        RECT 16.835 -103.810 19.455 -103.275 ;
        RECT 16.835 -103.910 17.450 -103.810 ;
        RECT 18.840 -103.900 19.455 -103.810 ;
        RECT 25.620 -103.310 26.235 -103.245 ;
        RECT 31.700 -103.310 32.315 -103.250 ;
        RECT 25.620 -103.835 32.315 -103.310 ;
        RECT 25.620 -103.925 26.235 -103.835 ;
        RECT 31.700 -103.930 32.315 -103.835 ;
        RECT 8.750 -104.030 9.365 -103.960 ;
        RECT 10.695 -104.025 11.310 -103.960 ;
        RECT -113.435 -107.575 -113.205 -106.075 ;
        RECT -112.455 -107.575 -112.225 -106.075 ;
        RECT -111.475 -107.575 -111.245 -106.075 ;
        RECT -110.390 -106.570 -110.160 -106.070 ;
        RECT -109.410 -106.570 -109.180 -106.070 ;
        RECT -108.430 -106.570 -108.200 -106.070 ;
        RECT -107.450 -106.570 -107.220 -106.070 ;
        RECT -104.570 -106.600 -104.340 -105.600 ;
        RECT -103.590 -106.600 -103.360 -105.600 ;
        RECT -102.610 -106.600 -102.380 -105.600 ;
        RECT -101.630 -106.600 -101.400 -105.600 ;
        RECT -98.920 -106.600 -98.690 -105.600 ;
        RECT -97.940 -106.600 -97.710 -105.600 ;
        RECT -95.415 -107.485 -95.185 -106.485 ;
        RECT -94.435 -107.485 -94.205 -106.485 ;
        RECT -93.455 -107.485 -93.225 -106.485 ;
        RECT -92.475 -107.485 -92.245 -106.485 ;
        RECT -90.550 -107.340 -90.320 -105.840 ;
        RECT -89.570 -107.340 -89.340 -105.840 ;
        RECT -88.590 -107.340 -88.360 -105.840 ;
        RECT -87.505 -106.335 -87.275 -105.835 ;
        RECT -86.525 -106.335 -86.295 -105.835 ;
        RECT -85.545 -106.335 -85.315 -105.835 ;
        RECT -84.565 -106.335 -84.335 -105.835 ;
        RECT -70.600 -107.720 -70.370 -106.220 ;
        RECT -69.620 -107.720 -69.390 -106.220 ;
        RECT -68.640 -107.720 -68.410 -106.220 ;
        RECT -67.555 -107.725 -67.325 -107.225 ;
        RECT -66.575 -107.725 -66.345 -107.225 ;
        RECT -65.595 -107.725 -65.365 -107.225 ;
        RECT -64.615 -107.725 -64.385 -107.225 ;
        RECT -63.365 -108.165 -63.135 -105.165 ;
        RECT -62.385 -108.165 -62.155 -105.165 ;
        RECT -60.270 -108.165 -60.040 -105.165 ;
        RECT -35.865 -105.175 -35.635 -104.175 ;
        RECT -34.885 -105.175 -34.655 -104.175 ;
        RECT -33.905 -105.175 -33.675 -104.175 ;
        RECT -27.150 -105.175 -26.920 -104.175 ;
        RECT -26.170 -105.175 -25.940 -104.175 ;
        RECT -25.190 -105.175 -24.960 -104.175 ;
        RECT -22.365 -105.175 -22.135 -104.175 ;
        RECT -21.385 -105.175 -21.155 -104.175 ;
        RECT -20.405 -105.175 -20.175 -104.175 ;
        RECT -13.650 -105.175 -13.420 -104.175 ;
        RECT -12.670 -105.175 -12.440 -104.175 ;
        RECT -11.690 -105.175 -11.460 -104.175 ;
        RECT -9.240 -105.175 -9.010 -104.175 ;
        RECT -8.260 -105.175 -8.030 -104.175 ;
        RECT -7.280 -105.175 -7.050 -104.175 ;
        RECT -5.570 -105.260 -5.340 -104.260 ;
        RECT -4.590 -105.260 -4.360 -104.260 ;
        RECT -1.880 -105.260 -1.650 -104.260 ;
        RECT -0.900 -105.260 -0.670 -104.260 ;
        RECT 0.080 -105.260 0.310 -104.260 ;
        RECT 1.060 -105.260 1.290 -104.260 ;
        RECT 3.095 -104.825 3.325 -104.325 ;
        RECT 4.075 -104.825 4.305 -104.325 ;
        RECT 5.055 -104.825 5.285 -104.325 ;
        RECT 6.035 -104.825 6.265 -104.325 ;
        RECT 7.120 -105.830 7.350 -104.330 ;
        RECT 8.100 -105.830 8.330 -104.330 ;
        RECT 9.080 -105.830 9.310 -104.330 ;
        RECT 11.120 -104.835 11.350 -104.335 ;
        RECT 12.100 -104.835 12.330 -104.335 ;
        RECT 13.080 -104.835 13.310 -104.335 ;
        RECT 14.060 -104.835 14.290 -104.335 ;
        RECT 15.145 -105.840 15.375 -104.340 ;
        RECT 16.125 -105.840 16.355 -104.340 ;
        RECT 17.105 -105.840 17.335 -104.340 ;
        RECT 19.240 -105.215 19.470 -104.215 ;
        RECT 20.220 -105.215 20.450 -104.215 ;
        RECT 22.930 -105.215 23.160 -104.215 ;
        RECT 23.910 -105.215 24.140 -104.215 ;
        RECT 24.890 -105.215 25.120 -104.215 ;
        RECT 25.870 -105.215 26.100 -104.215 ;
        RECT 31.675 -105.270 31.905 -104.270 ;
        RECT 32.655 -105.270 32.885 -104.270 ;
        RECT 33.635 -105.270 33.865 -104.270 ;
        RECT 34.205 -105.270 34.435 -104.270 ;
        RECT 35.185 -105.270 35.415 -104.270 ;
        RECT 35.750 -105.270 35.980 -104.270 ;
        RECT 36.730 -105.270 36.960 -104.270 ;
        RECT 134.760 -104.755 134.990 -103.755 ;
        RECT 135.740 -104.755 135.970 -103.755 ;
        RECT 136.720 -104.755 136.950 -103.755 ;
        RECT 137.700 -104.755 137.930 -103.755 ;
        RECT 139.625 -105.400 139.855 -103.900 ;
        RECT 140.605 -105.400 140.835 -103.900 ;
        RECT 141.585 -105.400 141.815 -103.900 ;
        RECT 176.960 -104.810 177.190 -103.810 ;
        RECT 177.940 -104.810 178.170 -103.810 ;
        RECT 178.920 -104.810 179.150 -103.810 ;
        RECT 179.900 -104.810 180.130 -103.810 ;
        RECT 142.670 -105.405 142.900 -104.905 ;
        RECT 143.650 -105.405 143.880 -104.905 ;
        RECT 144.630 -105.405 144.860 -104.905 ;
        RECT 145.610 -105.405 145.840 -104.905 ;
        RECT 181.825 -105.455 182.055 -103.955 ;
        RECT 182.805 -105.455 183.035 -103.955 ;
        RECT 183.785 -105.455 184.015 -103.955 ;
        RECT 184.870 -105.460 185.100 -104.960 ;
        RECT 185.850 -105.460 186.080 -104.960 ;
        RECT 186.830 -105.460 187.060 -104.960 ;
        RECT 187.810 -105.460 188.040 -104.960 ;
        RECT 221.275 -105.005 221.505 -104.005 ;
        RECT 222.255 -105.005 222.485 -104.005 ;
        RECT 223.235 -105.005 223.465 -104.005 ;
        RECT 224.215 -105.005 224.445 -104.005 ;
        RECT 102.900 -106.520 103.130 -105.520 ;
        RECT 103.880 -106.520 104.110 -105.520 ;
        RECT 104.860 -106.520 105.090 -105.520 ;
        RECT 107.085 -106.520 107.315 -105.520 ;
        RECT 108.065 -106.520 108.295 -105.520 ;
        RECT 109.045 -106.520 109.275 -105.520 ;
        RECT 116.400 -106.520 116.630 -105.520 ;
        RECT 117.380 -106.520 117.610 -105.520 ;
        RECT 118.360 -106.520 118.590 -105.520 ;
        RECT 120.585 -106.520 120.815 -105.520 ;
        RECT 121.565 -106.520 121.795 -105.520 ;
        RECT 122.545 -106.520 122.775 -105.520 ;
        RECT 226.140 -105.650 226.370 -104.150 ;
        RECT 227.120 -105.650 227.350 -104.150 ;
        RECT 228.100 -105.650 228.330 -104.150 ;
        RECT 267.265 -104.835 267.495 -103.835 ;
        RECT 268.245 -104.835 268.475 -103.835 ;
        RECT 269.225 -104.835 269.455 -103.835 ;
        RECT 270.205 -104.835 270.435 -103.835 ;
        RECT 229.185 -105.655 229.415 -105.155 ;
        RECT 230.165 -105.655 230.395 -105.155 ;
        RECT 231.145 -105.655 231.375 -105.155 ;
        RECT 232.125 -105.655 232.355 -105.155 ;
        RECT 272.130 -105.480 272.360 -103.980 ;
        RECT 273.110 -105.480 273.340 -103.980 ;
        RECT 274.090 -105.480 274.320 -103.980 ;
        RECT 311.035 -104.505 311.265 -103.505 ;
        RECT 312.015 -104.505 312.245 -103.505 ;
        RECT 312.995 -104.505 313.225 -103.505 ;
        RECT 313.975 -104.505 314.205 -103.505 ;
        RECT 275.175 -105.485 275.405 -104.985 ;
        RECT 276.155 -105.485 276.385 -104.985 ;
        RECT 277.135 -105.485 277.365 -104.985 ;
        RECT 278.115 -105.485 278.345 -104.985 ;
        RECT 315.900 -105.150 316.130 -103.650 ;
        RECT 316.880 -105.150 317.110 -103.650 ;
        RECT 317.860 -105.150 318.090 -103.650 ;
        RECT 356.800 -104.420 357.030 -103.420 ;
        RECT 357.780 -104.420 358.010 -103.420 ;
        RECT 358.760 -104.420 358.990 -103.420 ;
        RECT 359.740 -104.420 359.970 -103.420 ;
        RECT 318.945 -105.155 319.175 -104.655 ;
        RECT 319.925 -105.155 320.155 -104.655 ;
        RECT 320.905 -105.155 321.135 -104.655 ;
        RECT 321.885 -105.155 322.115 -104.655 ;
        RECT 361.665 -105.065 361.895 -103.565 ;
        RECT 362.645 -105.065 362.875 -103.565 ;
        RECT 363.625 -105.065 363.855 -103.565 ;
        RECT 403.620 -104.230 403.850 -103.230 ;
        RECT 404.600 -104.230 404.830 -103.230 ;
        RECT 405.580 -104.230 405.810 -103.230 ;
        RECT 406.560 -104.230 406.790 -103.230 ;
        RECT 364.710 -105.070 364.940 -104.570 ;
        RECT 365.690 -105.070 365.920 -104.570 ;
        RECT 366.670 -105.070 366.900 -104.570 ;
        RECT 367.650 -105.070 367.880 -104.570 ;
        RECT 408.485 -104.875 408.715 -103.375 ;
        RECT 409.465 -104.875 409.695 -103.375 ;
        RECT 410.445 -104.875 410.675 -103.375 ;
        RECT 411.530 -104.880 411.760 -104.380 ;
        RECT 412.510 -104.880 412.740 -104.380 ;
        RECT 413.490 -104.880 413.720 -104.380 ;
        RECT 414.470 -104.880 414.700 -104.380 ;
        RECT 414.880 -106.455 415.250 -106.375 ;
        RECT 416.020 -106.455 416.570 -106.275 ;
        RECT 322.295 -106.730 322.665 -106.650 ;
        RECT 323.435 -106.730 323.985 -106.550 ;
        RECT 146.020 -106.980 146.390 -106.900 ;
        RECT 147.160 -106.980 147.710 -106.800 ;
        RECT 146.020 -107.460 147.710 -106.980 ;
        RECT 188.220 -107.035 188.590 -106.955 ;
        RECT 189.360 -107.035 189.910 -106.855 ;
        RECT 146.020 -107.490 146.390 -107.460 ;
        RECT 147.160 -107.550 147.710 -107.460 ;
        RECT -70.470 -112.365 -70.240 -111.365 ;
        RECT -69.490 -112.365 -69.260 -111.365 ;
        RECT -68.510 -112.365 -68.280 -111.365 ;
        RECT -67.530 -112.365 -67.300 -111.365 ;
        RECT -65.605 -112.220 -65.375 -110.720 ;
        RECT -64.625 -112.220 -64.395 -110.720 ;
        RECT -63.645 -112.220 -63.415 -110.720 ;
        RECT -62.560 -111.215 -62.330 -110.715 ;
        RECT -61.580 -111.215 -61.350 -110.715 ;
        RECT -60.600 -111.215 -60.370 -110.715 ;
        RECT -59.620 -111.215 -59.390 -110.715 ;
        RECT -36.355 -111.765 -36.125 -110.765 ;
        RECT -35.375 -111.765 -35.145 -110.765 ;
        RECT -34.395 -111.765 -34.165 -110.765 ;
        RECT -32.170 -111.765 -31.940 -110.765 ;
        RECT -31.190 -111.765 -30.960 -110.765 ;
        RECT -30.210 -111.765 -29.980 -110.765 ;
        RECT -22.855 -111.765 -22.625 -110.765 ;
        RECT -21.875 -111.765 -21.645 -110.765 ;
        RECT -20.895 -111.765 -20.665 -110.765 ;
        RECT -18.670 -111.765 -18.440 -110.765 ;
        RECT -17.690 -111.765 -17.460 -110.765 ;
        RECT -16.710 -111.765 -16.480 -110.765 ;
        RECT 86.865 -112.510 87.095 -109.510 ;
        RECT 87.845 -112.510 88.075 -109.510 ;
        RECT 134.630 -109.900 134.860 -108.400 ;
        RECT 135.610 -109.900 135.840 -108.400 ;
        RECT 136.590 -109.900 136.820 -108.400 ;
        RECT 137.675 -108.895 137.905 -108.395 ;
        RECT 138.655 -108.895 138.885 -108.395 ;
        RECT 139.635 -108.895 139.865 -108.395 ;
        RECT 140.615 -108.895 140.845 -108.395 ;
        RECT 141.865 -110.955 142.095 -107.955 ;
        RECT 142.845 -110.955 143.075 -107.955 ;
        RECT 144.960 -110.955 145.190 -107.955 ;
        RECT 151.825 -109.745 152.055 -107.245 ;
        RECT 152.805 -109.745 153.035 -107.245 ;
        RECT 155.780 -109.745 156.010 -107.245 ;
        RECT 156.430 -109.745 156.660 -107.245 ;
        RECT 157.570 -108.745 157.800 -107.245 ;
        RECT 158.550 -108.745 158.780 -107.245 ;
        RECT 188.220 -107.515 189.910 -107.035 ;
        RECT 232.535 -107.230 232.905 -107.150 ;
        RECT 233.675 -107.230 234.225 -107.050 ;
        RECT 188.220 -107.545 188.590 -107.515 ;
        RECT 189.360 -107.605 189.910 -107.515 ;
        RECT 176.830 -109.955 177.060 -108.455 ;
        RECT 177.810 -109.955 178.040 -108.455 ;
        RECT 178.790 -109.955 179.020 -108.455 ;
        RECT 179.875 -108.950 180.105 -108.450 ;
        RECT 180.855 -108.950 181.085 -108.450 ;
        RECT 181.835 -108.950 182.065 -108.450 ;
        RECT 182.815 -108.950 183.045 -108.450 ;
        RECT 184.065 -111.010 184.295 -108.010 ;
        RECT 185.045 -111.010 185.275 -108.010 ;
        RECT 187.160 -111.010 187.390 -108.010 ;
        RECT 194.025 -109.800 194.255 -107.300 ;
        RECT 195.005 -109.800 195.235 -107.300 ;
        RECT 197.980 -109.800 198.210 -107.300 ;
        RECT 198.630 -109.800 198.860 -107.300 ;
        RECT 199.770 -108.800 200.000 -107.300 ;
        RECT 200.750 -108.800 200.980 -107.300 ;
        RECT 232.535 -107.710 234.225 -107.230 ;
        RECT 278.525 -107.060 278.895 -106.980 ;
        RECT 279.665 -107.060 280.215 -106.880 ;
        RECT 232.535 -107.740 232.905 -107.710 ;
        RECT 233.675 -107.800 234.225 -107.710 ;
        RECT 221.145 -110.150 221.375 -108.650 ;
        RECT 222.125 -110.150 222.355 -108.650 ;
        RECT 223.105 -110.150 223.335 -108.650 ;
        RECT 224.190 -109.145 224.420 -108.645 ;
        RECT 225.170 -109.145 225.400 -108.645 ;
        RECT 226.150 -109.145 226.380 -108.645 ;
        RECT 227.130 -109.145 227.360 -108.645 ;
        RECT 228.380 -111.205 228.610 -108.205 ;
        RECT 229.360 -111.205 229.590 -108.205 ;
        RECT 231.475 -111.205 231.705 -108.205 ;
        RECT 238.340 -109.995 238.570 -107.495 ;
        RECT 239.320 -109.995 239.550 -107.495 ;
        RECT 242.295 -109.995 242.525 -107.495 ;
        RECT 242.945 -109.995 243.175 -107.495 ;
        RECT 244.085 -108.995 244.315 -107.495 ;
        RECT 245.065 -108.995 245.295 -107.495 ;
        RECT 278.525 -107.540 280.215 -107.060 ;
        RECT 322.295 -107.210 323.985 -106.730 ;
        RECT 368.060 -106.645 368.430 -106.565 ;
        RECT 369.200 -106.645 369.750 -106.465 ;
        RECT 322.295 -107.240 322.665 -107.210 ;
        RECT 323.435 -107.300 323.985 -107.210 ;
        RECT 278.525 -107.570 278.895 -107.540 ;
        RECT 279.665 -107.630 280.215 -107.540 ;
        RECT 267.135 -109.980 267.365 -108.480 ;
        RECT 268.115 -109.980 268.345 -108.480 ;
        RECT 269.095 -109.980 269.325 -108.480 ;
        RECT 270.180 -108.975 270.410 -108.475 ;
        RECT 271.160 -108.975 271.390 -108.475 ;
        RECT 272.140 -108.975 272.370 -108.475 ;
        RECT 273.120 -108.975 273.350 -108.475 ;
        RECT 274.370 -111.035 274.600 -108.035 ;
        RECT 275.350 -111.035 275.580 -108.035 ;
        RECT 277.465 -111.035 277.695 -108.035 ;
        RECT 284.330 -109.825 284.560 -107.325 ;
        RECT 285.310 -109.825 285.540 -107.325 ;
        RECT 288.285 -109.825 288.515 -107.325 ;
        RECT 288.935 -109.825 289.165 -107.325 ;
        RECT 290.075 -108.825 290.305 -107.325 ;
        RECT 291.055 -108.825 291.285 -107.325 ;
        RECT 310.905 -109.650 311.135 -108.150 ;
        RECT 311.885 -109.650 312.115 -108.150 ;
        RECT 312.865 -109.650 313.095 -108.150 ;
        RECT 313.950 -108.645 314.180 -108.145 ;
        RECT 314.930 -108.645 315.160 -108.145 ;
        RECT 315.910 -108.645 316.140 -108.145 ;
        RECT 316.890 -108.645 317.120 -108.145 ;
        RECT 318.140 -110.705 318.370 -107.705 ;
        RECT 319.120 -110.705 319.350 -107.705 ;
        RECT 321.235 -110.705 321.465 -107.705 ;
        RECT 328.100 -109.495 328.330 -106.995 ;
        RECT 329.080 -109.495 329.310 -106.995 ;
        RECT 332.055 -109.495 332.285 -106.995 ;
        RECT 332.705 -109.495 332.935 -106.995 ;
        RECT 333.845 -108.495 334.075 -106.995 ;
        RECT 334.825 -108.495 335.055 -106.995 ;
        RECT 368.060 -107.125 369.750 -106.645 ;
        RECT 368.060 -107.155 368.430 -107.125 ;
        RECT 369.200 -107.215 369.750 -107.125 ;
        RECT 356.670 -109.565 356.900 -108.065 ;
        RECT 357.650 -109.565 357.880 -108.065 ;
        RECT 358.630 -109.565 358.860 -108.065 ;
        RECT 359.715 -108.560 359.945 -108.060 ;
        RECT 360.695 -108.560 360.925 -108.060 ;
        RECT 361.675 -108.560 361.905 -108.060 ;
        RECT 362.655 -108.560 362.885 -108.060 ;
        RECT 363.905 -110.620 364.135 -107.620 ;
        RECT 364.885 -110.620 365.115 -107.620 ;
        RECT 367.000 -110.620 367.230 -107.620 ;
        RECT 373.865 -109.410 374.095 -106.910 ;
        RECT 374.845 -109.410 375.075 -106.910 ;
        RECT 377.820 -109.410 378.050 -106.910 ;
        RECT 378.470 -109.410 378.700 -106.910 ;
        RECT 379.610 -108.410 379.840 -106.910 ;
        RECT 380.590 -108.410 380.820 -106.910 ;
        RECT 414.880 -106.935 416.570 -106.455 ;
        RECT 414.880 -106.965 415.250 -106.935 ;
        RECT 416.020 -107.025 416.570 -106.935 ;
        RECT 403.490 -109.375 403.720 -107.875 ;
        RECT 404.470 -109.375 404.700 -107.875 ;
        RECT 405.450 -109.375 405.680 -107.875 ;
        RECT 406.535 -108.370 406.765 -107.870 ;
        RECT 407.515 -108.370 407.745 -107.870 ;
        RECT 408.495 -108.370 408.725 -107.870 ;
        RECT 409.475 -108.370 409.705 -107.870 ;
        RECT 410.725 -110.430 410.955 -107.430 ;
        RECT 411.705 -110.430 411.935 -107.430 ;
        RECT 413.820 -110.430 414.050 -107.430 ;
        RECT 420.685 -109.220 420.915 -106.720 ;
        RECT 421.665 -109.220 421.895 -106.720 ;
        RECT 424.640 -109.220 424.870 -106.720 ;
        RECT 425.290 -109.220 425.520 -106.720 ;
        RECT 426.430 -108.220 426.660 -106.720 ;
        RECT 427.410 -108.220 427.640 -106.720 ;
        RECT 93.470 -113.110 93.700 -112.110 ;
        RECT 94.450 -113.110 94.680 -112.110 ;
        RECT 95.430 -113.110 95.660 -112.110 ;
        RECT 97.880 -113.110 98.110 -112.110 ;
        RECT 98.860 -113.110 99.090 -112.110 ;
        RECT 99.840 -113.110 100.070 -112.110 ;
        RECT 106.595 -113.110 106.825 -112.110 ;
        RECT 107.575 -113.110 107.805 -112.110 ;
        RECT 108.555 -113.110 108.785 -112.110 ;
        RECT 111.380 -113.110 111.610 -112.110 ;
        RECT 112.360 -113.110 112.590 -112.110 ;
        RECT 113.340 -113.110 113.570 -112.110 ;
        RECT 120.095 -113.110 120.325 -112.110 ;
        RECT 121.075 -113.110 121.305 -112.110 ;
        RECT 122.055 -113.110 122.285 -112.110 ;
        RECT -75.725 -117.620 -75.495 -116.620 ;
        RECT -74.745 -117.620 -74.515 -116.620 ;
        RECT -73.765 -117.620 -73.535 -116.620 ;
        RECT -71.540 -117.620 -71.310 -116.620 ;
        RECT -70.560 -117.620 -70.330 -116.620 ;
        RECT -69.580 -117.620 -69.350 -116.620 ;
        RECT -62.225 -117.620 -61.995 -116.620 ;
        RECT -61.245 -117.620 -61.015 -116.620 ;
        RECT -60.265 -117.620 -60.035 -116.620 ;
        RECT -58.040 -117.620 -57.810 -116.620 ;
        RECT -57.060 -117.620 -56.830 -116.620 ;
        RECT -56.080 -117.620 -55.850 -116.620 ;
        RECT -97.850 -120.145 -96.955 -119.310 ;
        RECT -43.780 -119.705 -43.550 -116.705 ;
        RECT -41.665 -119.705 -41.435 -116.705 ;
        RECT -40.685 -119.705 -40.455 -116.705 ;
        RECT 105.695 -117.870 105.925 -115.870 ;
        RECT 106.675 -117.870 106.905 -115.870 ;
        RECT 107.655 -117.870 107.885 -115.870 ;
        RECT -36.355 -118.955 -36.125 -117.955 ;
        RECT -35.375 -118.955 -35.145 -117.955 ;
        RECT -34.395 -118.955 -34.165 -117.955 ;
        RECT -32.170 -118.955 -31.940 -117.955 ;
        RECT -31.190 -118.955 -30.960 -117.955 ;
        RECT -30.210 -118.955 -29.980 -117.955 ;
        RECT -22.855 -118.955 -22.625 -117.955 ;
        RECT -21.875 -118.955 -21.645 -117.955 ;
        RECT -20.895 -118.955 -20.665 -117.955 ;
        RECT -18.670 -118.955 -18.440 -117.955 ;
        RECT -17.690 -118.955 -17.460 -117.955 ;
        RECT -16.710 -118.955 -16.480 -117.955 ;
        RECT -113.110 -125.045 -112.880 -122.045 ;
        RECT -112.130 -125.045 -111.900 -122.045 ;
        RECT -107.080 -123.690 -106.850 -121.690 ;
        RECT -106.100 -123.690 -105.870 -121.690 ;
        RECT -102.555 -123.695 -102.325 -121.695 ;
        RECT -101.575 -123.695 -101.345 -121.695 ;
        RECT -97.715 -128.965 -97.085 -120.145 ;
        RECT -75.235 -124.210 -75.005 -123.210 ;
        RECT -74.255 -124.210 -74.025 -123.210 ;
        RECT -73.275 -124.210 -73.045 -123.210 ;
        RECT -66.520 -124.210 -66.290 -123.210 ;
        RECT -65.540 -124.210 -65.310 -123.210 ;
        RECT -64.560 -124.210 -64.330 -123.210 ;
        RECT -61.735 -124.210 -61.505 -123.210 ;
        RECT -60.755 -124.210 -60.525 -123.210 ;
        RECT -59.775 -124.210 -59.545 -123.210 ;
        RECT -53.020 -124.210 -52.790 -123.210 ;
        RECT -52.040 -124.210 -51.810 -123.210 ;
        RECT -51.060 -124.210 -50.830 -123.210 ;
        RECT -48.610 -124.210 -48.380 -123.210 ;
        RECT -47.630 -124.210 -47.400 -123.210 ;
        RECT -46.650 -124.210 -46.420 -123.210 ;
        RECT -95.545 -127.840 -95.315 -126.340 ;
        RECT -94.565 -127.840 -94.335 -126.340 ;
        RECT -93.585 -127.840 -93.355 -126.340 ;
        RECT -92.500 -127.845 -92.270 -127.345 ;
        RECT -91.520 -127.845 -91.290 -127.345 ;
        RECT -90.540 -127.845 -90.310 -127.345 ;
        RECT -89.560 -127.845 -89.330 -127.345 ;
        RECT -88.310 -128.285 -88.080 -125.285 ;
        RECT -87.330 -128.285 -87.100 -125.285 ;
        RECT -85.215 -128.285 -84.985 -125.285 ;
        RECT -35.865 -125.545 -35.635 -124.545 ;
        RECT -34.885 -125.545 -34.655 -124.545 ;
        RECT -33.905 -125.545 -33.675 -124.545 ;
        RECT -27.150 -125.545 -26.920 -124.545 ;
        RECT -26.170 -125.545 -25.940 -124.545 ;
        RECT -25.190 -125.545 -24.960 -124.545 ;
        RECT -22.365 -125.545 -22.135 -124.545 ;
        RECT -21.385 -125.545 -21.155 -124.545 ;
        RECT -20.405 -125.545 -20.175 -124.545 ;
        RECT -13.650 -125.545 -13.420 -124.545 ;
        RECT -12.670 -125.545 -12.440 -124.545 ;
        RECT -11.690 -125.545 -11.460 -124.545 ;
        RECT -9.240 -125.545 -9.010 -124.545 ;
        RECT -8.260 -125.545 -8.030 -124.545 ;
        RECT -7.280 -125.545 -7.050 -124.545 ;
        RECT -5.570 -125.460 -5.340 -124.460 ;
        RECT -4.590 -125.460 -4.360 -124.460 ;
        RECT -1.880 -125.460 -1.650 -124.460 ;
        RECT -0.900 -125.460 -0.670 -124.460 ;
        RECT 0.080 -125.460 0.310 -124.460 ;
        RECT 1.060 -125.460 1.290 -124.460 ;
        RECT 3.095 -125.395 3.325 -124.895 ;
        RECT 4.075 -125.395 4.305 -124.895 ;
        RECT 5.055 -125.395 5.285 -124.895 ;
        RECT 6.035 -125.395 6.265 -124.895 ;
        RECT 7.120 -125.390 7.350 -123.890 ;
        RECT 8.100 -125.390 8.330 -123.890 ;
        RECT 9.080 -125.390 9.310 -123.890 ;
        RECT 11.120 -125.385 11.350 -124.885 ;
        RECT 12.100 -125.385 12.330 -124.885 ;
        RECT 13.080 -125.385 13.310 -124.885 ;
        RECT 14.060 -125.385 14.290 -124.885 ;
        RECT 15.145 -125.380 15.375 -123.880 ;
        RECT 16.125 -125.380 16.355 -123.880 ;
        RECT 17.105 -125.380 17.335 -123.880 ;
        RECT 86.840 -124.240 87.070 -122.240 ;
        RECT 87.820 -124.240 88.050 -122.240 ;
        RECT 91.570 -124.240 91.800 -122.240 ;
        RECT 92.550 -124.240 92.780 -122.240 ;
        RECT 96.150 -124.410 96.380 -123.410 ;
        RECT 97.130 -124.410 97.360 -123.410 ;
        RECT 98.110 -124.410 98.340 -123.410 ;
        RECT 99.090 -124.410 99.320 -123.410 ;
        RECT 101.800 -124.410 102.030 -123.410 ;
        RECT 102.780 -124.410 103.010 -123.410 ;
        RECT 105.445 -124.375 105.675 -123.375 ;
        RECT 106.425 -124.375 106.655 -123.375 ;
        RECT 107.405 -124.375 107.635 -123.375 ;
        RECT 109.845 -124.020 110.075 -120.520 ;
        RECT 110.825 -124.020 111.055 -120.520 ;
        RECT 111.845 -124.020 112.075 -120.520 ;
        RECT 112.825 -124.020 113.055 -120.520 ;
        RECT 114.845 -124.020 115.075 -120.520 ;
        RECT 115.825 -124.020 116.055 -120.520 ;
        RECT 116.845 -124.020 117.075 -120.520 ;
        RECT 117.825 -124.020 118.055 -120.520 ;
        RECT 119.845 -124.020 120.075 -120.520 ;
        RECT 120.825 -124.020 121.055 -120.520 ;
        RECT 121.845 -124.020 122.075 -120.520 ;
        RECT 122.825 -124.020 123.055 -120.520 ;
        RECT 134.720 -122.020 134.950 -121.020 ;
        RECT 135.700 -122.020 135.930 -121.020 ;
        RECT 136.680 -122.020 136.910 -121.020 ;
        RECT 137.660 -122.020 137.890 -121.020 ;
        RECT 139.585 -122.665 139.815 -121.165 ;
        RECT 140.565 -122.665 140.795 -121.165 ;
        RECT 141.545 -122.665 141.775 -121.165 ;
        RECT 142.630 -122.670 142.860 -122.170 ;
        RECT 143.610 -122.670 143.840 -122.170 ;
        RECT 144.590 -122.670 144.820 -122.170 ;
        RECT 145.570 -122.670 145.800 -122.170 ;
        RECT 153.060 -122.175 153.290 -121.175 ;
        RECT 154.040 -122.175 154.270 -121.175 ;
        RECT 155.020 -122.175 155.250 -121.175 ;
        RECT 156.000 -122.175 156.230 -121.175 ;
        RECT 157.925 -122.820 158.155 -121.320 ;
        RECT 158.905 -122.820 159.135 -121.320 ;
        RECT 159.885 -122.820 160.115 -121.320 ;
        RECT 176.920 -122.075 177.150 -121.075 ;
        RECT 177.900 -122.075 178.130 -121.075 ;
        RECT 178.880 -122.075 179.110 -121.075 ;
        RECT 179.860 -122.075 180.090 -121.075 ;
        RECT 160.970 -122.825 161.200 -122.325 ;
        RECT 161.950 -122.825 162.180 -122.325 ;
        RECT 162.930 -122.825 163.160 -122.325 ;
        RECT 163.910 -122.825 164.140 -122.325 ;
        RECT 181.785 -122.720 182.015 -121.220 ;
        RECT 182.765 -122.720 182.995 -121.220 ;
        RECT 183.745 -122.720 183.975 -121.220 ;
        RECT 184.830 -122.725 185.060 -122.225 ;
        RECT 185.810 -122.725 186.040 -122.225 ;
        RECT 186.790 -122.725 187.020 -122.225 ;
        RECT 187.770 -122.725 188.000 -122.225 ;
        RECT 195.260 -122.230 195.490 -121.230 ;
        RECT 196.240 -122.230 196.470 -121.230 ;
        RECT 197.220 -122.230 197.450 -121.230 ;
        RECT 198.200 -122.230 198.430 -121.230 ;
        RECT 200.125 -122.875 200.355 -121.375 ;
        RECT 201.105 -122.875 201.335 -121.375 ;
        RECT 202.085 -122.875 202.315 -121.375 ;
        RECT 221.235 -122.270 221.465 -121.270 ;
        RECT 222.215 -122.270 222.445 -121.270 ;
        RECT 223.195 -122.270 223.425 -121.270 ;
        RECT 224.175 -122.270 224.405 -121.270 ;
        RECT 203.170 -122.880 203.400 -122.380 ;
        RECT 204.150 -122.880 204.380 -122.380 ;
        RECT 205.130 -122.880 205.360 -122.380 ;
        RECT 206.110 -122.880 206.340 -122.380 ;
        RECT 226.100 -122.915 226.330 -121.415 ;
        RECT 227.080 -122.915 227.310 -121.415 ;
        RECT 228.060 -122.915 228.290 -121.415 ;
        RECT 229.145 -122.920 229.375 -122.420 ;
        RECT 230.125 -122.920 230.355 -122.420 ;
        RECT 231.105 -122.920 231.335 -122.420 ;
        RECT 232.085 -122.920 232.315 -122.420 ;
        RECT 239.575 -122.425 239.805 -121.425 ;
        RECT 240.555 -122.425 240.785 -121.425 ;
        RECT 241.535 -122.425 241.765 -121.425 ;
        RECT 242.515 -122.425 242.745 -121.425 ;
        RECT 244.440 -123.070 244.670 -121.570 ;
        RECT 245.420 -123.070 245.650 -121.570 ;
        RECT 246.400 -123.070 246.630 -121.570 ;
        RECT 267.225 -122.100 267.455 -121.100 ;
        RECT 268.205 -122.100 268.435 -121.100 ;
        RECT 269.185 -122.100 269.415 -121.100 ;
        RECT 270.165 -122.100 270.395 -121.100 ;
        RECT 247.485 -123.075 247.715 -122.575 ;
        RECT 248.465 -123.075 248.695 -122.575 ;
        RECT 249.445 -123.075 249.675 -122.575 ;
        RECT 250.425 -123.075 250.655 -122.575 ;
        RECT 272.090 -122.745 272.320 -121.245 ;
        RECT 273.070 -122.745 273.300 -121.245 ;
        RECT 274.050 -122.745 274.280 -121.245 ;
        RECT 275.135 -122.750 275.365 -122.250 ;
        RECT 276.115 -122.750 276.345 -122.250 ;
        RECT 277.095 -122.750 277.325 -122.250 ;
        RECT 278.075 -122.750 278.305 -122.250 ;
        RECT 285.565 -122.255 285.795 -121.255 ;
        RECT 286.545 -122.255 286.775 -121.255 ;
        RECT 287.525 -122.255 287.755 -121.255 ;
        RECT 288.505 -122.255 288.735 -121.255 ;
        RECT 290.430 -122.900 290.660 -121.400 ;
        RECT 291.410 -122.900 291.640 -121.400 ;
        RECT 292.390 -122.900 292.620 -121.400 ;
        RECT 310.995 -121.770 311.225 -120.770 ;
        RECT 311.975 -121.770 312.205 -120.770 ;
        RECT 312.955 -121.770 313.185 -120.770 ;
        RECT 313.935 -121.770 314.165 -120.770 ;
        RECT 293.475 -122.905 293.705 -122.405 ;
        RECT 294.455 -122.905 294.685 -122.405 ;
        RECT 295.435 -122.905 295.665 -122.405 ;
        RECT 296.415 -122.905 296.645 -122.405 ;
        RECT 315.860 -122.415 316.090 -120.915 ;
        RECT 316.840 -122.415 317.070 -120.915 ;
        RECT 317.820 -122.415 318.050 -120.915 ;
        RECT 318.905 -122.420 319.135 -121.920 ;
        RECT 319.885 -122.420 320.115 -121.920 ;
        RECT 320.865 -122.420 321.095 -121.920 ;
        RECT 321.845 -122.420 322.075 -121.920 ;
        RECT 329.335 -121.925 329.565 -120.925 ;
        RECT 330.315 -121.925 330.545 -120.925 ;
        RECT 331.295 -121.925 331.525 -120.925 ;
        RECT 332.275 -121.925 332.505 -120.925 ;
        RECT 334.200 -122.570 334.430 -121.070 ;
        RECT 335.180 -122.570 335.410 -121.070 ;
        RECT 336.160 -122.570 336.390 -121.070 ;
        RECT 356.760 -121.685 356.990 -120.685 ;
        RECT 357.740 -121.685 357.970 -120.685 ;
        RECT 358.720 -121.685 358.950 -120.685 ;
        RECT 359.700 -121.685 359.930 -120.685 ;
        RECT 337.245 -122.575 337.475 -122.075 ;
        RECT 338.225 -122.575 338.455 -122.075 ;
        RECT 339.205 -122.575 339.435 -122.075 ;
        RECT 340.185 -122.575 340.415 -122.075 ;
        RECT 361.625 -122.330 361.855 -120.830 ;
        RECT 362.605 -122.330 362.835 -120.830 ;
        RECT 363.585 -122.330 363.815 -120.830 ;
        RECT 364.670 -122.335 364.900 -121.835 ;
        RECT 365.650 -122.335 365.880 -121.835 ;
        RECT 366.630 -122.335 366.860 -121.835 ;
        RECT 367.610 -122.335 367.840 -121.835 ;
        RECT 375.100 -121.840 375.330 -120.840 ;
        RECT 376.080 -121.840 376.310 -120.840 ;
        RECT 377.060 -121.840 377.290 -120.840 ;
        RECT 378.040 -121.840 378.270 -120.840 ;
        RECT 379.965 -122.485 380.195 -120.985 ;
        RECT 380.945 -122.485 381.175 -120.985 ;
        RECT 381.925 -122.485 382.155 -120.985 ;
        RECT 403.580 -121.495 403.810 -120.495 ;
        RECT 404.560 -121.495 404.790 -120.495 ;
        RECT 405.540 -121.495 405.770 -120.495 ;
        RECT 406.520 -121.495 406.750 -120.495 ;
        RECT 383.010 -122.490 383.240 -121.990 ;
        RECT 383.990 -122.490 384.220 -121.990 ;
        RECT 384.970 -122.490 385.200 -121.990 ;
        RECT 385.950 -122.490 386.180 -121.990 ;
        RECT 408.445 -122.140 408.675 -120.640 ;
        RECT 409.425 -122.140 409.655 -120.640 ;
        RECT 410.405 -122.140 410.635 -120.640 ;
        RECT 411.490 -122.145 411.720 -121.645 ;
        RECT 412.470 -122.145 412.700 -121.645 ;
        RECT 413.450 -122.145 413.680 -121.645 ;
        RECT 414.430 -122.145 414.660 -121.645 ;
        RECT 421.920 -121.650 422.150 -120.650 ;
        RECT 422.900 -121.650 423.130 -120.650 ;
        RECT 423.880 -121.650 424.110 -120.650 ;
        RECT 424.860 -121.650 425.090 -120.650 ;
        RECT 426.785 -122.295 427.015 -120.795 ;
        RECT 427.765 -122.295 427.995 -120.795 ;
        RECT 428.745 -122.295 428.975 -120.795 ;
        RECT 429.830 -122.300 430.060 -121.800 ;
        RECT 430.810 -122.300 431.040 -121.800 ;
        RECT 431.790 -122.300 432.020 -121.800 ;
        RECT 432.770 -122.300 433.000 -121.800 ;
        RECT 316.870 -123.790 317.785 -123.585 ;
        RECT 323.385 -123.790 323.865 -123.645 ;
        RECT 362.635 -123.705 363.550 -123.500 ;
        RECT 409.455 -123.515 410.370 -123.310 ;
        RECT 415.970 -123.515 416.450 -123.370 ;
        RECT 369.150 -123.705 369.630 -123.560 ;
        RECT 140.595 -124.040 141.510 -123.835 ;
        RECT 147.110 -124.040 147.590 -123.895 ;
        RECT 140.595 -124.450 147.590 -124.040 ;
        RECT 19.240 -125.505 19.470 -124.505 ;
        RECT 20.220 -125.505 20.450 -124.505 ;
        RECT 22.930 -125.505 23.160 -124.505 ;
        RECT 23.910 -125.505 24.140 -124.505 ;
        RECT 24.890 -125.505 25.120 -124.505 ;
        RECT 25.870 -125.505 26.100 -124.505 ;
        RECT 31.675 -125.450 31.905 -124.450 ;
        RECT 32.655 -125.450 32.885 -124.450 ;
        RECT 33.635 -125.450 33.865 -124.450 ;
        RECT 34.205 -125.450 34.435 -124.450 ;
        RECT 35.185 -125.450 35.415 -124.450 ;
        RECT 35.750 -125.450 35.980 -124.450 ;
        RECT 36.730 -125.450 36.960 -124.450 ;
        RECT 140.595 -124.485 141.510 -124.450 ;
        RECT 147.110 -124.580 147.590 -124.450 ;
        RECT 164.210 -124.150 164.665 -124.090 ;
        RECT 165.460 -124.150 166.215 -124.015 ;
        RECT 164.210 -124.845 166.215 -124.150 ;
        RECT 182.795 -124.095 183.710 -123.890 ;
        RECT 189.310 -124.095 189.790 -123.950 ;
        RECT 182.795 -124.505 189.790 -124.095 ;
        RECT 182.795 -124.540 183.710 -124.505 ;
        RECT 189.310 -124.635 189.790 -124.505 ;
        RECT 206.410 -124.205 206.865 -124.145 ;
        RECT 207.660 -124.205 208.415 -124.070 ;
        RECT 164.210 -124.905 164.665 -124.845 ;
        RECT 165.460 -124.970 166.215 -124.845 ;
        RECT 206.410 -124.900 208.415 -124.205 ;
        RECT 227.110 -124.290 228.025 -124.085 ;
        RECT 273.100 -124.120 274.015 -123.915 ;
        RECT 279.615 -124.120 280.095 -123.975 ;
        RECT 233.625 -124.290 234.105 -124.145 ;
        RECT 227.110 -124.700 234.105 -124.290 ;
        RECT 227.110 -124.735 228.025 -124.700 ;
        RECT 233.625 -124.830 234.105 -124.700 ;
        RECT 250.725 -124.400 251.180 -124.340 ;
        RECT 251.975 -124.400 252.730 -124.265 ;
        RECT 206.410 -124.960 206.865 -124.900 ;
        RECT 207.660 -125.025 208.415 -124.900 ;
        RECT 250.725 -125.095 252.730 -124.400 ;
        RECT 273.100 -124.530 280.095 -124.120 ;
        RECT 273.100 -124.565 274.015 -124.530 ;
        RECT 279.615 -124.660 280.095 -124.530 ;
        RECT 296.715 -124.230 297.170 -124.170 ;
        RECT 297.965 -124.230 298.720 -124.095 ;
        RECT 296.715 -124.925 298.720 -124.230 ;
        RECT 316.870 -124.200 323.865 -123.790 ;
        RECT 316.870 -124.235 317.785 -124.200 ;
        RECT 323.385 -124.330 323.865 -124.200 ;
        RECT 340.485 -123.900 340.940 -123.840 ;
        RECT 341.735 -123.900 342.490 -123.765 ;
        RECT 340.485 -124.595 342.490 -123.900 ;
        RECT 362.635 -124.115 369.630 -123.705 ;
        RECT 362.635 -124.150 363.550 -124.115 ;
        RECT 369.150 -124.245 369.630 -124.115 ;
        RECT 386.250 -123.815 386.705 -123.755 ;
        RECT 387.500 -123.815 388.255 -123.680 ;
        RECT 386.250 -124.510 388.255 -123.815 ;
        RECT 409.455 -123.925 416.450 -123.515 ;
        RECT 409.455 -123.960 410.370 -123.925 ;
        RECT 415.970 -124.055 416.450 -123.925 ;
        RECT 433.070 -123.625 433.525 -123.565 ;
        RECT 434.320 -123.625 435.075 -123.490 ;
        RECT 433.070 -124.320 435.075 -123.625 ;
        RECT 433.070 -124.380 433.525 -124.320 ;
        RECT 434.320 -124.445 435.075 -124.320 ;
        RECT 386.250 -124.570 386.705 -124.510 ;
        RECT 340.485 -124.655 340.940 -124.595 ;
        RECT 341.735 -124.720 342.490 -124.595 ;
        RECT 387.500 -124.635 388.255 -124.510 ;
        RECT 296.715 -124.985 297.170 -124.925 ;
        RECT 297.965 -125.050 298.720 -124.925 ;
        RECT 250.725 -125.155 251.180 -125.095 ;
        RECT 251.975 -125.220 252.730 -125.095 ;
        RECT -7.610 -125.795 -6.995 -125.750 ;
        RECT -6.140 -125.795 -5.525 -125.755 ;
        RECT -7.610 -126.370 -5.525 -125.795 ;
        RECT 8.750 -125.760 9.365 -125.690 ;
        RECT 10.695 -125.760 11.310 -125.695 ;
        RECT 8.750 -126.295 11.310 -125.760 ;
        RECT 8.750 -126.370 9.365 -126.295 ;
        RECT -7.610 -126.430 -6.995 -126.370 ;
        RECT -6.140 -126.435 -5.525 -126.370 ;
        RECT 10.695 -126.375 11.310 -126.295 ;
        RECT 16.835 -125.910 17.450 -125.810 ;
        RECT 18.840 -125.910 19.455 -125.820 ;
        RECT 16.835 -126.445 19.455 -125.910 ;
        RECT 16.835 -126.490 17.450 -126.445 ;
        RECT 18.840 -126.500 19.455 -126.445 ;
        RECT 25.620 -125.885 26.235 -125.795 ;
        RECT 31.700 -125.885 32.315 -125.790 ;
        RECT 25.620 -126.410 32.315 -125.885 ;
        RECT 25.620 -126.475 26.235 -126.410 ;
        RECT 31.700 -126.470 32.315 -126.410 ;
        RECT 134.590 -127.165 134.820 -125.665 ;
        RECT 135.570 -127.165 135.800 -125.665 ;
        RECT 136.550 -127.165 136.780 -125.665 ;
        RECT 137.635 -126.160 137.865 -125.660 ;
        RECT 138.615 -126.160 138.845 -125.660 ;
        RECT 139.595 -126.160 139.825 -125.660 ;
        RECT 140.575 -126.160 140.805 -125.660 ;
        RECT 141.825 -128.220 142.055 -125.220 ;
        RECT 142.805 -128.220 143.035 -125.220 ;
        RECT 144.920 -128.220 145.150 -125.220 ;
        RECT 152.930 -127.320 153.160 -125.820 ;
        RECT 153.910 -127.320 154.140 -125.820 ;
        RECT 154.890 -127.320 155.120 -125.820 ;
        RECT 155.975 -126.315 156.205 -125.815 ;
        RECT 156.955 -126.315 157.185 -125.815 ;
        RECT 157.935 -126.315 158.165 -125.815 ;
        RECT 158.915 -126.315 159.145 -125.815 ;
        RECT -97.720 -129.825 -96.760 -128.965 ;
        RECT -26.740 -129.760 -26.125 -129.080 ;
        RECT 52.830 -129.300 53.060 -128.300 ;
        RECT 53.810 -129.300 54.040 -128.300 ;
        RECT 54.790 -129.300 55.020 -128.300 ;
        RECT 57.240 -129.300 57.470 -128.300 ;
        RECT 58.220 -129.300 58.450 -128.300 ;
        RECT 59.200 -129.300 59.430 -128.300 ;
        RECT 65.955 -129.300 66.185 -128.300 ;
        RECT 66.935 -129.300 67.165 -128.300 ;
        RECT 67.915 -129.300 68.145 -128.300 ;
        RECT 70.740 -129.300 70.970 -128.300 ;
        RECT 71.720 -129.300 71.950 -128.300 ;
        RECT 72.700 -129.300 72.930 -128.300 ;
        RECT 79.455 -129.300 79.685 -128.300 ;
        RECT 80.435 -129.300 80.665 -128.300 ;
        RECT 81.415 -129.300 81.645 -128.300 ;
        RECT 160.165 -128.375 160.395 -125.375 ;
        RECT 161.145 -128.375 161.375 -125.375 ;
        RECT 163.260 -128.375 163.490 -125.375 ;
        RECT 176.790 -127.220 177.020 -125.720 ;
        RECT 177.770 -127.220 178.000 -125.720 ;
        RECT 178.750 -127.220 178.980 -125.720 ;
        RECT 179.835 -126.215 180.065 -125.715 ;
        RECT 180.815 -126.215 181.045 -125.715 ;
        RECT 181.795 -126.215 182.025 -125.715 ;
        RECT 182.775 -126.215 183.005 -125.715 ;
        RECT 184.025 -128.275 184.255 -125.275 ;
        RECT 185.005 -128.275 185.235 -125.275 ;
        RECT 187.120 -128.275 187.350 -125.275 ;
        RECT 195.130 -127.375 195.360 -125.875 ;
        RECT 196.110 -127.375 196.340 -125.875 ;
        RECT 197.090 -127.375 197.320 -125.875 ;
        RECT 198.175 -126.370 198.405 -125.870 ;
        RECT 199.155 -126.370 199.385 -125.870 ;
        RECT 200.135 -126.370 200.365 -125.870 ;
        RECT 201.115 -126.370 201.345 -125.870 ;
        RECT 202.365 -128.430 202.595 -125.430 ;
        RECT 203.345 -128.430 203.575 -125.430 ;
        RECT 205.460 -128.430 205.690 -125.430 ;
        RECT 221.105 -127.415 221.335 -125.915 ;
        RECT 222.085 -127.415 222.315 -125.915 ;
        RECT 223.065 -127.415 223.295 -125.915 ;
        RECT 224.150 -126.410 224.380 -125.910 ;
        RECT 225.130 -126.410 225.360 -125.910 ;
        RECT 226.110 -126.410 226.340 -125.910 ;
        RECT 227.090 -126.410 227.320 -125.910 ;
        RECT 228.340 -128.470 228.570 -125.470 ;
        RECT 229.320 -128.470 229.550 -125.470 ;
        RECT 231.435 -128.470 231.665 -125.470 ;
        RECT 239.445 -127.570 239.675 -126.070 ;
        RECT 240.425 -127.570 240.655 -126.070 ;
        RECT 241.405 -127.570 241.635 -126.070 ;
        RECT 242.490 -126.565 242.720 -126.065 ;
        RECT 243.470 -126.565 243.700 -126.065 ;
        RECT 244.450 -126.565 244.680 -126.065 ;
        RECT 245.430 -126.565 245.660 -126.065 ;
        RECT 246.680 -128.625 246.910 -125.625 ;
        RECT 247.660 -128.625 247.890 -125.625 ;
        RECT 249.775 -128.625 250.005 -125.625 ;
        RECT 267.095 -127.245 267.325 -125.745 ;
        RECT 268.075 -127.245 268.305 -125.745 ;
        RECT 269.055 -127.245 269.285 -125.745 ;
        RECT 270.140 -126.240 270.370 -125.740 ;
        RECT 271.120 -126.240 271.350 -125.740 ;
        RECT 272.100 -126.240 272.330 -125.740 ;
        RECT 273.080 -126.240 273.310 -125.740 ;
        RECT 274.330 -128.300 274.560 -125.300 ;
        RECT 275.310 -128.300 275.540 -125.300 ;
        RECT 277.425 -128.300 277.655 -125.300 ;
        RECT 285.435 -127.400 285.665 -125.900 ;
        RECT 286.415 -127.400 286.645 -125.900 ;
        RECT 287.395 -127.400 287.625 -125.900 ;
        RECT 288.480 -126.395 288.710 -125.895 ;
        RECT 289.460 -126.395 289.690 -125.895 ;
        RECT 290.440 -126.395 290.670 -125.895 ;
        RECT 291.420 -126.395 291.650 -125.895 ;
        RECT 292.670 -128.455 292.900 -125.455 ;
        RECT 293.650 -128.455 293.880 -125.455 ;
        RECT 295.765 -128.455 295.995 -125.455 ;
        RECT 310.865 -126.915 311.095 -125.415 ;
        RECT 311.845 -126.915 312.075 -125.415 ;
        RECT 312.825 -126.915 313.055 -125.415 ;
        RECT 313.910 -125.910 314.140 -125.410 ;
        RECT 314.890 -125.910 315.120 -125.410 ;
        RECT 315.870 -125.910 316.100 -125.410 ;
        RECT 316.850 -125.910 317.080 -125.410 ;
        RECT 318.100 -127.970 318.330 -124.970 ;
        RECT 319.080 -127.970 319.310 -124.970 ;
        RECT 321.195 -127.970 321.425 -124.970 ;
        RECT 329.205 -127.070 329.435 -125.570 ;
        RECT 330.185 -127.070 330.415 -125.570 ;
        RECT 331.165 -127.070 331.395 -125.570 ;
        RECT 332.250 -126.065 332.480 -125.565 ;
        RECT 333.230 -126.065 333.460 -125.565 ;
        RECT 334.210 -126.065 334.440 -125.565 ;
        RECT 335.190 -126.065 335.420 -125.565 ;
        RECT 336.440 -128.125 336.670 -125.125 ;
        RECT 337.420 -128.125 337.650 -125.125 ;
        RECT 339.535 -128.125 339.765 -125.125 ;
        RECT 356.630 -126.830 356.860 -125.330 ;
        RECT 357.610 -126.830 357.840 -125.330 ;
        RECT 358.590 -126.830 358.820 -125.330 ;
        RECT 359.675 -125.825 359.905 -125.325 ;
        RECT 360.655 -125.825 360.885 -125.325 ;
        RECT 361.635 -125.825 361.865 -125.325 ;
        RECT 362.615 -125.825 362.845 -125.325 ;
        RECT 363.865 -127.885 364.095 -124.885 ;
        RECT 364.845 -127.885 365.075 -124.885 ;
        RECT 366.960 -127.885 367.190 -124.885 ;
        RECT 374.970 -126.985 375.200 -125.485 ;
        RECT 375.950 -126.985 376.180 -125.485 ;
        RECT 376.930 -126.985 377.160 -125.485 ;
        RECT 378.015 -125.980 378.245 -125.480 ;
        RECT 378.995 -125.980 379.225 -125.480 ;
        RECT 379.975 -125.980 380.205 -125.480 ;
        RECT 380.955 -125.980 381.185 -125.480 ;
        RECT 382.205 -128.040 382.435 -125.040 ;
        RECT 383.185 -128.040 383.415 -125.040 ;
        RECT 385.300 -128.040 385.530 -125.040 ;
        RECT 403.450 -126.640 403.680 -125.140 ;
        RECT 404.430 -126.640 404.660 -125.140 ;
        RECT 405.410 -126.640 405.640 -125.140 ;
        RECT 406.495 -125.635 406.725 -125.135 ;
        RECT 407.475 -125.635 407.705 -125.135 ;
        RECT 408.455 -125.635 408.685 -125.135 ;
        RECT 409.435 -125.635 409.665 -125.135 ;
        RECT 410.685 -127.695 410.915 -124.695 ;
        RECT 411.665 -127.695 411.895 -124.695 ;
        RECT 413.780 -127.695 414.010 -124.695 ;
        RECT 421.790 -126.795 422.020 -125.295 ;
        RECT 422.770 -126.795 423.000 -125.295 ;
        RECT 423.750 -126.795 423.980 -125.295 ;
        RECT 424.835 -125.790 425.065 -125.290 ;
        RECT 425.815 -125.790 426.045 -125.290 ;
        RECT 426.795 -125.790 427.025 -125.290 ;
        RECT 427.775 -125.790 428.005 -125.290 ;
        RECT 429.025 -127.850 429.255 -124.850 ;
        RECT 430.005 -127.850 430.235 -124.850 ;
        RECT 432.120 -127.850 432.350 -124.850 ;
        RECT -95.415 -132.485 -95.185 -131.485 ;
        RECT -94.435 -132.485 -94.205 -131.485 ;
        RECT -93.455 -132.485 -93.225 -131.485 ;
        RECT -92.475 -132.485 -92.245 -131.485 ;
        RECT -90.550 -132.340 -90.320 -130.840 ;
        RECT -89.570 -132.340 -89.340 -130.840 ;
        RECT -88.590 -132.340 -88.360 -130.840 ;
        RECT -87.505 -131.335 -87.275 -130.835 ;
        RECT -86.525 -131.335 -86.295 -130.835 ;
        RECT -85.545 -131.335 -85.315 -130.835 ;
        RECT -84.565 -131.335 -84.335 -130.835 ;
        RECT -26.715 -132.915 -26.145 -129.760 ;
        RECT -13.905 -130.480 -13.290 -129.800 ;
        RECT -13.880 -132.740 -13.310 -130.480 ;
        RECT -1.490 -130.650 0.040 -130.340 ;
        RECT -1.490 -130.655 -0.875 -130.650 ;
        RECT -1.465 -132.740 -0.895 -130.655 ;
        RECT -26.735 -133.595 -26.120 -132.915 ;
        RECT -13.900 -133.420 -13.285 -132.740 ;
        RECT -1.485 -133.420 -0.870 -132.740 ;
        RECT -114.795 -137.135 -114.565 -136.135 ;
        RECT -113.815 -137.135 -113.585 -136.135 ;
        RECT -111.105 -137.135 -110.875 -136.135 ;
        RECT -110.125 -137.135 -109.895 -136.135 ;
        RECT -109.145 -137.135 -108.915 -136.135 ;
        RECT -108.165 -137.135 -107.935 -136.135 ;
        RECT -101.745 -137.955 -100.865 -134.800 ;
        RECT -33.375 -136.705 -33.145 -135.705 ;
        RECT -32.395 -136.705 -32.165 -135.705 ;
        RECT -31.415 -136.705 -31.185 -135.705 ;
        RECT -30.845 -136.705 -30.615 -135.705 ;
        RECT -29.865 -136.705 -29.635 -135.705 ;
        RECT -29.300 -136.705 -29.070 -135.705 ;
        RECT -28.320 -136.705 -28.090 -135.705 ;
        RECT -20.875 -136.705 -20.645 -135.705 ;
        RECT -19.895 -136.705 -19.665 -135.705 ;
        RECT -18.915 -136.705 -18.685 -135.705 ;
        RECT -18.345 -136.705 -18.115 -135.705 ;
        RECT -17.365 -136.705 -17.135 -135.705 ;
        RECT -16.800 -136.705 -16.570 -135.705 ;
        RECT -15.820 -136.705 -15.590 -135.705 ;
        RECT -8.375 -136.705 -8.145 -135.705 ;
        RECT -7.395 -136.705 -7.165 -135.705 ;
        RECT -6.415 -136.705 -6.185 -135.705 ;
        RECT -5.845 -136.705 -5.615 -135.705 ;
        RECT -4.865 -136.705 -4.635 -135.705 ;
        RECT -4.300 -136.705 -4.070 -135.705 ;
        RECT -3.320 -136.705 -3.090 -135.705 ;
        RECT 4.125 -136.705 4.355 -135.705 ;
        RECT 5.105 -136.705 5.335 -135.705 ;
        RECT 6.085 -136.705 6.315 -135.705 ;
        RECT 6.655 -136.705 6.885 -135.705 ;
        RECT 7.635 -136.705 7.865 -135.705 ;
        RECT 8.200 -136.705 8.430 -135.705 ;
        RECT 9.180 -136.705 9.410 -135.705 ;
        RECT 16.625 -136.705 16.855 -135.705 ;
        RECT 17.605 -136.705 17.835 -135.705 ;
        RECT 18.585 -136.705 18.815 -135.705 ;
        RECT 19.155 -136.705 19.385 -135.705 ;
        RECT 20.135 -136.705 20.365 -135.705 ;
        RECT 20.700 -136.705 20.930 -135.705 ;
        RECT 21.680 -136.705 21.910 -135.705 ;
        RECT 31.625 -136.705 31.855 -135.705 ;
        RECT 32.605 -136.705 32.835 -135.705 ;
        RECT 33.585 -136.705 33.815 -135.705 ;
        RECT 34.155 -136.705 34.385 -135.705 ;
        RECT 35.135 -136.705 35.365 -135.705 ;
        RECT 35.700 -136.705 35.930 -135.705 ;
        RECT 36.680 -136.705 36.910 -135.705 ;
        RECT 62.260 -135.890 62.490 -134.890 ;
        RECT 63.240 -135.890 63.470 -134.890 ;
        RECT 64.220 -135.890 64.450 -134.890 ;
        RECT 66.445 -135.890 66.675 -134.890 ;
        RECT 67.425 -135.890 67.655 -134.890 ;
        RECT 68.405 -135.890 68.635 -134.890 ;
        RECT 75.760 -135.890 75.990 -134.890 ;
        RECT 76.740 -135.890 76.970 -134.890 ;
        RECT 77.720 -135.890 77.950 -134.890 ;
        RECT 79.945 -135.890 80.175 -134.890 ;
        RECT 80.925 -135.890 81.155 -134.890 ;
        RECT 81.905 -135.890 82.135 -134.890 ;
        RECT -130.060 -170.885 -128.060 -170.655 ;
        RECT -130.060 -172.065 -128.060 -171.835 ;
        RECT -130.060 -173.245 -128.060 -173.015 ;
        RECT -130.060 -174.425 -128.060 -174.195 ;
        RECT -130.060 -175.605 -128.060 -175.375 ;
        RECT -72.235 -175.940 -72.005 -174.940 ;
        RECT -71.255 -175.940 -71.025 -174.940 ;
        RECT -70.275 -175.940 -70.045 -174.940 ;
        RECT -68.050 -175.940 -67.820 -174.940 ;
        RECT -67.070 -175.940 -66.840 -174.940 ;
        RECT -66.090 -175.940 -65.860 -174.940 ;
        RECT -58.735 -175.940 -58.505 -174.940 ;
        RECT -57.755 -175.940 -57.525 -174.940 ;
        RECT -56.775 -175.940 -56.545 -174.940 ;
        RECT -54.550 -175.940 -54.320 -174.940 ;
        RECT -53.570 -175.940 -53.340 -174.940 ;
        RECT -52.590 -175.940 -52.360 -174.940 ;
        RECT -130.060 -176.785 -128.060 -176.555 ;
        RECT -130.060 -177.965 -128.060 -177.735 ;
        RECT -40.425 -177.990 -40.195 -174.990 ;
        RECT -38.310 -177.990 -38.080 -174.990 ;
        RECT -37.330 -177.990 -37.100 -174.990 ;
        RECT -29.885 -176.970 -29.655 -175.970 ;
        RECT -28.905 -176.970 -28.675 -175.970 ;
        RECT -27.925 -176.970 -27.695 -175.970 ;
        RECT -27.355 -176.970 -27.125 -175.970 ;
        RECT -26.375 -176.970 -26.145 -175.970 ;
        RECT -25.810 -176.970 -25.580 -175.970 ;
        RECT -24.830 -176.970 -24.600 -175.970 ;
        RECT -17.385 -176.970 -17.155 -175.970 ;
        RECT -16.405 -176.970 -16.175 -175.970 ;
        RECT -15.425 -176.970 -15.195 -175.970 ;
        RECT -14.855 -176.970 -14.625 -175.970 ;
        RECT -13.875 -176.970 -13.645 -175.970 ;
        RECT -13.310 -176.970 -13.080 -175.970 ;
        RECT -12.330 -176.970 -12.100 -175.970 ;
        RECT -4.885 -176.970 -4.655 -175.970 ;
        RECT -3.905 -176.970 -3.675 -175.970 ;
        RECT -2.925 -176.970 -2.695 -175.970 ;
        RECT -2.355 -176.970 -2.125 -175.970 ;
        RECT -1.375 -176.970 -1.145 -175.970 ;
        RECT -0.810 -176.970 -0.580 -175.970 ;
        RECT 0.170 -176.970 0.400 -175.970 ;
        RECT 7.615 -176.970 7.845 -175.970 ;
        RECT 8.595 -176.970 8.825 -175.970 ;
        RECT 9.575 -176.970 9.805 -175.970 ;
        RECT 10.145 -176.970 10.375 -175.970 ;
        RECT 11.125 -176.970 11.355 -175.970 ;
        RECT 11.690 -176.970 11.920 -175.970 ;
        RECT 12.670 -176.970 12.900 -175.970 ;
        RECT 20.115 -176.970 20.345 -175.970 ;
        RECT 21.095 -176.970 21.325 -175.970 ;
        RECT 22.075 -176.970 22.305 -175.970 ;
        RECT 22.645 -176.970 22.875 -175.970 ;
        RECT 23.625 -176.970 23.855 -175.970 ;
        RECT 24.190 -176.970 24.420 -175.970 ;
        RECT 25.170 -176.970 25.400 -175.970 ;
        RECT 35.115 -176.970 35.345 -175.970 ;
        RECT 36.095 -176.970 36.325 -175.970 ;
        RECT 37.075 -176.970 37.305 -175.970 ;
        RECT 37.645 -176.970 37.875 -175.970 ;
        RECT 38.625 -176.970 38.855 -175.970 ;
        RECT 39.190 -176.970 39.420 -175.970 ;
        RECT 40.170 -176.970 40.400 -175.970 ;
        RECT -130.060 -179.145 -128.060 -178.915 ;
        RECT -110.230 -179.875 -110.000 -178.875 ;
        RECT -109.250 -179.875 -109.020 -178.875 ;
        RECT -108.270 -179.875 -108.040 -178.875 ;
        RECT -107.290 -179.875 -107.060 -178.875 ;
        RECT -104.580 -179.875 -104.350 -178.875 ;
        RECT -103.600 -179.875 -103.370 -178.875 ;
        RECT -130.060 -180.325 -128.060 -180.095 ;
        RECT -100.235 -180.985 -100.005 -179.485 ;
        RECT -99.255 -180.985 -99.025 -179.485 ;
        RECT -98.275 -180.985 -98.045 -179.485 ;
        RECT -97.190 -179.980 -96.960 -179.480 ;
        RECT -96.210 -179.980 -95.980 -179.480 ;
        RECT -95.230 -179.980 -95.000 -179.480 ;
        RECT -94.250 -179.980 -94.020 -179.480 ;
        RECT -23.245 -179.760 -22.630 -179.080 ;
        RECT -130.060 -181.505 -128.060 -181.275 ;
        RECT -130.060 -182.685 -128.060 -182.455 ;
        RECT -71.745 -182.530 -71.515 -181.530 ;
        RECT -70.765 -182.530 -70.535 -181.530 ;
        RECT -69.785 -182.530 -69.555 -181.530 ;
        RECT -63.030 -182.530 -62.800 -181.530 ;
        RECT -62.050 -182.530 -61.820 -181.530 ;
        RECT -61.070 -182.530 -60.840 -181.530 ;
        RECT -58.245 -182.530 -58.015 -181.530 ;
        RECT -57.265 -182.530 -57.035 -181.530 ;
        RECT -56.285 -182.530 -56.055 -181.530 ;
        RECT -49.530 -182.530 -49.300 -181.530 ;
        RECT -48.550 -182.530 -48.320 -181.530 ;
        RECT -47.570 -182.530 -47.340 -181.530 ;
        RECT -45.120 -182.530 -44.890 -181.530 ;
        RECT -44.140 -182.530 -43.910 -181.530 ;
        RECT -43.160 -182.530 -42.930 -181.530 ;
        RECT -130.060 -183.865 -128.060 -183.635 ;
        RECT -130.060 -185.045 -128.060 -184.815 ;
        RECT -92.055 -185.795 -91.825 -184.295 ;
        RECT -91.075 -185.795 -90.845 -184.295 ;
        RECT -90.095 -185.795 -89.865 -184.295 ;
        RECT -89.010 -185.800 -88.780 -185.300 ;
        RECT -88.030 -185.800 -87.800 -185.300 ;
        RECT -87.050 -185.800 -86.820 -185.300 ;
        RECT -86.070 -185.800 -85.840 -185.300 ;
        RECT -130.060 -186.225 -128.060 -185.995 ;
        RECT -84.820 -186.240 -84.590 -183.240 ;
        RECT -83.840 -186.240 -83.610 -183.240 ;
        RECT -81.725 -186.240 -81.495 -183.240 ;
        RECT -31.580 -183.615 -31.350 -182.615 ;
        RECT -30.600 -183.615 -30.370 -182.615 ;
        RECT -29.620 -183.615 -29.390 -182.615 ;
        RECT -23.225 -182.915 -22.655 -179.760 ;
        RECT -10.410 -179.935 -9.795 -179.255 ;
        RECT 2.005 -179.935 2.620 -179.255 ;
        RECT -10.390 -182.195 -9.820 -179.935 ;
        RECT 2.025 -182.020 2.595 -179.935 ;
        RECT 2.000 -182.025 2.615 -182.020 ;
        RECT -10.415 -182.875 -9.800 -182.195 ;
        RECT 2.000 -182.335 3.530 -182.025 ;
        RECT -23.250 -183.595 -22.635 -182.915 ;
        RECT 20.325 -186.230 20.940 -186.185 ;
        RECT 22.330 -186.230 22.945 -186.175 ;
        RECT -4.120 -186.305 -3.505 -186.245 ;
        RECT -2.650 -186.305 -2.035 -186.240 ;
        RECT -4.120 -186.880 -2.035 -186.305 ;
        RECT -4.120 -186.925 -3.505 -186.880 ;
        RECT -2.650 -186.920 -2.035 -186.880 ;
        RECT 12.240 -186.380 12.855 -186.305 ;
        RECT 14.185 -186.380 14.800 -186.300 ;
        RECT 12.240 -186.915 14.800 -186.380 ;
        RECT 20.325 -186.765 22.945 -186.230 ;
        RECT 20.325 -186.865 20.940 -186.765 ;
        RECT 22.330 -186.855 22.945 -186.765 ;
        RECT 29.110 -186.265 29.725 -186.200 ;
        RECT 35.190 -186.265 35.805 -186.205 ;
        RECT 29.110 -186.790 35.805 -186.265 ;
        RECT 29.110 -186.880 29.725 -186.790 ;
        RECT 35.190 -186.885 35.805 -186.790 ;
        RECT 12.240 -186.985 12.855 -186.915 ;
        RECT 14.185 -186.980 14.800 -186.915 ;
        RECT -130.060 -187.405 -128.060 -187.175 ;
        RECT -130.060 -188.585 -128.060 -188.355 ;
        RECT -130.060 -189.825 -128.060 -189.595 ;
        RECT -109.945 -190.530 -109.715 -189.030 ;
        RECT -108.965 -190.530 -108.735 -189.030 ;
        RECT -107.985 -190.530 -107.755 -189.030 ;
        RECT -106.900 -189.525 -106.670 -189.025 ;
        RECT -105.920 -189.525 -105.690 -189.025 ;
        RECT -104.940 -189.525 -104.710 -189.025 ;
        RECT -103.960 -189.525 -103.730 -189.025 ;
        RECT -101.080 -189.555 -100.850 -188.555 ;
        RECT -100.100 -189.555 -99.870 -188.555 ;
        RECT -99.120 -189.555 -98.890 -188.555 ;
        RECT -98.140 -189.555 -97.910 -188.555 ;
        RECT -95.430 -189.555 -95.200 -188.555 ;
        RECT -94.450 -189.555 -94.220 -188.555 ;
        RECT -91.925 -190.440 -91.695 -189.440 ;
        RECT -90.945 -190.440 -90.715 -189.440 ;
        RECT -89.965 -190.440 -89.735 -189.440 ;
        RECT -88.985 -190.440 -88.755 -189.440 ;
        RECT -87.060 -190.295 -86.830 -188.795 ;
        RECT -86.080 -190.295 -85.850 -188.795 ;
        RECT -85.100 -190.295 -84.870 -188.795 ;
        RECT -84.015 -189.290 -83.785 -188.790 ;
        RECT -83.035 -189.290 -82.805 -188.790 ;
        RECT -82.055 -189.290 -81.825 -188.790 ;
        RECT -81.075 -189.290 -80.845 -188.790 ;
        RECT -67.110 -190.675 -66.880 -189.175 ;
        RECT -66.130 -190.675 -65.900 -189.175 ;
        RECT -65.150 -190.675 -64.920 -189.175 ;
        RECT -64.065 -190.680 -63.835 -190.180 ;
        RECT -63.085 -190.680 -62.855 -190.180 ;
        RECT -62.105 -190.680 -61.875 -190.180 ;
        RECT -61.125 -190.680 -60.895 -190.180 ;
        RECT -130.060 -191.005 -128.060 -190.775 ;
        RECT -59.875 -191.120 -59.645 -188.120 ;
        RECT -58.895 -191.120 -58.665 -188.120 ;
        RECT -56.780 -191.120 -56.550 -188.120 ;
        RECT -32.375 -188.130 -32.145 -187.130 ;
        RECT -31.395 -188.130 -31.165 -187.130 ;
        RECT -30.415 -188.130 -30.185 -187.130 ;
        RECT -23.660 -188.130 -23.430 -187.130 ;
        RECT -22.680 -188.130 -22.450 -187.130 ;
        RECT -21.700 -188.130 -21.470 -187.130 ;
        RECT -18.875 -188.130 -18.645 -187.130 ;
        RECT -17.895 -188.130 -17.665 -187.130 ;
        RECT -16.915 -188.130 -16.685 -187.130 ;
        RECT -10.160 -188.130 -9.930 -187.130 ;
        RECT -9.180 -188.130 -8.950 -187.130 ;
        RECT -8.200 -188.130 -7.970 -187.130 ;
        RECT -5.750 -188.130 -5.520 -187.130 ;
        RECT -4.770 -188.130 -4.540 -187.130 ;
        RECT -3.790 -188.130 -3.560 -187.130 ;
        RECT -2.080 -188.215 -1.850 -187.215 ;
        RECT -1.100 -188.215 -0.870 -187.215 ;
        RECT 1.610 -188.215 1.840 -187.215 ;
        RECT 2.590 -188.215 2.820 -187.215 ;
        RECT 3.570 -188.215 3.800 -187.215 ;
        RECT 4.550 -188.215 4.780 -187.215 ;
        RECT 6.585 -187.780 6.815 -187.280 ;
        RECT 7.565 -187.780 7.795 -187.280 ;
        RECT 8.545 -187.780 8.775 -187.280 ;
        RECT 9.525 -187.780 9.755 -187.280 ;
        RECT 10.610 -188.785 10.840 -187.285 ;
        RECT 11.590 -188.785 11.820 -187.285 ;
        RECT 12.570 -188.785 12.800 -187.285 ;
        RECT 14.610 -187.790 14.840 -187.290 ;
        RECT 15.590 -187.790 15.820 -187.290 ;
        RECT 16.570 -187.790 16.800 -187.290 ;
        RECT 17.550 -187.790 17.780 -187.290 ;
        RECT 18.635 -188.795 18.865 -187.295 ;
        RECT 19.615 -188.795 19.845 -187.295 ;
        RECT 20.595 -188.795 20.825 -187.295 ;
        RECT 22.730 -188.170 22.960 -187.170 ;
        RECT 23.710 -188.170 23.940 -187.170 ;
        RECT 26.420 -188.170 26.650 -187.170 ;
        RECT 27.400 -188.170 27.630 -187.170 ;
        RECT 28.380 -188.170 28.610 -187.170 ;
        RECT 29.360 -188.170 29.590 -187.170 ;
        RECT 35.165 -188.225 35.395 -187.225 ;
        RECT 36.145 -188.225 36.375 -187.225 ;
        RECT 37.125 -188.225 37.355 -187.225 ;
        RECT 37.695 -188.225 37.925 -187.225 ;
        RECT 38.675 -188.225 38.905 -187.225 ;
        RECT 39.240 -188.225 39.470 -187.225 ;
        RECT 40.220 -188.225 40.450 -187.225 ;
        RECT 138.250 -187.710 138.480 -186.710 ;
        RECT 139.230 -187.710 139.460 -186.710 ;
        RECT 140.210 -187.710 140.440 -186.710 ;
        RECT 141.190 -187.710 141.420 -186.710 ;
        RECT 143.115 -188.355 143.345 -186.855 ;
        RECT 144.095 -188.355 144.325 -186.855 ;
        RECT 145.075 -188.355 145.305 -186.855 ;
        RECT 180.450 -187.765 180.680 -186.765 ;
        RECT 181.430 -187.765 181.660 -186.765 ;
        RECT 182.410 -187.765 182.640 -186.765 ;
        RECT 183.390 -187.765 183.620 -186.765 ;
        RECT 146.160 -188.360 146.390 -187.860 ;
        RECT 147.140 -188.360 147.370 -187.860 ;
        RECT 148.120 -188.360 148.350 -187.860 ;
        RECT 149.100 -188.360 149.330 -187.860 ;
        RECT 185.315 -188.410 185.545 -186.910 ;
        RECT 186.295 -188.410 186.525 -186.910 ;
        RECT 187.275 -188.410 187.505 -186.910 ;
        RECT 188.360 -188.415 188.590 -187.915 ;
        RECT 189.340 -188.415 189.570 -187.915 ;
        RECT 190.320 -188.415 190.550 -187.915 ;
        RECT 191.300 -188.415 191.530 -187.915 ;
        RECT 224.765 -187.960 224.995 -186.960 ;
        RECT 225.745 -187.960 225.975 -186.960 ;
        RECT 226.725 -187.960 226.955 -186.960 ;
        RECT 227.705 -187.960 227.935 -186.960 ;
        RECT 106.390 -189.475 106.620 -188.475 ;
        RECT 107.370 -189.475 107.600 -188.475 ;
        RECT 108.350 -189.475 108.580 -188.475 ;
        RECT 110.575 -189.475 110.805 -188.475 ;
        RECT 111.555 -189.475 111.785 -188.475 ;
        RECT 112.535 -189.475 112.765 -188.475 ;
        RECT 119.890 -189.475 120.120 -188.475 ;
        RECT 120.870 -189.475 121.100 -188.475 ;
        RECT 121.850 -189.475 122.080 -188.475 ;
        RECT 124.075 -189.475 124.305 -188.475 ;
        RECT 125.055 -189.475 125.285 -188.475 ;
        RECT 126.035 -189.475 126.265 -188.475 ;
        RECT 229.630 -188.605 229.860 -187.105 ;
        RECT 230.610 -188.605 230.840 -187.105 ;
        RECT 231.590 -188.605 231.820 -187.105 ;
        RECT 270.755 -187.790 270.985 -186.790 ;
        RECT 271.735 -187.790 271.965 -186.790 ;
        RECT 272.715 -187.790 272.945 -186.790 ;
        RECT 273.695 -187.790 273.925 -186.790 ;
        RECT 232.675 -188.610 232.905 -188.110 ;
        RECT 233.655 -188.610 233.885 -188.110 ;
        RECT 234.635 -188.610 234.865 -188.110 ;
        RECT 235.615 -188.610 235.845 -188.110 ;
        RECT 275.620 -188.435 275.850 -186.935 ;
        RECT 276.600 -188.435 276.830 -186.935 ;
        RECT 277.580 -188.435 277.810 -186.935 ;
        RECT 314.525 -187.460 314.755 -186.460 ;
        RECT 315.505 -187.460 315.735 -186.460 ;
        RECT 316.485 -187.460 316.715 -186.460 ;
        RECT 317.465 -187.460 317.695 -186.460 ;
        RECT 278.665 -188.440 278.895 -187.940 ;
        RECT 279.645 -188.440 279.875 -187.940 ;
        RECT 280.625 -188.440 280.855 -187.940 ;
        RECT 281.605 -188.440 281.835 -187.940 ;
        RECT 319.390 -188.105 319.620 -186.605 ;
        RECT 320.370 -188.105 320.600 -186.605 ;
        RECT 321.350 -188.105 321.580 -186.605 ;
        RECT 360.290 -187.375 360.520 -186.375 ;
        RECT 361.270 -187.375 361.500 -186.375 ;
        RECT 362.250 -187.375 362.480 -186.375 ;
        RECT 363.230 -187.375 363.460 -186.375 ;
        RECT 322.435 -188.110 322.665 -187.610 ;
        RECT 323.415 -188.110 323.645 -187.610 ;
        RECT 324.395 -188.110 324.625 -187.610 ;
        RECT 325.375 -188.110 325.605 -187.610 ;
        RECT 365.155 -188.020 365.385 -186.520 ;
        RECT 366.135 -188.020 366.365 -186.520 ;
        RECT 367.115 -188.020 367.345 -186.520 ;
        RECT 407.110 -187.185 407.340 -186.185 ;
        RECT 408.090 -187.185 408.320 -186.185 ;
        RECT 409.070 -187.185 409.300 -186.185 ;
        RECT 410.050 -187.185 410.280 -186.185 ;
        RECT 368.200 -188.025 368.430 -187.525 ;
        RECT 369.180 -188.025 369.410 -187.525 ;
        RECT 370.160 -188.025 370.390 -187.525 ;
        RECT 371.140 -188.025 371.370 -187.525 ;
        RECT 411.975 -187.830 412.205 -186.330 ;
        RECT 412.955 -187.830 413.185 -186.330 ;
        RECT 413.935 -187.830 414.165 -186.330 ;
        RECT 415.020 -187.835 415.250 -187.335 ;
        RECT 416.000 -187.835 416.230 -187.335 ;
        RECT 416.980 -187.835 417.210 -187.335 ;
        RECT 417.960 -187.835 418.190 -187.335 ;
        RECT 418.370 -189.410 418.740 -189.330 ;
        RECT 419.510 -189.410 420.060 -189.230 ;
        RECT 325.785 -189.685 326.155 -189.605 ;
        RECT 326.925 -189.685 327.475 -189.505 ;
        RECT 149.510 -189.935 149.880 -189.855 ;
        RECT 150.650 -189.935 151.200 -189.755 ;
        RECT 149.510 -190.415 151.200 -189.935 ;
        RECT 191.710 -189.990 192.080 -189.910 ;
        RECT 192.850 -189.990 193.400 -189.810 ;
        RECT 149.510 -190.445 149.880 -190.415 ;
        RECT 150.650 -190.505 151.200 -190.415 ;
        RECT -130.060 -192.185 -128.060 -191.955 ;
        RECT -130.060 -193.365 -128.060 -193.135 ;
        RECT -130.060 -194.545 -128.060 -194.315 ;
        RECT -66.980 -195.320 -66.750 -194.320 ;
        RECT -66.000 -195.320 -65.770 -194.320 ;
        RECT -65.020 -195.320 -64.790 -194.320 ;
        RECT -64.040 -195.320 -63.810 -194.320 ;
        RECT -62.115 -195.175 -61.885 -193.675 ;
        RECT -61.135 -195.175 -60.905 -193.675 ;
        RECT -60.155 -195.175 -59.925 -193.675 ;
        RECT -59.070 -194.170 -58.840 -193.670 ;
        RECT -58.090 -194.170 -57.860 -193.670 ;
        RECT -57.110 -194.170 -56.880 -193.670 ;
        RECT -56.130 -194.170 -55.900 -193.670 ;
        RECT -32.865 -194.720 -32.635 -193.720 ;
        RECT -31.885 -194.720 -31.655 -193.720 ;
        RECT -30.905 -194.720 -30.675 -193.720 ;
        RECT -28.680 -194.720 -28.450 -193.720 ;
        RECT -27.700 -194.720 -27.470 -193.720 ;
        RECT -26.720 -194.720 -26.490 -193.720 ;
        RECT -19.365 -194.720 -19.135 -193.720 ;
        RECT -18.385 -194.720 -18.155 -193.720 ;
        RECT -17.405 -194.720 -17.175 -193.720 ;
        RECT -15.180 -194.720 -14.950 -193.720 ;
        RECT -14.200 -194.720 -13.970 -193.720 ;
        RECT -13.220 -194.720 -12.990 -193.720 ;
        RECT 90.355 -195.465 90.585 -192.465 ;
        RECT 91.335 -195.465 91.565 -192.465 ;
        RECT 138.120 -192.855 138.350 -191.355 ;
        RECT 139.100 -192.855 139.330 -191.355 ;
        RECT 140.080 -192.855 140.310 -191.355 ;
        RECT 141.165 -191.850 141.395 -191.350 ;
        RECT 142.145 -191.850 142.375 -191.350 ;
        RECT 143.125 -191.850 143.355 -191.350 ;
        RECT 144.105 -191.850 144.335 -191.350 ;
        RECT 145.355 -193.910 145.585 -190.910 ;
        RECT 146.335 -193.910 146.565 -190.910 ;
        RECT 148.450 -193.910 148.680 -190.910 ;
        RECT 155.315 -192.700 155.545 -190.200 ;
        RECT 156.295 -192.700 156.525 -190.200 ;
        RECT 159.270 -192.700 159.500 -190.200 ;
        RECT 159.920 -192.700 160.150 -190.200 ;
        RECT 161.060 -191.700 161.290 -190.200 ;
        RECT 162.040 -191.700 162.270 -190.200 ;
        RECT 191.710 -190.470 193.400 -189.990 ;
        RECT 236.025 -190.185 236.395 -190.105 ;
        RECT 237.165 -190.185 237.715 -190.005 ;
        RECT 191.710 -190.500 192.080 -190.470 ;
        RECT 192.850 -190.560 193.400 -190.470 ;
        RECT 180.320 -192.910 180.550 -191.410 ;
        RECT 181.300 -192.910 181.530 -191.410 ;
        RECT 182.280 -192.910 182.510 -191.410 ;
        RECT 183.365 -191.905 183.595 -191.405 ;
        RECT 184.345 -191.905 184.575 -191.405 ;
        RECT 185.325 -191.905 185.555 -191.405 ;
        RECT 186.305 -191.905 186.535 -191.405 ;
        RECT 187.555 -193.965 187.785 -190.965 ;
        RECT 188.535 -193.965 188.765 -190.965 ;
        RECT 190.650 -193.965 190.880 -190.965 ;
        RECT 197.515 -192.755 197.745 -190.255 ;
        RECT 198.495 -192.755 198.725 -190.255 ;
        RECT 201.470 -192.755 201.700 -190.255 ;
        RECT 202.120 -192.755 202.350 -190.255 ;
        RECT 203.260 -191.755 203.490 -190.255 ;
        RECT 204.240 -191.755 204.470 -190.255 ;
        RECT 236.025 -190.665 237.715 -190.185 ;
        RECT 282.015 -190.015 282.385 -189.935 ;
        RECT 283.155 -190.015 283.705 -189.835 ;
        RECT 236.025 -190.695 236.395 -190.665 ;
        RECT 237.165 -190.755 237.715 -190.665 ;
        RECT 224.635 -193.105 224.865 -191.605 ;
        RECT 225.615 -193.105 225.845 -191.605 ;
        RECT 226.595 -193.105 226.825 -191.605 ;
        RECT 227.680 -192.100 227.910 -191.600 ;
        RECT 228.660 -192.100 228.890 -191.600 ;
        RECT 229.640 -192.100 229.870 -191.600 ;
        RECT 230.620 -192.100 230.850 -191.600 ;
        RECT 231.870 -194.160 232.100 -191.160 ;
        RECT 232.850 -194.160 233.080 -191.160 ;
        RECT 234.965 -194.160 235.195 -191.160 ;
        RECT 241.830 -192.950 242.060 -190.450 ;
        RECT 242.810 -192.950 243.040 -190.450 ;
        RECT 245.785 -192.950 246.015 -190.450 ;
        RECT 246.435 -192.950 246.665 -190.450 ;
        RECT 247.575 -191.950 247.805 -190.450 ;
        RECT 248.555 -191.950 248.785 -190.450 ;
        RECT 282.015 -190.495 283.705 -190.015 ;
        RECT 325.785 -190.165 327.475 -189.685 ;
        RECT 371.550 -189.600 371.920 -189.520 ;
        RECT 372.690 -189.600 373.240 -189.420 ;
        RECT 325.785 -190.195 326.155 -190.165 ;
        RECT 326.925 -190.255 327.475 -190.165 ;
        RECT 282.015 -190.525 282.385 -190.495 ;
        RECT 283.155 -190.585 283.705 -190.495 ;
        RECT 270.625 -192.935 270.855 -191.435 ;
        RECT 271.605 -192.935 271.835 -191.435 ;
        RECT 272.585 -192.935 272.815 -191.435 ;
        RECT 273.670 -191.930 273.900 -191.430 ;
        RECT 274.650 -191.930 274.880 -191.430 ;
        RECT 275.630 -191.930 275.860 -191.430 ;
        RECT 276.610 -191.930 276.840 -191.430 ;
        RECT 277.860 -193.990 278.090 -190.990 ;
        RECT 278.840 -193.990 279.070 -190.990 ;
        RECT 280.955 -193.990 281.185 -190.990 ;
        RECT 287.820 -192.780 288.050 -190.280 ;
        RECT 288.800 -192.780 289.030 -190.280 ;
        RECT 291.775 -192.780 292.005 -190.280 ;
        RECT 292.425 -192.780 292.655 -190.280 ;
        RECT 293.565 -191.780 293.795 -190.280 ;
        RECT 294.545 -191.780 294.775 -190.280 ;
        RECT 314.395 -192.605 314.625 -191.105 ;
        RECT 315.375 -192.605 315.605 -191.105 ;
        RECT 316.355 -192.605 316.585 -191.105 ;
        RECT 317.440 -191.600 317.670 -191.100 ;
        RECT 318.420 -191.600 318.650 -191.100 ;
        RECT 319.400 -191.600 319.630 -191.100 ;
        RECT 320.380 -191.600 320.610 -191.100 ;
        RECT 321.630 -193.660 321.860 -190.660 ;
        RECT 322.610 -193.660 322.840 -190.660 ;
        RECT 324.725 -193.660 324.955 -190.660 ;
        RECT 331.590 -192.450 331.820 -189.950 ;
        RECT 332.570 -192.450 332.800 -189.950 ;
        RECT 335.545 -192.450 335.775 -189.950 ;
        RECT 336.195 -192.450 336.425 -189.950 ;
        RECT 337.335 -191.450 337.565 -189.950 ;
        RECT 338.315 -191.450 338.545 -189.950 ;
        RECT 371.550 -190.080 373.240 -189.600 ;
        RECT 371.550 -190.110 371.920 -190.080 ;
        RECT 372.690 -190.170 373.240 -190.080 ;
        RECT 360.160 -192.520 360.390 -191.020 ;
        RECT 361.140 -192.520 361.370 -191.020 ;
        RECT 362.120 -192.520 362.350 -191.020 ;
        RECT 363.205 -191.515 363.435 -191.015 ;
        RECT 364.185 -191.515 364.415 -191.015 ;
        RECT 365.165 -191.515 365.395 -191.015 ;
        RECT 366.145 -191.515 366.375 -191.015 ;
        RECT 367.395 -193.575 367.625 -190.575 ;
        RECT 368.375 -193.575 368.605 -190.575 ;
        RECT 370.490 -193.575 370.720 -190.575 ;
        RECT 377.355 -192.365 377.585 -189.865 ;
        RECT 378.335 -192.365 378.565 -189.865 ;
        RECT 381.310 -192.365 381.540 -189.865 ;
        RECT 381.960 -192.365 382.190 -189.865 ;
        RECT 383.100 -191.365 383.330 -189.865 ;
        RECT 384.080 -191.365 384.310 -189.865 ;
        RECT 418.370 -189.890 420.060 -189.410 ;
        RECT 418.370 -189.920 418.740 -189.890 ;
        RECT 419.510 -189.980 420.060 -189.890 ;
        RECT 406.980 -192.330 407.210 -190.830 ;
        RECT 407.960 -192.330 408.190 -190.830 ;
        RECT 408.940 -192.330 409.170 -190.830 ;
        RECT 410.025 -191.325 410.255 -190.825 ;
        RECT 411.005 -191.325 411.235 -190.825 ;
        RECT 411.985 -191.325 412.215 -190.825 ;
        RECT 412.965 -191.325 413.195 -190.825 ;
        RECT 414.215 -193.385 414.445 -190.385 ;
        RECT 415.195 -193.385 415.425 -190.385 ;
        RECT 417.310 -193.385 417.540 -190.385 ;
        RECT 424.175 -192.175 424.405 -189.675 ;
        RECT 425.155 -192.175 425.385 -189.675 ;
        RECT 428.130 -192.175 428.360 -189.675 ;
        RECT 428.780 -192.175 429.010 -189.675 ;
        RECT 429.920 -191.175 430.150 -189.675 ;
        RECT 430.900 -191.175 431.130 -189.675 ;
        RECT -130.060 -195.725 -128.060 -195.495 ;
        RECT 96.960 -196.065 97.190 -195.065 ;
        RECT 97.940 -196.065 98.170 -195.065 ;
        RECT 98.920 -196.065 99.150 -195.065 ;
        RECT 101.370 -196.065 101.600 -195.065 ;
        RECT 102.350 -196.065 102.580 -195.065 ;
        RECT 103.330 -196.065 103.560 -195.065 ;
        RECT 110.085 -196.065 110.315 -195.065 ;
        RECT 111.065 -196.065 111.295 -195.065 ;
        RECT 112.045 -196.065 112.275 -195.065 ;
        RECT 114.870 -196.065 115.100 -195.065 ;
        RECT 115.850 -196.065 116.080 -195.065 ;
        RECT 116.830 -196.065 117.060 -195.065 ;
        RECT 123.585 -196.065 123.815 -195.065 ;
        RECT 124.565 -196.065 124.795 -195.065 ;
        RECT 125.545 -196.065 125.775 -195.065 ;
        RECT -130.060 -196.905 -128.060 -196.675 ;
        RECT -130.060 -198.085 -128.060 -197.855 ;
        RECT -130.060 -199.265 -128.060 -199.035 ;
        RECT -130.060 -199.915 -128.060 -199.685 ;
        RECT -72.235 -200.575 -72.005 -199.575 ;
        RECT -71.255 -200.575 -71.025 -199.575 ;
        RECT -70.275 -200.575 -70.045 -199.575 ;
        RECT -68.050 -200.575 -67.820 -199.575 ;
        RECT -67.070 -200.575 -66.840 -199.575 ;
        RECT -66.090 -200.575 -65.860 -199.575 ;
        RECT -58.735 -200.575 -58.505 -199.575 ;
        RECT -57.755 -200.575 -57.525 -199.575 ;
        RECT -56.775 -200.575 -56.545 -199.575 ;
        RECT -54.550 -200.575 -54.320 -199.575 ;
        RECT -53.570 -200.575 -53.340 -199.575 ;
        RECT -52.590 -200.575 -52.360 -199.575 ;
        RECT -130.060 -201.095 -128.060 -200.865 ;
        RECT -130.060 -202.275 -128.060 -202.045 ;
        RECT -94.360 -203.100 -93.465 -202.265 ;
        RECT -40.290 -202.660 -40.060 -199.660 ;
        RECT -38.175 -202.660 -37.945 -199.660 ;
        RECT -37.195 -202.660 -36.965 -199.660 ;
        RECT 109.185 -200.825 109.415 -198.825 ;
        RECT 110.165 -200.825 110.395 -198.825 ;
        RECT 111.145 -200.825 111.375 -198.825 ;
        RECT -32.865 -201.910 -32.635 -200.910 ;
        RECT -31.885 -201.910 -31.655 -200.910 ;
        RECT -30.905 -201.910 -30.675 -200.910 ;
        RECT -28.680 -201.910 -28.450 -200.910 ;
        RECT -27.700 -201.910 -27.470 -200.910 ;
        RECT -26.720 -201.910 -26.490 -200.910 ;
        RECT -19.365 -201.910 -19.135 -200.910 ;
        RECT -18.385 -201.910 -18.155 -200.910 ;
        RECT -17.405 -201.910 -17.175 -200.910 ;
        RECT -15.180 -201.910 -14.950 -200.910 ;
        RECT -14.200 -201.910 -13.970 -200.910 ;
        RECT -13.220 -201.910 -12.990 -200.910 ;
        RECT -130.060 -203.455 -128.060 -203.225 ;
        RECT -130.060 -204.635 -128.060 -204.405 ;
        RECT -130.060 -205.285 -128.060 -205.055 ;
        RECT -130.060 -206.465 -128.060 -206.235 ;
        RECT -130.060 -207.645 -128.060 -207.415 ;
        RECT -109.620 -208.000 -109.390 -205.000 ;
        RECT -108.640 -208.000 -108.410 -205.000 ;
        RECT -103.590 -206.645 -103.360 -204.645 ;
        RECT -102.610 -206.645 -102.380 -204.645 ;
        RECT -99.065 -206.650 -98.835 -204.650 ;
        RECT -98.085 -206.650 -97.855 -204.650 ;
        RECT -94.225 -211.920 -93.595 -203.100 ;
        RECT -71.745 -207.165 -71.515 -206.165 ;
        RECT -70.765 -207.165 -70.535 -206.165 ;
        RECT -69.785 -207.165 -69.555 -206.165 ;
        RECT -63.030 -207.165 -62.800 -206.165 ;
        RECT -62.050 -207.165 -61.820 -206.165 ;
        RECT -61.070 -207.165 -60.840 -206.165 ;
        RECT -58.245 -207.165 -58.015 -206.165 ;
        RECT -57.265 -207.165 -57.035 -206.165 ;
        RECT -56.285 -207.165 -56.055 -206.165 ;
        RECT -49.530 -207.165 -49.300 -206.165 ;
        RECT -48.550 -207.165 -48.320 -206.165 ;
        RECT -47.570 -207.165 -47.340 -206.165 ;
        RECT -45.120 -207.165 -44.890 -206.165 ;
        RECT -44.140 -207.165 -43.910 -206.165 ;
        RECT -43.160 -207.165 -42.930 -206.165 ;
        RECT -92.055 -210.795 -91.825 -209.295 ;
        RECT -91.075 -210.795 -90.845 -209.295 ;
        RECT -90.095 -210.795 -89.865 -209.295 ;
        RECT -89.010 -210.800 -88.780 -210.300 ;
        RECT -88.030 -210.800 -87.800 -210.300 ;
        RECT -87.050 -210.800 -86.820 -210.300 ;
        RECT -86.070 -210.800 -85.840 -210.300 ;
        RECT -84.820 -211.240 -84.590 -208.240 ;
        RECT -83.840 -211.240 -83.610 -208.240 ;
        RECT -81.725 -211.240 -81.495 -208.240 ;
        RECT -32.375 -208.500 -32.145 -207.500 ;
        RECT -31.395 -208.500 -31.165 -207.500 ;
        RECT -30.415 -208.500 -30.185 -207.500 ;
        RECT -23.660 -208.500 -23.430 -207.500 ;
        RECT -22.680 -208.500 -22.450 -207.500 ;
        RECT -21.700 -208.500 -21.470 -207.500 ;
        RECT -18.875 -208.500 -18.645 -207.500 ;
        RECT -17.895 -208.500 -17.665 -207.500 ;
        RECT -16.915 -208.500 -16.685 -207.500 ;
        RECT -10.160 -208.500 -9.930 -207.500 ;
        RECT -9.180 -208.500 -8.950 -207.500 ;
        RECT -8.200 -208.500 -7.970 -207.500 ;
        RECT -5.750 -208.500 -5.520 -207.500 ;
        RECT -4.770 -208.500 -4.540 -207.500 ;
        RECT -3.790 -208.500 -3.560 -207.500 ;
        RECT -2.080 -208.415 -1.850 -207.415 ;
        RECT -1.100 -208.415 -0.870 -207.415 ;
        RECT 1.610 -208.415 1.840 -207.415 ;
        RECT 2.590 -208.415 2.820 -207.415 ;
        RECT 3.570 -208.415 3.800 -207.415 ;
        RECT 4.550 -208.415 4.780 -207.415 ;
        RECT 6.585 -208.350 6.815 -207.850 ;
        RECT 7.565 -208.350 7.795 -207.850 ;
        RECT 8.545 -208.350 8.775 -207.850 ;
        RECT 9.525 -208.350 9.755 -207.850 ;
        RECT 10.610 -208.345 10.840 -206.845 ;
        RECT 11.590 -208.345 11.820 -206.845 ;
        RECT 12.570 -208.345 12.800 -206.845 ;
        RECT 14.610 -208.340 14.840 -207.840 ;
        RECT 15.590 -208.340 15.820 -207.840 ;
        RECT 16.570 -208.340 16.800 -207.840 ;
        RECT 17.550 -208.340 17.780 -207.840 ;
        RECT 18.635 -208.335 18.865 -206.835 ;
        RECT 19.615 -208.335 19.845 -206.835 ;
        RECT 20.595 -208.335 20.825 -206.835 ;
        RECT 90.330 -207.195 90.560 -205.195 ;
        RECT 91.310 -207.195 91.540 -205.195 ;
        RECT 95.060 -207.195 95.290 -205.195 ;
        RECT 96.040 -207.195 96.270 -205.195 ;
        RECT 99.640 -207.365 99.870 -206.365 ;
        RECT 100.620 -207.365 100.850 -206.365 ;
        RECT 101.600 -207.365 101.830 -206.365 ;
        RECT 102.580 -207.365 102.810 -206.365 ;
        RECT 105.290 -207.365 105.520 -206.365 ;
        RECT 106.270 -207.365 106.500 -206.365 ;
        RECT 108.935 -207.330 109.165 -206.330 ;
        RECT 109.915 -207.330 110.145 -206.330 ;
        RECT 110.895 -207.330 111.125 -206.330 ;
        RECT 113.335 -206.975 113.565 -203.475 ;
        RECT 114.315 -206.975 114.545 -203.475 ;
        RECT 115.335 -206.975 115.565 -203.475 ;
        RECT 116.315 -206.975 116.545 -203.475 ;
        RECT 118.335 -206.975 118.565 -203.475 ;
        RECT 119.315 -206.975 119.545 -203.475 ;
        RECT 120.335 -206.975 120.565 -203.475 ;
        RECT 121.315 -206.975 121.545 -203.475 ;
        RECT 123.335 -206.975 123.565 -203.475 ;
        RECT 124.315 -206.975 124.545 -203.475 ;
        RECT 125.335 -206.975 125.565 -203.475 ;
        RECT 126.315 -206.975 126.545 -203.475 ;
        RECT 138.210 -204.975 138.440 -203.975 ;
        RECT 139.190 -204.975 139.420 -203.975 ;
        RECT 140.170 -204.975 140.400 -203.975 ;
        RECT 141.150 -204.975 141.380 -203.975 ;
        RECT 143.075 -205.620 143.305 -204.120 ;
        RECT 144.055 -205.620 144.285 -204.120 ;
        RECT 145.035 -205.620 145.265 -204.120 ;
        RECT 146.120 -205.625 146.350 -205.125 ;
        RECT 147.100 -205.625 147.330 -205.125 ;
        RECT 148.080 -205.625 148.310 -205.125 ;
        RECT 149.060 -205.625 149.290 -205.125 ;
        RECT 156.550 -205.130 156.780 -204.130 ;
        RECT 157.530 -205.130 157.760 -204.130 ;
        RECT 158.510 -205.130 158.740 -204.130 ;
        RECT 159.490 -205.130 159.720 -204.130 ;
        RECT 161.415 -205.775 161.645 -204.275 ;
        RECT 162.395 -205.775 162.625 -204.275 ;
        RECT 163.375 -205.775 163.605 -204.275 ;
        RECT 180.410 -205.030 180.640 -204.030 ;
        RECT 181.390 -205.030 181.620 -204.030 ;
        RECT 182.370 -205.030 182.600 -204.030 ;
        RECT 183.350 -205.030 183.580 -204.030 ;
        RECT 164.460 -205.780 164.690 -205.280 ;
        RECT 165.440 -205.780 165.670 -205.280 ;
        RECT 166.420 -205.780 166.650 -205.280 ;
        RECT 167.400 -205.780 167.630 -205.280 ;
        RECT 185.275 -205.675 185.505 -204.175 ;
        RECT 186.255 -205.675 186.485 -204.175 ;
        RECT 187.235 -205.675 187.465 -204.175 ;
        RECT 188.320 -205.680 188.550 -205.180 ;
        RECT 189.300 -205.680 189.530 -205.180 ;
        RECT 190.280 -205.680 190.510 -205.180 ;
        RECT 191.260 -205.680 191.490 -205.180 ;
        RECT 198.750 -205.185 198.980 -204.185 ;
        RECT 199.730 -205.185 199.960 -204.185 ;
        RECT 200.710 -205.185 200.940 -204.185 ;
        RECT 201.690 -205.185 201.920 -204.185 ;
        RECT 203.615 -205.830 203.845 -204.330 ;
        RECT 204.595 -205.830 204.825 -204.330 ;
        RECT 205.575 -205.830 205.805 -204.330 ;
        RECT 224.725 -205.225 224.955 -204.225 ;
        RECT 225.705 -205.225 225.935 -204.225 ;
        RECT 226.685 -205.225 226.915 -204.225 ;
        RECT 227.665 -205.225 227.895 -204.225 ;
        RECT 206.660 -205.835 206.890 -205.335 ;
        RECT 207.640 -205.835 207.870 -205.335 ;
        RECT 208.620 -205.835 208.850 -205.335 ;
        RECT 209.600 -205.835 209.830 -205.335 ;
        RECT 229.590 -205.870 229.820 -204.370 ;
        RECT 230.570 -205.870 230.800 -204.370 ;
        RECT 231.550 -205.870 231.780 -204.370 ;
        RECT 232.635 -205.875 232.865 -205.375 ;
        RECT 233.615 -205.875 233.845 -205.375 ;
        RECT 234.595 -205.875 234.825 -205.375 ;
        RECT 235.575 -205.875 235.805 -205.375 ;
        RECT 243.065 -205.380 243.295 -204.380 ;
        RECT 244.045 -205.380 244.275 -204.380 ;
        RECT 245.025 -205.380 245.255 -204.380 ;
        RECT 246.005 -205.380 246.235 -204.380 ;
        RECT 247.930 -206.025 248.160 -204.525 ;
        RECT 248.910 -206.025 249.140 -204.525 ;
        RECT 249.890 -206.025 250.120 -204.525 ;
        RECT 270.715 -205.055 270.945 -204.055 ;
        RECT 271.695 -205.055 271.925 -204.055 ;
        RECT 272.675 -205.055 272.905 -204.055 ;
        RECT 273.655 -205.055 273.885 -204.055 ;
        RECT 250.975 -206.030 251.205 -205.530 ;
        RECT 251.955 -206.030 252.185 -205.530 ;
        RECT 252.935 -206.030 253.165 -205.530 ;
        RECT 253.915 -206.030 254.145 -205.530 ;
        RECT 275.580 -205.700 275.810 -204.200 ;
        RECT 276.560 -205.700 276.790 -204.200 ;
        RECT 277.540 -205.700 277.770 -204.200 ;
        RECT 278.625 -205.705 278.855 -205.205 ;
        RECT 279.605 -205.705 279.835 -205.205 ;
        RECT 280.585 -205.705 280.815 -205.205 ;
        RECT 281.565 -205.705 281.795 -205.205 ;
        RECT 289.055 -205.210 289.285 -204.210 ;
        RECT 290.035 -205.210 290.265 -204.210 ;
        RECT 291.015 -205.210 291.245 -204.210 ;
        RECT 291.995 -205.210 292.225 -204.210 ;
        RECT 293.920 -205.855 294.150 -204.355 ;
        RECT 294.900 -205.855 295.130 -204.355 ;
        RECT 295.880 -205.855 296.110 -204.355 ;
        RECT 314.485 -204.725 314.715 -203.725 ;
        RECT 315.465 -204.725 315.695 -203.725 ;
        RECT 316.445 -204.725 316.675 -203.725 ;
        RECT 317.425 -204.725 317.655 -203.725 ;
        RECT 296.965 -205.860 297.195 -205.360 ;
        RECT 297.945 -205.860 298.175 -205.360 ;
        RECT 298.925 -205.860 299.155 -205.360 ;
        RECT 299.905 -205.860 300.135 -205.360 ;
        RECT 319.350 -205.370 319.580 -203.870 ;
        RECT 320.330 -205.370 320.560 -203.870 ;
        RECT 321.310 -205.370 321.540 -203.870 ;
        RECT 322.395 -205.375 322.625 -204.875 ;
        RECT 323.375 -205.375 323.605 -204.875 ;
        RECT 324.355 -205.375 324.585 -204.875 ;
        RECT 325.335 -205.375 325.565 -204.875 ;
        RECT 332.825 -204.880 333.055 -203.880 ;
        RECT 333.805 -204.880 334.035 -203.880 ;
        RECT 334.785 -204.880 335.015 -203.880 ;
        RECT 335.765 -204.880 335.995 -203.880 ;
        RECT 337.690 -205.525 337.920 -204.025 ;
        RECT 338.670 -205.525 338.900 -204.025 ;
        RECT 339.650 -205.525 339.880 -204.025 ;
        RECT 360.250 -204.640 360.480 -203.640 ;
        RECT 361.230 -204.640 361.460 -203.640 ;
        RECT 362.210 -204.640 362.440 -203.640 ;
        RECT 363.190 -204.640 363.420 -203.640 ;
        RECT 340.735 -205.530 340.965 -205.030 ;
        RECT 341.715 -205.530 341.945 -205.030 ;
        RECT 342.695 -205.530 342.925 -205.030 ;
        RECT 343.675 -205.530 343.905 -205.030 ;
        RECT 365.115 -205.285 365.345 -203.785 ;
        RECT 366.095 -205.285 366.325 -203.785 ;
        RECT 367.075 -205.285 367.305 -203.785 ;
        RECT 368.160 -205.290 368.390 -204.790 ;
        RECT 369.140 -205.290 369.370 -204.790 ;
        RECT 370.120 -205.290 370.350 -204.790 ;
        RECT 371.100 -205.290 371.330 -204.790 ;
        RECT 378.590 -204.795 378.820 -203.795 ;
        RECT 379.570 -204.795 379.800 -203.795 ;
        RECT 380.550 -204.795 380.780 -203.795 ;
        RECT 381.530 -204.795 381.760 -203.795 ;
        RECT 383.455 -205.440 383.685 -203.940 ;
        RECT 384.435 -205.440 384.665 -203.940 ;
        RECT 385.415 -205.440 385.645 -203.940 ;
        RECT 407.070 -204.450 407.300 -203.450 ;
        RECT 408.050 -204.450 408.280 -203.450 ;
        RECT 409.030 -204.450 409.260 -203.450 ;
        RECT 410.010 -204.450 410.240 -203.450 ;
        RECT 386.500 -205.445 386.730 -204.945 ;
        RECT 387.480 -205.445 387.710 -204.945 ;
        RECT 388.460 -205.445 388.690 -204.945 ;
        RECT 389.440 -205.445 389.670 -204.945 ;
        RECT 411.935 -205.095 412.165 -203.595 ;
        RECT 412.915 -205.095 413.145 -203.595 ;
        RECT 413.895 -205.095 414.125 -203.595 ;
        RECT 414.980 -205.100 415.210 -204.600 ;
        RECT 415.960 -205.100 416.190 -204.600 ;
        RECT 416.940 -205.100 417.170 -204.600 ;
        RECT 417.920 -205.100 418.150 -204.600 ;
        RECT 425.410 -204.605 425.640 -203.605 ;
        RECT 426.390 -204.605 426.620 -203.605 ;
        RECT 427.370 -204.605 427.600 -203.605 ;
        RECT 428.350 -204.605 428.580 -203.605 ;
        RECT 430.275 -205.250 430.505 -203.750 ;
        RECT 431.255 -205.250 431.485 -203.750 ;
        RECT 432.235 -205.250 432.465 -203.750 ;
        RECT 433.320 -205.255 433.550 -204.755 ;
        RECT 434.300 -205.255 434.530 -204.755 ;
        RECT 435.280 -205.255 435.510 -204.755 ;
        RECT 436.260 -205.255 436.490 -204.755 ;
        RECT 320.360 -206.745 321.275 -206.540 ;
        RECT 326.875 -206.745 327.355 -206.600 ;
        RECT 366.125 -206.660 367.040 -206.455 ;
        RECT 412.945 -206.470 413.860 -206.265 ;
        RECT 419.460 -206.470 419.940 -206.325 ;
        RECT 372.640 -206.660 373.120 -206.515 ;
        RECT 144.085 -206.995 145.000 -206.790 ;
        RECT 150.600 -206.995 151.080 -206.850 ;
        RECT 144.085 -207.405 151.080 -206.995 ;
        RECT 22.730 -208.460 22.960 -207.460 ;
        RECT 23.710 -208.460 23.940 -207.460 ;
        RECT 26.420 -208.460 26.650 -207.460 ;
        RECT 27.400 -208.460 27.630 -207.460 ;
        RECT 28.380 -208.460 28.610 -207.460 ;
        RECT 29.360 -208.460 29.590 -207.460 ;
        RECT 35.165 -208.405 35.395 -207.405 ;
        RECT 36.145 -208.405 36.375 -207.405 ;
        RECT 37.125 -208.405 37.355 -207.405 ;
        RECT 37.695 -208.405 37.925 -207.405 ;
        RECT 38.675 -208.405 38.905 -207.405 ;
        RECT 39.240 -208.405 39.470 -207.405 ;
        RECT 40.220 -208.405 40.450 -207.405 ;
        RECT 144.085 -207.440 145.000 -207.405 ;
        RECT 150.600 -207.535 151.080 -207.405 ;
        RECT 167.700 -207.105 168.155 -207.045 ;
        RECT 168.950 -207.105 169.705 -206.970 ;
        RECT 167.700 -207.800 169.705 -207.105 ;
        RECT 186.285 -207.050 187.200 -206.845 ;
        RECT 192.800 -207.050 193.280 -206.905 ;
        RECT 186.285 -207.460 193.280 -207.050 ;
        RECT 186.285 -207.495 187.200 -207.460 ;
        RECT 192.800 -207.590 193.280 -207.460 ;
        RECT 209.900 -207.160 210.355 -207.100 ;
        RECT 211.150 -207.160 211.905 -207.025 ;
        RECT 167.700 -207.860 168.155 -207.800 ;
        RECT 168.950 -207.925 169.705 -207.800 ;
        RECT 209.900 -207.855 211.905 -207.160 ;
        RECT 230.600 -207.245 231.515 -207.040 ;
        RECT 276.590 -207.075 277.505 -206.870 ;
        RECT 283.105 -207.075 283.585 -206.930 ;
        RECT 237.115 -207.245 237.595 -207.100 ;
        RECT 230.600 -207.655 237.595 -207.245 ;
        RECT 230.600 -207.690 231.515 -207.655 ;
        RECT 237.115 -207.785 237.595 -207.655 ;
        RECT 254.215 -207.355 254.670 -207.295 ;
        RECT 255.465 -207.355 256.220 -207.220 ;
        RECT 209.900 -207.915 210.355 -207.855 ;
        RECT 211.150 -207.980 211.905 -207.855 ;
        RECT 254.215 -208.050 256.220 -207.355 ;
        RECT 276.590 -207.485 283.585 -207.075 ;
        RECT 276.590 -207.520 277.505 -207.485 ;
        RECT 283.105 -207.615 283.585 -207.485 ;
        RECT 300.205 -207.185 300.660 -207.125 ;
        RECT 301.455 -207.185 302.210 -207.050 ;
        RECT 300.205 -207.880 302.210 -207.185 ;
        RECT 320.360 -207.155 327.355 -206.745 ;
        RECT 320.360 -207.190 321.275 -207.155 ;
        RECT 326.875 -207.285 327.355 -207.155 ;
        RECT 343.975 -206.855 344.430 -206.795 ;
        RECT 345.225 -206.855 345.980 -206.720 ;
        RECT 343.975 -207.550 345.980 -206.855 ;
        RECT 366.125 -207.070 373.120 -206.660 ;
        RECT 366.125 -207.105 367.040 -207.070 ;
        RECT 372.640 -207.200 373.120 -207.070 ;
        RECT 389.740 -206.770 390.195 -206.710 ;
        RECT 390.990 -206.770 391.745 -206.635 ;
        RECT 389.740 -207.465 391.745 -206.770 ;
        RECT 412.945 -206.880 419.940 -206.470 ;
        RECT 412.945 -206.915 413.860 -206.880 ;
        RECT 419.460 -207.010 419.940 -206.880 ;
        RECT 436.560 -206.580 437.015 -206.520 ;
        RECT 437.810 -206.580 438.565 -206.445 ;
        RECT 436.560 -207.275 438.565 -206.580 ;
        RECT 436.560 -207.335 437.015 -207.275 ;
        RECT 437.810 -207.400 438.565 -207.275 ;
        RECT 389.740 -207.525 390.195 -207.465 ;
        RECT 343.975 -207.610 344.430 -207.550 ;
        RECT 345.225 -207.675 345.980 -207.550 ;
        RECT 390.990 -207.590 391.745 -207.465 ;
        RECT 300.205 -207.940 300.660 -207.880 ;
        RECT 301.455 -208.005 302.210 -207.880 ;
        RECT 254.215 -208.110 254.670 -208.050 ;
        RECT 255.465 -208.175 256.220 -208.050 ;
        RECT -4.120 -208.750 -3.505 -208.705 ;
        RECT -2.650 -208.750 -2.035 -208.710 ;
        RECT -4.120 -209.325 -2.035 -208.750 ;
        RECT 12.240 -208.715 12.855 -208.645 ;
        RECT 14.185 -208.715 14.800 -208.650 ;
        RECT 12.240 -209.250 14.800 -208.715 ;
        RECT 12.240 -209.325 12.855 -209.250 ;
        RECT -4.120 -209.385 -3.505 -209.325 ;
        RECT -2.650 -209.390 -2.035 -209.325 ;
        RECT 14.185 -209.330 14.800 -209.250 ;
        RECT 20.325 -208.865 20.940 -208.765 ;
        RECT 22.330 -208.865 22.945 -208.775 ;
        RECT 20.325 -209.400 22.945 -208.865 ;
        RECT 20.325 -209.445 20.940 -209.400 ;
        RECT 22.330 -209.455 22.945 -209.400 ;
        RECT 29.110 -208.840 29.725 -208.750 ;
        RECT 35.190 -208.840 35.805 -208.745 ;
        RECT 29.110 -209.365 35.805 -208.840 ;
        RECT 29.110 -209.430 29.725 -209.365 ;
        RECT 35.190 -209.425 35.805 -209.365 ;
        RECT 138.080 -210.120 138.310 -208.620 ;
        RECT 139.060 -210.120 139.290 -208.620 ;
        RECT 140.040 -210.120 140.270 -208.620 ;
        RECT 141.125 -209.115 141.355 -208.615 ;
        RECT 142.105 -209.115 142.335 -208.615 ;
        RECT 143.085 -209.115 143.315 -208.615 ;
        RECT 144.065 -209.115 144.295 -208.615 ;
        RECT 145.315 -211.175 145.545 -208.175 ;
        RECT 146.295 -211.175 146.525 -208.175 ;
        RECT 148.410 -211.175 148.640 -208.175 ;
        RECT 156.420 -210.275 156.650 -208.775 ;
        RECT 157.400 -210.275 157.630 -208.775 ;
        RECT 158.380 -210.275 158.610 -208.775 ;
        RECT 159.465 -209.270 159.695 -208.770 ;
        RECT 160.445 -209.270 160.675 -208.770 ;
        RECT 161.425 -209.270 161.655 -208.770 ;
        RECT 162.405 -209.270 162.635 -208.770 ;
        RECT -94.230 -212.780 -93.270 -211.920 ;
        RECT -23.250 -212.715 -22.635 -212.035 ;
        RECT 56.320 -212.255 56.550 -211.255 ;
        RECT 57.300 -212.255 57.530 -211.255 ;
        RECT 58.280 -212.255 58.510 -211.255 ;
        RECT 60.730 -212.255 60.960 -211.255 ;
        RECT 61.710 -212.255 61.940 -211.255 ;
        RECT 62.690 -212.255 62.920 -211.255 ;
        RECT 69.445 -212.255 69.675 -211.255 ;
        RECT 70.425 -212.255 70.655 -211.255 ;
        RECT 71.405 -212.255 71.635 -211.255 ;
        RECT 74.230 -212.255 74.460 -211.255 ;
        RECT 75.210 -212.255 75.440 -211.255 ;
        RECT 76.190 -212.255 76.420 -211.255 ;
        RECT 82.945 -212.255 83.175 -211.255 ;
        RECT 83.925 -212.255 84.155 -211.255 ;
        RECT 84.905 -212.255 85.135 -211.255 ;
        RECT 163.655 -211.330 163.885 -208.330 ;
        RECT 164.635 -211.330 164.865 -208.330 ;
        RECT 166.750 -211.330 166.980 -208.330 ;
        RECT 180.280 -210.175 180.510 -208.675 ;
        RECT 181.260 -210.175 181.490 -208.675 ;
        RECT 182.240 -210.175 182.470 -208.675 ;
        RECT 183.325 -209.170 183.555 -208.670 ;
        RECT 184.305 -209.170 184.535 -208.670 ;
        RECT 185.285 -209.170 185.515 -208.670 ;
        RECT 186.265 -209.170 186.495 -208.670 ;
        RECT 187.515 -211.230 187.745 -208.230 ;
        RECT 188.495 -211.230 188.725 -208.230 ;
        RECT 190.610 -211.230 190.840 -208.230 ;
        RECT 198.620 -210.330 198.850 -208.830 ;
        RECT 199.600 -210.330 199.830 -208.830 ;
        RECT 200.580 -210.330 200.810 -208.830 ;
        RECT 201.665 -209.325 201.895 -208.825 ;
        RECT 202.645 -209.325 202.875 -208.825 ;
        RECT 203.625 -209.325 203.855 -208.825 ;
        RECT 204.605 -209.325 204.835 -208.825 ;
        RECT 205.855 -211.385 206.085 -208.385 ;
        RECT 206.835 -211.385 207.065 -208.385 ;
        RECT 208.950 -211.385 209.180 -208.385 ;
        RECT 224.595 -210.370 224.825 -208.870 ;
        RECT 225.575 -210.370 225.805 -208.870 ;
        RECT 226.555 -210.370 226.785 -208.870 ;
        RECT 227.640 -209.365 227.870 -208.865 ;
        RECT 228.620 -209.365 228.850 -208.865 ;
        RECT 229.600 -209.365 229.830 -208.865 ;
        RECT 230.580 -209.365 230.810 -208.865 ;
        RECT 231.830 -211.425 232.060 -208.425 ;
        RECT 232.810 -211.425 233.040 -208.425 ;
        RECT 234.925 -211.425 235.155 -208.425 ;
        RECT 242.935 -210.525 243.165 -209.025 ;
        RECT 243.915 -210.525 244.145 -209.025 ;
        RECT 244.895 -210.525 245.125 -209.025 ;
        RECT 245.980 -209.520 246.210 -209.020 ;
        RECT 246.960 -209.520 247.190 -209.020 ;
        RECT 247.940 -209.520 248.170 -209.020 ;
        RECT 248.920 -209.520 249.150 -209.020 ;
        RECT 250.170 -211.580 250.400 -208.580 ;
        RECT 251.150 -211.580 251.380 -208.580 ;
        RECT 253.265 -211.580 253.495 -208.580 ;
        RECT 270.585 -210.200 270.815 -208.700 ;
        RECT 271.565 -210.200 271.795 -208.700 ;
        RECT 272.545 -210.200 272.775 -208.700 ;
        RECT 273.630 -209.195 273.860 -208.695 ;
        RECT 274.610 -209.195 274.840 -208.695 ;
        RECT 275.590 -209.195 275.820 -208.695 ;
        RECT 276.570 -209.195 276.800 -208.695 ;
        RECT 277.820 -211.255 278.050 -208.255 ;
        RECT 278.800 -211.255 279.030 -208.255 ;
        RECT 280.915 -211.255 281.145 -208.255 ;
        RECT 288.925 -210.355 289.155 -208.855 ;
        RECT 289.905 -210.355 290.135 -208.855 ;
        RECT 290.885 -210.355 291.115 -208.855 ;
        RECT 291.970 -209.350 292.200 -208.850 ;
        RECT 292.950 -209.350 293.180 -208.850 ;
        RECT 293.930 -209.350 294.160 -208.850 ;
        RECT 294.910 -209.350 295.140 -208.850 ;
        RECT 296.160 -211.410 296.390 -208.410 ;
        RECT 297.140 -211.410 297.370 -208.410 ;
        RECT 299.255 -211.410 299.485 -208.410 ;
        RECT 314.355 -209.870 314.585 -208.370 ;
        RECT 315.335 -209.870 315.565 -208.370 ;
        RECT 316.315 -209.870 316.545 -208.370 ;
        RECT 317.400 -208.865 317.630 -208.365 ;
        RECT 318.380 -208.865 318.610 -208.365 ;
        RECT 319.360 -208.865 319.590 -208.365 ;
        RECT 320.340 -208.865 320.570 -208.365 ;
        RECT 321.590 -210.925 321.820 -207.925 ;
        RECT 322.570 -210.925 322.800 -207.925 ;
        RECT 324.685 -210.925 324.915 -207.925 ;
        RECT 332.695 -210.025 332.925 -208.525 ;
        RECT 333.675 -210.025 333.905 -208.525 ;
        RECT 334.655 -210.025 334.885 -208.525 ;
        RECT 335.740 -209.020 335.970 -208.520 ;
        RECT 336.720 -209.020 336.950 -208.520 ;
        RECT 337.700 -209.020 337.930 -208.520 ;
        RECT 338.680 -209.020 338.910 -208.520 ;
        RECT 339.930 -211.080 340.160 -208.080 ;
        RECT 340.910 -211.080 341.140 -208.080 ;
        RECT 343.025 -211.080 343.255 -208.080 ;
        RECT 360.120 -209.785 360.350 -208.285 ;
        RECT 361.100 -209.785 361.330 -208.285 ;
        RECT 362.080 -209.785 362.310 -208.285 ;
        RECT 363.165 -208.780 363.395 -208.280 ;
        RECT 364.145 -208.780 364.375 -208.280 ;
        RECT 365.125 -208.780 365.355 -208.280 ;
        RECT 366.105 -208.780 366.335 -208.280 ;
        RECT 367.355 -210.840 367.585 -207.840 ;
        RECT 368.335 -210.840 368.565 -207.840 ;
        RECT 370.450 -210.840 370.680 -207.840 ;
        RECT 378.460 -209.940 378.690 -208.440 ;
        RECT 379.440 -209.940 379.670 -208.440 ;
        RECT 380.420 -209.940 380.650 -208.440 ;
        RECT 381.505 -208.935 381.735 -208.435 ;
        RECT 382.485 -208.935 382.715 -208.435 ;
        RECT 383.465 -208.935 383.695 -208.435 ;
        RECT 384.445 -208.935 384.675 -208.435 ;
        RECT 385.695 -210.995 385.925 -207.995 ;
        RECT 386.675 -210.995 386.905 -207.995 ;
        RECT 388.790 -210.995 389.020 -207.995 ;
        RECT 406.940 -209.595 407.170 -208.095 ;
        RECT 407.920 -209.595 408.150 -208.095 ;
        RECT 408.900 -209.595 409.130 -208.095 ;
        RECT 409.985 -208.590 410.215 -208.090 ;
        RECT 410.965 -208.590 411.195 -208.090 ;
        RECT 411.945 -208.590 412.175 -208.090 ;
        RECT 412.925 -208.590 413.155 -208.090 ;
        RECT 414.175 -210.650 414.405 -207.650 ;
        RECT 415.155 -210.650 415.385 -207.650 ;
        RECT 417.270 -210.650 417.500 -207.650 ;
        RECT 425.280 -209.750 425.510 -208.250 ;
        RECT 426.260 -209.750 426.490 -208.250 ;
        RECT 427.240 -209.750 427.470 -208.250 ;
        RECT 428.325 -208.745 428.555 -208.245 ;
        RECT 429.305 -208.745 429.535 -208.245 ;
        RECT 430.285 -208.745 430.515 -208.245 ;
        RECT 431.265 -208.745 431.495 -208.245 ;
        RECT 432.515 -210.805 432.745 -207.805 ;
        RECT 433.495 -210.805 433.725 -207.805 ;
        RECT 435.610 -210.805 435.840 -207.805 ;
        RECT -91.925 -215.440 -91.695 -214.440 ;
        RECT -90.945 -215.440 -90.715 -214.440 ;
        RECT -89.965 -215.440 -89.735 -214.440 ;
        RECT -88.985 -215.440 -88.755 -214.440 ;
        RECT -87.060 -215.295 -86.830 -213.795 ;
        RECT -86.080 -215.295 -85.850 -213.795 ;
        RECT -85.100 -215.295 -84.870 -213.795 ;
        RECT -84.015 -214.290 -83.785 -213.790 ;
        RECT -83.035 -214.290 -82.805 -213.790 ;
        RECT -82.055 -214.290 -81.825 -213.790 ;
        RECT -81.075 -214.290 -80.845 -213.790 ;
        RECT -23.225 -215.870 -22.655 -212.715 ;
        RECT -10.415 -213.435 -9.800 -212.755 ;
        RECT -10.390 -215.695 -9.820 -213.435 ;
        RECT 2.000 -213.605 3.530 -213.295 ;
        RECT 2.000 -213.610 2.615 -213.605 ;
        RECT 2.025 -215.695 2.595 -213.610 ;
        RECT -23.245 -216.550 -22.630 -215.870 ;
        RECT -10.410 -216.375 -9.795 -215.695 ;
        RECT 2.005 -216.375 2.620 -215.695 ;
        RECT -111.305 -220.090 -111.075 -219.090 ;
        RECT -110.325 -220.090 -110.095 -219.090 ;
        RECT -107.615 -220.090 -107.385 -219.090 ;
        RECT -106.635 -220.090 -106.405 -219.090 ;
        RECT -105.655 -220.090 -105.425 -219.090 ;
        RECT -104.675 -220.090 -104.445 -219.090 ;
        RECT -98.255 -220.910 -97.375 -217.755 ;
        RECT -29.885 -219.660 -29.655 -218.660 ;
        RECT -28.905 -219.660 -28.675 -218.660 ;
        RECT -27.925 -219.660 -27.695 -218.660 ;
        RECT -27.355 -219.660 -27.125 -218.660 ;
        RECT -26.375 -219.660 -26.145 -218.660 ;
        RECT -25.810 -219.660 -25.580 -218.660 ;
        RECT -24.830 -219.660 -24.600 -218.660 ;
        RECT -17.385 -219.660 -17.155 -218.660 ;
        RECT -16.405 -219.660 -16.175 -218.660 ;
        RECT -15.425 -219.660 -15.195 -218.660 ;
        RECT -14.855 -219.660 -14.625 -218.660 ;
        RECT -13.875 -219.660 -13.645 -218.660 ;
        RECT -13.310 -219.660 -13.080 -218.660 ;
        RECT -12.330 -219.660 -12.100 -218.660 ;
        RECT -4.885 -219.660 -4.655 -218.660 ;
        RECT -3.905 -219.660 -3.675 -218.660 ;
        RECT -2.925 -219.660 -2.695 -218.660 ;
        RECT -2.355 -219.660 -2.125 -218.660 ;
        RECT -1.375 -219.660 -1.145 -218.660 ;
        RECT -0.810 -219.660 -0.580 -218.660 ;
        RECT 0.170 -219.660 0.400 -218.660 ;
        RECT 7.615 -219.660 7.845 -218.660 ;
        RECT 8.595 -219.660 8.825 -218.660 ;
        RECT 9.575 -219.660 9.805 -218.660 ;
        RECT 10.145 -219.660 10.375 -218.660 ;
        RECT 11.125 -219.660 11.355 -218.660 ;
        RECT 11.690 -219.660 11.920 -218.660 ;
        RECT 12.670 -219.660 12.900 -218.660 ;
        RECT 20.115 -219.660 20.345 -218.660 ;
        RECT 21.095 -219.660 21.325 -218.660 ;
        RECT 22.075 -219.660 22.305 -218.660 ;
        RECT 22.645 -219.660 22.875 -218.660 ;
        RECT 23.625 -219.660 23.855 -218.660 ;
        RECT 24.190 -219.660 24.420 -218.660 ;
        RECT 25.170 -219.660 25.400 -218.660 ;
        RECT 35.115 -219.660 35.345 -218.660 ;
        RECT 36.095 -219.660 36.325 -218.660 ;
        RECT 37.075 -219.660 37.305 -218.660 ;
        RECT 37.645 -219.660 37.875 -218.660 ;
        RECT 38.625 -219.660 38.855 -218.660 ;
        RECT 39.190 -219.660 39.420 -218.660 ;
        RECT 40.170 -219.660 40.400 -218.660 ;
        RECT 65.750 -218.845 65.980 -217.845 ;
        RECT 66.730 -218.845 66.960 -217.845 ;
        RECT 67.710 -218.845 67.940 -217.845 ;
        RECT 69.935 -218.845 70.165 -217.845 ;
        RECT 70.915 -218.845 71.145 -217.845 ;
        RECT 71.895 -218.845 72.125 -217.845 ;
        RECT 79.250 -218.845 79.480 -217.845 ;
        RECT 80.230 -218.845 80.460 -217.845 ;
        RECT 81.210 -218.845 81.440 -217.845 ;
        RECT 83.435 -218.845 83.665 -217.845 ;
        RECT 84.415 -218.845 84.645 -217.845 ;
        RECT 85.395 -218.845 85.625 -217.845 ;
        RECT -139.160 -261.610 -137.160 -261.380 ;
        RECT -139.160 -262.790 -137.160 -262.560 ;
        RECT -139.160 -263.970 -137.160 -263.740 ;
        RECT -139.160 -265.150 -137.160 -264.920 ;
        RECT -139.160 -266.330 -137.160 -266.100 ;
        RECT -68.720 -266.495 -68.490 -265.495 ;
        RECT -67.740 -266.495 -67.510 -265.495 ;
        RECT -66.760 -266.495 -66.530 -265.495 ;
        RECT -64.535 -266.495 -64.305 -265.495 ;
        RECT -63.555 -266.495 -63.325 -265.495 ;
        RECT -62.575 -266.495 -62.345 -265.495 ;
        RECT -55.220 -266.495 -54.990 -265.495 ;
        RECT -54.240 -266.495 -54.010 -265.495 ;
        RECT -53.260 -266.495 -53.030 -265.495 ;
        RECT -51.035 -266.495 -50.805 -265.495 ;
        RECT -50.055 -266.495 -49.825 -265.495 ;
        RECT -49.075 -266.495 -48.845 -265.495 ;
        RECT -139.160 -267.510 -137.160 -267.280 ;
        RECT -139.160 -268.690 -137.160 -268.460 ;
        RECT -36.910 -268.545 -36.680 -265.545 ;
        RECT -34.795 -268.545 -34.565 -265.545 ;
        RECT -33.815 -268.545 -33.585 -265.545 ;
        RECT -26.370 -267.525 -26.140 -266.525 ;
        RECT -25.390 -267.525 -25.160 -266.525 ;
        RECT -24.410 -267.525 -24.180 -266.525 ;
        RECT -23.840 -267.525 -23.610 -266.525 ;
        RECT -22.860 -267.525 -22.630 -266.525 ;
        RECT -22.295 -267.525 -22.065 -266.525 ;
        RECT -21.315 -267.525 -21.085 -266.525 ;
        RECT -13.870 -267.525 -13.640 -266.525 ;
        RECT -12.890 -267.525 -12.660 -266.525 ;
        RECT -11.910 -267.525 -11.680 -266.525 ;
        RECT -11.340 -267.525 -11.110 -266.525 ;
        RECT -10.360 -267.525 -10.130 -266.525 ;
        RECT -9.795 -267.525 -9.565 -266.525 ;
        RECT -8.815 -267.525 -8.585 -266.525 ;
        RECT -1.370 -267.525 -1.140 -266.525 ;
        RECT -0.390 -267.525 -0.160 -266.525 ;
        RECT 0.590 -267.525 0.820 -266.525 ;
        RECT 1.160 -267.525 1.390 -266.525 ;
        RECT 2.140 -267.525 2.370 -266.525 ;
        RECT 2.705 -267.525 2.935 -266.525 ;
        RECT 3.685 -267.525 3.915 -266.525 ;
        RECT 11.130 -267.525 11.360 -266.525 ;
        RECT 12.110 -267.525 12.340 -266.525 ;
        RECT 13.090 -267.525 13.320 -266.525 ;
        RECT 13.660 -267.525 13.890 -266.525 ;
        RECT 14.640 -267.525 14.870 -266.525 ;
        RECT 15.205 -267.525 15.435 -266.525 ;
        RECT 16.185 -267.525 16.415 -266.525 ;
        RECT 23.630 -267.525 23.860 -266.525 ;
        RECT 24.610 -267.525 24.840 -266.525 ;
        RECT 25.590 -267.525 25.820 -266.525 ;
        RECT 26.160 -267.525 26.390 -266.525 ;
        RECT 27.140 -267.525 27.370 -266.525 ;
        RECT 27.705 -267.525 27.935 -266.525 ;
        RECT 28.685 -267.525 28.915 -266.525 ;
        RECT 38.630 -267.525 38.860 -266.525 ;
        RECT 39.610 -267.525 39.840 -266.525 ;
        RECT 40.590 -267.525 40.820 -266.525 ;
        RECT 41.160 -267.525 41.390 -266.525 ;
        RECT 42.140 -267.525 42.370 -266.525 ;
        RECT 42.705 -267.525 42.935 -266.525 ;
        RECT 43.685 -267.525 43.915 -266.525 ;
        RECT -139.160 -269.870 -137.160 -269.640 ;
        RECT -106.715 -270.430 -106.485 -269.430 ;
        RECT -105.735 -270.430 -105.505 -269.430 ;
        RECT -104.755 -270.430 -104.525 -269.430 ;
        RECT -103.775 -270.430 -103.545 -269.430 ;
        RECT -101.065 -270.430 -100.835 -269.430 ;
        RECT -100.085 -270.430 -99.855 -269.430 ;
        RECT -139.160 -271.050 -137.160 -270.820 ;
        RECT -96.720 -271.540 -96.490 -270.040 ;
        RECT -95.740 -271.540 -95.510 -270.040 ;
        RECT -94.760 -271.540 -94.530 -270.040 ;
        RECT -93.675 -270.535 -93.445 -270.035 ;
        RECT -92.695 -270.535 -92.465 -270.035 ;
        RECT -91.715 -270.535 -91.485 -270.035 ;
        RECT -90.735 -270.535 -90.505 -270.035 ;
        RECT -19.730 -270.315 -19.115 -269.635 ;
        RECT -139.160 -272.230 -137.160 -272.000 ;
        RECT -68.230 -273.085 -68.000 -272.085 ;
        RECT -67.250 -273.085 -67.020 -272.085 ;
        RECT -66.270 -273.085 -66.040 -272.085 ;
        RECT -59.515 -273.085 -59.285 -272.085 ;
        RECT -58.535 -273.085 -58.305 -272.085 ;
        RECT -57.555 -273.085 -57.325 -272.085 ;
        RECT -54.730 -273.085 -54.500 -272.085 ;
        RECT -53.750 -273.085 -53.520 -272.085 ;
        RECT -52.770 -273.085 -52.540 -272.085 ;
        RECT -46.015 -273.085 -45.785 -272.085 ;
        RECT -45.035 -273.085 -44.805 -272.085 ;
        RECT -44.055 -273.085 -43.825 -272.085 ;
        RECT -41.605 -273.085 -41.375 -272.085 ;
        RECT -40.625 -273.085 -40.395 -272.085 ;
        RECT -39.645 -273.085 -39.415 -272.085 ;
        RECT -139.160 -273.410 -137.160 -273.180 ;
        RECT -139.160 -274.590 -137.160 -274.360 ;
        RECT -139.160 -275.770 -137.160 -275.540 ;
        RECT -88.540 -276.350 -88.310 -274.850 ;
        RECT -87.560 -276.350 -87.330 -274.850 ;
        RECT -86.580 -276.350 -86.350 -274.850 ;
        RECT -85.495 -276.355 -85.265 -275.855 ;
        RECT -84.515 -276.355 -84.285 -275.855 ;
        RECT -83.535 -276.355 -83.305 -275.855 ;
        RECT -82.555 -276.355 -82.325 -275.855 ;
        RECT -139.160 -276.950 -137.160 -276.720 ;
        RECT -81.305 -276.795 -81.075 -273.795 ;
        RECT -80.325 -276.795 -80.095 -273.795 ;
        RECT -78.210 -276.795 -77.980 -273.795 ;
        RECT -28.065 -274.170 -27.835 -273.170 ;
        RECT -27.085 -274.170 -26.855 -273.170 ;
        RECT -26.105 -274.170 -25.875 -273.170 ;
        RECT -19.710 -273.470 -19.140 -270.315 ;
        RECT -6.895 -270.490 -6.280 -269.810 ;
        RECT 5.520 -270.490 6.135 -269.810 ;
        RECT -6.875 -272.750 -6.305 -270.490 ;
        RECT 5.540 -272.575 6.110 -270.490 ;
        RECT 5.515 -272.580 6.130 -272.575 ;
        RECT -6.900 -273.430 -6.285 -272.750 ;
        RECT 5.515 -272.890 7.045 -272.580 ;
        RECT -19.735 -274.150 -19.120 -273.470 ;
        RECT 23.840 -276.785 24.455 -276.740 ;
        RECT 25.845 -276.785 26.460 -276.730 ;
        RECT -0.605 -276.860 0.010 -276.800 ;
        RECT 0.865 -276.860 1.480 -276.795 ;
        RECT -0.605 -277.435 1.480 -276.860 ;
        RECT -0.605 -277.480 0.010 -277.435 ;
        RECT 0.865 -277.475 1.480 -277.435 ;
        RECT 15.755 -276.935 16.370 -276.860 ;
        RECT 17.700 -276.935 18.315 -276.855 ;
        RECT 15.755 -277.470 18.315 -276.935 ;
        RECT 23.840 -277.320 26.460 -276.785 ;
        RECT 23.840 -277.420 24.455 -277.320 ;
        RECT 25.845 -277.410 26.460 -277.320 ;
        RECT 32.625 -276.820 33.240 -276.755 ;
        RECT 38.705 -276.820 39.320 -276.760 ;
        RECT 32.625 -277.345 39.320 -276.820 ;
        RECT 32.625 -277.435 33.240 -277.345 ;
        RECT 38.705 -277.440 39.320 -277.345 ;
        RECT 15.755 -277.540 16.370 -277.470 ;
        RECT 17.700 -277.535 18.315 -277.470 ;
        RECT -139.160 -278.130 -137.160 -277.900 ;
        RECT -139.160 -279.310 -137.160 -279.080 ;
        RECT -139.160 -280.550 -137.160 -280.320 ;
        RECT -106.430 -281.085 -106.200 -279.585 ;
        RECT -105.450 -281.085 -105.220 -279.585 ;
        RECT -104.470 -281.085 -104.240 -279.585 ;
        RECT -103.385 -280.080 -103.155 -279.580 ;
        RECT -102.405 -280.080 -102.175 -279.580 ;
        RECT -101.425 -280.080 -101.195 -279.580 ;
        RECT -100.445 -280.080 -100.215 -279.580 ;
        RECT -97.565 -280.110 -97.335 -279.110 ;
        RECT -96.585 -280.110 -96.355 -279.110 ;
        RECT -95.605 -280.110 -95.375 -279.110 ;
        RECT -94.625 -280.110 -94.395 -279.110 ;
        RECT -91.915 -280.110 -91.685 -279.110 ;
        RECT -90.935 -280.110 -90.705 -279.110 ;
        RECT -88.410 -280.995 -88.180 -279.995 ;
        RECT -87.430 -280.995 -87.200 -279.995 ;
        RECT -86.450 -280.995 -86.220 -279.995 ;
        RECT -85.470 -280.995 -85.240 -279.995 ;
        RECT -83.545 -280.850 -83.315 -279.350 ;
        RECT -82.565 -280.850 -82.335 -279.350 ;
        RECT -81.585 -280.850 -81.355 -279.350 ;
        RECT -80.500 -279.845 -80.270 -279.345 ;
        RECT -79.520 -279.845 -79.290 -279.345 ;
        RECT -78.540 -279.845 -78.310 -279.345 ;
        RECT -77.560 -279.845 -77.330 -279.345 ;
        RECT -63.595 -281.230 -63.365 -279.730 ;
        RECT -62.615 -281.230 -62.385 -279.730 ;
        RECT -61.635 -281.230 -61.405 -279.730 ;
        RECT -60.550 -281.235 -60.320 -280.735 ;
        RECT -59.570 -281.235 -59.340 -280.735 ;
        RECT -58.590 -281.235 -58.360 -280.735 ;
        RECT -57.610 -281.235 -57.380 -280.735 ;
        RECT -139.160 -281.730 -137.160 -281.500 ;
        RECT -56.360 -281.675 -56.130 -278.675 ;
        RECT -55.380 -281.675 -55.150 -278.675 ;
        RECT -53.265 -281.675 -53.035 -278.675 ;
        RECT -28.860 -278.685 -28.630 -277.685 ;
        RECT -27.880 -278.685 -27.650 -277.685 ;
        RECT -26.900 -278.685 -26.670 -277.685 ;
        RECT -20.145 -278.685 -19.915 -277.685 ;
        RECT -19.165 -278.685 -18.935 -277.685 ;
        RECT -18.185 -278.685 -17.955 -277.685 ;
        RECT -15.360 -278.685 -15.130 -277.685 ;
        RECT -14.380 -278.685 -14.150 -277.685 ;
        RECT -13.400 -278.685 -13.170 -277.685 ;
        RECT -6.645 -278.685 -6.415 -277.685 ;
        RECT -5.665 -278.685 -5.435 -277.685 ;
        RECT -4.685 -278.685 -4.455 -277.685 ;
        RECT -2.235 -278.685 -2.005 -277.685 ;
        RECT -1.255 -278.685 -1.025 -277.685 ;
        RECT -0.275 -278.685 -0.045 -277.685 ;
        RECT 1.435 -278.770 1.665 -277.770 ;
        RECT 2.415 -278.770 2.645 -277.770 ;
        RECT 5.125 -278.770 5.355 -277.770 ;
        RECT 6.105 -278.770 6.335 -277.770 ;
        RECT 7.085 -278.770 7.315 -277.770 ;
        RECT 8.065 -278.770 8.295 -277.770 ;
        RECT 10.100 -278.335 10.330 -277.835 ;
        RECT 11.080 -278.335 11.310 -277.835 ;
        RECT 12.060 -278.335 12.290 -277.835 ;
        RECT 13.040 -278.335 13.270 -277.835 ;
        RECT 14.125 -279.340 14.355 -277.840 ;
        RECT 15.105 -279.340 15.335 -277.840 ;
        RECT 16.085 -279.340 16.315 -277.840 ;
        RECT 18.125 -278.345 18.355 -277.845 ;
        RECT 19.105 -278.345 19.335 -277.845 ;
        RECT 20.085 -278.345 20.315 -277.845 ;
        RECT 21.065 -278.345 21.295 -277.845 ;
        RECT 22.150 -279.350 22.380 -277.850 ;
        RECT 23.130 -279.350 23.360 -277.850 ;
        RECT 24.110 -279.350 24.340 -277.850 ;
        RECT 26.245 -278.725 26.475 -277.725 ;
        RECT 27.225 -278.725 27.455 -277.725 ;
        RECT 29.935 -278.725 30.165 -277.725 ;
        RECT 30.915 -278.725 31.145 -277.725 ;
        RECT 31.895 -278.725 32.125 -277.725 ;
        RECT 32.875 -278.725 33.105 -277.725 ;
        RECT 38.680 -278.780 38.910 -277.780 ;
        RECT 39.660 -278.780 39.890 -277.780 ;
        RECT 40.640 -278.780 40.870 -277.780 ;
        RECT 41.210 -278.780 41.440 -277.780 ;
        RECT 42.190 -278.780 42.420 -277.780 ;
        RECT 42.755 -278.780 42.985 -277.780 ;
        RECT 43.735 -278.780 43.965 -277.780 ;
        RECT 141.765 -278.265 141.995 -277.265 ;
        RECT 142.745 -278.265 142.975 -277.265 ;
        RECT 143.725 -278.265 143.955 -277.265 ;
        RECT 144.705 -278.265 144.935 -277.265 ;
        RECT 146.630 -278.910 146.860 -277.410 ;
        RECT 147.610 -278.910 147.840 -277.410 ;
        RECT 148.590 -278.910 148.820 -277.410 ;
        RECT 183.965 -278.320 184.195 -277.320 ;
        RECT 184.945 -278.320 185.175 -277.320 ;
        RECT 185.925 -278.320 186.155 -277.320 ;
        RECT 186.905 -278.320 187.135 -277.320 ;
        RECT 149.675 -278.915 149.905 -278.415 ;
        RECT 150.655 -278.915 150.885 -278.415 ;
        RECT 151.635 -278.915 151.865 -278.415 ;
        RECT 152.615 -278.915 152.845 -278.415 ;
        RECT 188.830 -278.965 189.060 -277.465 ;
        RECT 189.810 -278.965 190.040 -277.465 ;
        RECT 190.790 -278.965 191.020 -277.465 ;
        RECT 191.875 -278.970 192.105 -278.470 ;
        RECT 192.855 -278.970 193.085 -278.470 ;
        RECT 193.835 -278.970 194.065 -278.470 ;
        RECT 194.815 -278.970 195.045 -278.470 ;
        RECT 228.280 -278.515 228.510 -277.515 ;
        RECT 229.260 -278.515 229.490 -277.515 ;
        RECT 230.240 -278.515 230.470 -277.515 ;
        RECT 231.220 -278.515 231.450 -277.515 ;
        RECT 109.905 -280.030 110.135 -279.030 ;
        RECT 110.885 -280.030 111.115 -279.030 ;
        RECT 111.865 -280.030 112.095 -279.030 ;
        RECT 114.090 -280.030 114.320 -279.030 ;
        RECT 115.070 -280.030 115.300 -279.030 ;
        RECT 116.050 -280.030 116.280 -279.030 ;
        RECT 123.405 -280.030 123.635 -279.030 ;
        RECT 124.385 -280.030 124.615 -279.030 ;
        RECT 125.365 -280.030 125.595 -279.030 ;
        RECT 127.590 -280.030 127.820 -279.030 ;
        RECT 128.570 -280.030 128.800 -279.030 ;
        RECT 129.550 -280.030 129.780 -279.030 ;
        RECT 233.145 -279.160 233.375 -277.660 ;
        RECT 234.125 -279.160 234.355 -277.660 ;
        RECT 235.105 -279.160 235.335 -277.660 ;
        RECT 274.270 -278.345 274.500 -277.345 ;
        RECT 275.250 -278.345 275.480 -277.345 ;
        RECT 276.230 -278.345 276.460 -277.345 ;
        RECT 277.210 -278.345 277.440 -277.345 ;
        RECT 236.190 -279.165 236.420 -278.665 ;
        RECT 237.170 -279.165 237.400 -278.665 ;
        RECT 238.150 -279.165 238.380 -278.665 ;
        RECT 239.130 -279.165 239.360 -278.665 ;
        RECT 279.135 -278.990 279.365 -277.490 ;
        RECT 280.115 -278.990 280.345 -277.490 ;
        RECT 281.095 -278.990 281.325 -277.490 ;
        RECT 318.040 -278.015 318.270 -277.015 ;
        RECT 319.020 -278.015 319.250 -277.015 ;
        RECT 320.000 -278.015 320.230 -277.015 ;
        RECT 320.980 -278.015 321.210 -277.015 ;
        RECT 282.180 -278.995 282.410 -278.495 ;
        RECT 283.160 -278.995 283.390 -278.495 ;
        RECT 284.140 -278.995 284.370 -278.495 ;
        RECT 285.120 -278.995 285.350 -278.495 ;
        RECT 322.905 -278.660 323.135 -277.160 ;
        RECT 323.885 -278.660 324.115 -277.160 ;
        RECT 324.865 -278.660 325.095 -277.160 ;
        RECT 363.805 -277.930 364.035 -276.930 ;
        RECT 364.785 -277.930 365.015 -276.930 ;
        RECT 365.765 -277.930 365.995 -276.930 ;
        RECT 366.745 -277.930 366.975 -276.930 ;
        RECT 325.950 -278.665 326.180 -278.165 ;
        RECT 326.930 -278.665 327.160 -278.165 ;
        RECT 327.910 -278.665 328.140 -278.165 ;
        RECT 328.890 -278.665 329.120 -278.165 ;
        RECT 368.670 -278.575 368.900 -277.075 ;
        RECT 369.650 -278.575 369.880 -277.075 ;
        RECT 370.630 -278.575 370.860 -277.075 ;
        RECT 410.625 -277.740 410.855 -276.740 ;
        RECT 411.605 -277.740 411.835 -276.740 ;
        RECT 412.585 -277.740 412.815 -276.740 ;
        RECT 413.565 -277.740 413.795 -276.740 ;
        RECT 371.715 -278.580 371.945 -278.080 ;
        RECT 372.695 -278.580 372.925 -278.080 ;
        RECT 373.675 -278.580 373.905 -278.080 ;
        RECT 374.655 -278.580 374.885 -278.080 ;
        RECT 415.490 -278.385 415.720 -276.885 ;
        RECT 416.470 -278.385 416.700 -276.885 ;
        RECT 417.450 -278.385 417.680 -276.885 ;
        RECT 418.535 -278.390 418.765 -277.890 ;
        RECT 419.515 -278.390 419.745 -277.890 ;
        RECT 420.495 -278.390 420.725 -277.890 ;
        RECT 421.475 -278.390 421.705 -277.890 ;
        RECT 421.885 -279.965 422.255 -279.885 ;
        RECT 423.025 -279.965 423.575 -279.785 ;
        RECT 329.300 -280.240 329.670 -280.160 ;
        RECT 330.440 -280.240 330.990 -280.060 ;
        RECT 153.025 -280.490 153.395 -280.410 ;
        RECT 154.165 -280.490 154.715 -280.310 ;
        RECT 153.025 -280.970 154.715 -280.490 ;
        RECT 195.225 -280.545 195.595 -280.465 ;
        RECT 196.365 -280.545 196.915 -280.365 ;
        RECT 153.025 -281.000 153.395 -280.970 ;
        RECT 154.165 -281.060 154.715 -280.970 ;
        RECT -139.160 -282.910 -137.160 -282.680 ;
        RECT -139.160 -284.090 -137.160 -283.860 ;
        RECT -139.160 -285.270 -137.160 -285.040 ;
        RECT -63.465 -285.875 -63.235 -284.875 ;
        RECT -62.485 -285.875 -62.255 -284.875 ;
        RECT -61.505 -285.875 -61.275 -284.875 ;
        RECT -60.525 -285.875 -60.295 -284.875 ;
        RECT -58.600 -285.730 -58.370 -284.230 ;
        RECT -57.620 -285.730 -57.390 -284.230 ;
        RECT -56.640 -285.730 -56.410 -284.230 ;
        RECT -55.555 -284.725 -55.325 -284.225 ;
        RECT -54.575 -284.725 -54.345 -284.225 ;
        RECT -53.595 -284.725 -53.365 -284.225 ;
        RECT -52.615 -284.725 -52.385 -284.225 ;
        RECT -29.350 -285.275 -29.120 -284.275 ;
        RECT -28.370 -285.275 -28.140 -284.275 ;
        RECT -27.390 -285.275 -27.160 -284.275 ;
        RECT -25.165 -285.275 -24.935 -284.275 ;
        RECT -24.185 -285.275 -23.955 -284.275 ;
        RECT -23.205 -285.275 -22.975 -284.275 ;
        RECT -15.850 -285.275 -15.620 -284.275 ;
        RECT -14.870 -285.275 -14.640 -284.275 ;
        RECT -13.890 -285.275 -13.660 -284.275 ;
        RECT -11.665 -285.275 -11.435 -284.275 ;
        RECT -10.685 -285.275 -10.455 -284.275 ;
        RECT -9.705 -285.275 -9.475 -284.275 ;
        RECT 93.870 -286.020 94.100 -283.020 ;
        RECT 94.850 -286.020 95.080 -283.020 ;
        RECT 141.635 -283.410 141.865 -281.910 ;
        RECT 142.615 -283.410 142.845 -281.910 ;
        RECT 143.595 -283.410 143.825 -281.910 ;
        RECT 144.680 -282.405 144.910 -281.905 ;
        RECT 145.660 -282.405 145.890 -281.905 ;
        RECT 146.640 -282.405 146.870 -281.905 ;
        RECT 147.620 -282.405 147.850 -281.905 ;
        RECT 148.870 -284.465 149.100 -281.465 ;
        RECT 149.850 -284.465 150.080 -281.465 ;
        RECT 151.965 -284.465 152.195 -281.465 ;
        RECT 158.830 -283.255 159.060 -280.755 ;
        RECT 159.810 -283.255 160.040 -280.755 ;
        RECT 162.785 -283.255 163.015 -280.755 ;
        RECT 163.435 -283.255 163.665 -280.755 ;
        RECT 164.575 -282.255 164.805 -280.755 ;
        RECT 165.555 -282.255 165.785 -280.755 ;
        RECT 195.225 -281.025 196.915 -280.545 ;
        RECT 239.540 -280.740 239.910 -280.660 ;
        RECT 240.680 -280.740 241.230 -280.560 ;
        RECT 195.225 -281.055 195.595 -281.025 ;
        RECT 196.365 -281.115 196.915 -281.025 ;
        RECT 183.835 -283.465 184.065 -281.965 ;
        RECT 184.815 -283.465 185.045 -281.965 ;
        RECT 185.795 -283.465 186.025 -281.965 ;
        RECT 186.880 -282.460 187.110 -281.960 ;
        RECT 187.860 -282.460 188.090 -281.960 ;
        RECT 188.840 -282.460 189.070 -281.960 ;
        RECT 189.820 -282.460 190.050 -281.960 ;
        RECT 191.070 -284.520 191.300 -281.520 ;
        RECT 192.050 -284.520 192.280 -281.520 ;
        RECT 194.165 -284.520 194.395 -281.520 ;
        RECT 201.030 -283.310 201.260 -280.810 ;
        RECT 202.010 -283.310 202.240 -280.810 ;
        RECT 204.985 -283.310 205.215 -280.810 ;
        RECT 205.635 -283.310 205.865 -280.810 ;
        RECT 206.775 -282.310 207.005 -280.810 ;
        RECT 207.755 -282.310 207.985 -280.810 ;
        RECT 239.540 -281.220 241.230 -280.740 ;
        RECT 285.530 -280.570 285.900 -280.490 ;
        RECT 286.670 -280.570 287.220 -280.390 ;
        RECT 239.540 -281.250 239.910 -281.220 ;
        RECT 240.680 -281.310 241.230 -281.220 ;
        RECT 228.150 -283.660 228.380 -282.160 ;
        RECT 229.130 -283.660 229.360 -282.160 ;
        RECT 230.110 -283.660 230.340 -282.160 ;
        RECT 231.195 -282.655 231.425 -282.155 ;
        RECT 232.175 -282.655 232.405 -282.155 ;
        RECT 233.155 -282.655 233.385 -282.155 ;
        RECT 234.135 -282.655 234.365 -282.155 ;
        RECT 235.385 -284.715 235.615 -281.715 ;
        RECT 236.365 -284.715 236.595 -281.715 ;
        RECT 238.480 -284.715 238.710 -281.715 ;
        RECT 245.345 -283.505 245.575 -281.005 ;
        RECT 246.325 -283.505 246.555 -281.005 ;
        RECT 249.300 -283.505 249.530 -281.005 ;
        RECT 249.950 -283.505 250.180 -281.005 ;
        RECT 251.090 -282.505 251.320 -281.005 ;
        RECT 252.070 -282.505 252.300 -281.005 ;
        RECT 285.530 -281.050 287.220 -280.570 ;
        RECT 329.300 -280.720 330.990 -280.240 ;
        RECT 375.065 -280.155 375.435 -280.075 ;
        RECT 376.205 -280.155 376.755 -279.975 ;
        RECT 329.300 -280.750 329.670 -280.720 ;
        RECT 330.440 -280.810 330.990 -280.720 ;
        RECT 285.530 -281.080 285.900 -281.050 ;
        RECT 286.670 -281.140 287.220 -281.050 ;
        RECT 274.140 -283.490 274.370 -281.990 ;
        RECT 275.120 -283.490 275.350 -281.990 ;
        RECT 276.100 -283.490 276.330 -281.990 ;
        RECT 277.185 -282.485 277.415 -281.985 ;
        RECT 278.165 -282.485 278.395 -281.985 ;
        RECT 279.145 -282.485 279.375 -281.985 ;
        RECT 280.125 -282.485 280.355 -281.985 ;
        RECT 281.375 -284.545 281.605 -281.545 ;
        RECT 282.355 -284.545 282.585 -281.545 ;
        RECT 284.470 -284.545 284.700 -281.545 ;
        RECT 291.335 -283.335 291.565 -280.835 ;
        RECT 292.315 -283.335 292.545 -280.835 ;
        RECT 295.290 -283.335 295.520 -280.835 ;
        RECT 295.940 -283.335 296.170 -280.835 ;
        RECT 297.080 -282.335 297.310 -280.835 ;
        RECT 298.060 -282.335 298.290 -280.835 ;
        RECT 317.910 -283.160 318.140 -281.660 ;
        RECT 318.890 -283.160 319.120 -281.660 ;
        RECT 319.870 -283.160 320.100 -281.660 ;
        RECT 320.955 -282.155 321.185 -281.655 ;
        RECT 321.935 -282.155 322.165 -281.655 ;
        RECT 322.915 -282.155 323.145 -281.655 ;
        RECT 323.895 -282.155 324.125 -281.655 ;
        RECT 325.145 -284.215 325.375 -281.215 ;
        RECT 326.125 -284.215 326.355 -281.215 ;
        RECT 328.240 -284.215 328.470 -281.215 ;
        RECT 335.105 -283.005 335.335 -280.505 ;
        RECT 336.085 -283.005 336.315 -280.505 ;
        RECT 339.060 -283.005 339.290 -280.505 ;
        RECT 339.710 -283.005 339.940 -280.505 ;
        RECT 340.850 -282.005 341.080 -280.505 ;
        RECT 341.830 -282.005 342.060 -280.505 ;
        RECT 375.065 -280.635 376.755 -280.155 ;
        RECT 375.065 -280.665 375.435 -280.635 ;
        RECT 376.205 -280.725 376.755 -280.635 ;
        RECT 363.675 -283.075 363.905 -281.575 ;
        RECT 364.655 -283.075 364.885 -281.575 ;
        RECT 365.635 -283.075 365.865 -281.575 ;
        RECT 366.720 -282.070 366.950 -281.570 ;
        RECT 367.700 -282.070 367.930 -281.570 ;
        RECT 368.680 -282.070 368.910 -281.570 ;
        RECT 369.660 -282.070 369.890 -281.570 ;
        RECT 370.910 -284.130 371.140 -281.130 ;
        RECT 371.890 -284.130 372.120 -281.130 ;
        RECT 374.005 -284.130 374.235 -281.130 ;
        RECT 380.870 -282.920 381.100 -280.420 ;
        RECT 381.850 -282.920 382.080 -280.420 ;
        RECT 384.825 -282.920 385.055 -280.420 ;
        RECT 385.475 -282.920 385.705 -280.420 ;
        RECT 386.615 -281.920 386.845 -280.420 ;
        RECT 387.595 -281.920 387.825 -280.420 ;
        RECT 421.885 -280.445 423.575 -279.965 ;
        RECT 421.885 -280.475 422.255 -280.445 ;
        RECT 423.025 -280.535 423.575 -280.445 ;
        RECT 410.495 -282.885 410.725 -281.385 ;
        RECT 411.475 -282.885 411.705 -281.385 ;
        RECT 412.455 -282.885 412.685 -281.385 ;
        RECT 413.540 -281.880 413.770 -281.380 ;
        RECT 414.520 -281.880 414.750 -281.380 ;
        RECT 415.500 -281.880 415.730 -281.380 ;
        RECT 416.480 -281.880 416.710 -281.380 ;
        RECT 417.730 -283.940 417.960 -280.940 ;
        RECT 418.710 -283.940 418.940 -280.940 ;
        RECT 420.825 -283.940 421.055 -280.940 ;
        RECT 427.690 -282.730 427.920 -280.230 ;
        RECT 428.670 -282.730 428.900 -280.230 ;
        RECT 431.645 -282.730 431.875 -280.230 ;
        RECT 432.295 -282.730 432.525 -280.230 ;
        RECT 433.435 -281.730 433.665 -280.230 ;
        RECT 434.415 -281.730 434.645 -280.230 ;
        RECT -139.160 -286.450 -137.160 -286.220 ;
        RECT 100.475 -286.620 100.705 -285.620 ;
        RECT 101.455 -286.620 101.685 -285.620 ;
        RECT 102.435 -286.620 102.665 -285.620 ;
        RECT 104.885 -286.620 105.115 -285.620 ;
        RECT 105.865 -286.620 106.095 -285.620 ;
        RECT 106.845 -286.620 107.075 -285.620 ;
        RECT 113.600 -286.620 113.830 -285.620 ;
        RECT 114.580 -286.620 114.810 -285.620 ;
        RECT 115.560 -286.620 115.790 -285.620 ;
        RECT 118.385 -286.620 118.615 -285.620 ;
        RECT 119.365 -286.620 119.595 -285.620 ;
        RECT 120.345 -286.620 120.575 -285.620 ;
        RECT 127.100 -286.620 127.330 -285.620 ;
        RECT 128.080 -286.620 128.310 -285.620 ;
        RECT 129.060 -286.620 129.290 -285.620 ;
        RECT -139.160 -287.630 -137.160 -287.400 ;
        RECT -139.160 -288.810 -137.160 -288.580 ;
        RECT -139.160 -289.990 -137.160 -289.760 ;
        RECT -139.160 -290.640 -137.160 -290.410 ;
        RECT -68.720 -291.130 -68.490 -290.130 ;
        RECT -67.740 -291.130 -67.510 -290.130 ;
        RECT -66.760 -291.130 -66.530 -290.130 ;
        RECT -64.535 -291.130 -64.305 -290.130 ;
        RECT -63.555 -291.130 -63.325 -290.130 ;
        RECT -62.575 -291.130 -62.345 -290.130 ;
        RECT -55.220 -291.130 -54.990 -290.130 ;
        RECT -54.240 -291.130 -54.010 -290.130 ;
        RECT -53.260 -291.130 -53.030 -290.130 ;
        RECT -51.035 -291.130 -50.805 -290.130 ;
        RECT -50.055 -291.130 -49.825 -290.130 ;
        RECT -49.075 -291.130 -48.845 -290.130 ;
        RECT -139.160 -291.820 -137.160 -291.590 ;
        RECT -139.160 -293.000 -137.160 -292.770 ;
        RECT -90.845 -293.655 -89.950 -292.820 ;
        RECT -36.775 -293.215 -36.545 -290.215 ;
        RECT -34.660 -293.215 -34.430 -290.215 ;
        RECT -33.680 -293.215 -33.450 -290.215 ;
        RECT 112.700 -291.380 112.930 -289.380 ;
        RECT 113.680 -291.380 113.910 -289.380 ;
        RECT 114.660 -291.380 114.890 -289.380 ;
        RECT -29.350 -292.465 -29.120 -291.465 ;
        RECT -28.370 -292.465 -28.140 -291.465 ;
        RECT -27.390 -292.465 -27.160 -291.465 ;
        RECT -25.165 -292.465 -24.935 -291.465 ;
        RECT -24.185 -292.465 -23.955 -291.465 ;
        RECT -23.205 -292.465 -22.975 -291.465 ;
        RECT -15.850 -292.465 -15.620 -291.465 ;
        RECT -14.870 -292.465 -14.640 -291.465 ;
        RECT -13.890 -292.465 -13.660 -291.465 ;
        RECT -11.665 -292.465 -11.435 -291.465 ;
        RECT -10.685 -292.465 -10.455 -291.465 ;
        RECT -9.705 -292.465 -9.475 -291.465 ;
        RECT -139.160 -294.180 -137.160 -293.950 ;
        RECT -139.160 -295.360 -137.160 -295.130 ;
        RECT -139.160 -296.010 -137.160 -295.780 ;
        RECT -139.160 -297.190 -137.160 -296.960 ;
        RECT -139.160 -298.370 -137.160 -298.140 ;
        RECT -106.105 -298.555 -105.875 -295.555 ;
        RECT -105.125 -298.555 -104.895 -295.555 ;
        RECT -100.075 -297.200 -99.845 -295.200 ;
        RECT -99.095 -297.200 -98.865 -295.200 ;
        RECT -95.550 -297.205 -95.320 -295.205 ;
        RECT -94.570 -297.205 -94.340 -295.205 ;
        RECT -90.710 -302.475 -90.080 -293.655 ;
        RECT -68.230 -297.720 -68.000 -296.720 ;
        RECT -67.250 -297.720 -67.020 -296.720 ;
        RECT -66.270 -297.720 -66.040 -296.720 ;
        RECT -59.515 -297.720 -59.285 -296.720 ;
        RECT -58.535 -297.720 -58.305 -296.720 ;
        RECT -57.555 -297.720 -57.325 -296.720 ;
        RECT -54.730 -297.720 -54.500 -296.720 ;
        RECT -53.750 -297.720 -53.520 -296.720 ;
        RECT -52.770 -297.720 -52.540 -296.720 ;
        RECT -46.015 -297.720 -45.785 -296.720 ;
        RECT -45.035 -297.720 -44.805 -296.720 ;
        RECT -44.055 -297.720 -43.825 -296.720 ;
        RECT -41.605 -297.720 -41.375 -296.720 ;
        RECT -40.625 -297.720 -40.395 -296.720 ;
        RECT -39.645 -297.720 -39.415 -296.720 ;
        RECT -88.540 -301.350 -88.310 -299.850 ;
        RECT -87.560 -301.350 -87.330 -299.850 ;
        RECT -86.580 -301.350 -86.350 -299.850 ;
        RECT -85.495 -301.355 -85.265 -300.855 ;
        RECT -84.515 -301.355 -84.285 -300.855 ;
        RECT -83.535 -301.355 -83.305 -300.855 ;
        RECT -82.555 -301.355 -82.325 -300.855 ;
        RECT -81.305 -301.795 -81.075 -298.795 ;
        RECT -80.325 -301.795 -80.095 -298.795 ;
        RECT -78.210 -301.795 -77.980 -298.795 ;
        RECT -28.860 -299.055 -28.630 -298.055 ;
        RECT -27.880 -299.055 -27.650 -298.055 ;
        RECT -26.900 -299.055 -26.670 -298.055 ;
        RECT -20.145 -299.055 -19.915 -298.055 ;
        RECT -19.165 -299.055 -18.935 -298.055 ;
        RECT -18.185 -299.055 -17.955 -298.055 ;
        RECT -15.360 -299.055 -15.130 -298.055 ;
        RECT -14.380 -299.055 -14.150 -298.055 ;
        RECT -13.400 -299.055 -13.170 -298.055 ;
        RECT -6.645 -299.055 -6.415 -298.055 ;
        RECT -5.665 -299.055 -5.435 -298.055 ;
        RECT -4.685 -299.055 -4.455 -298.055 ;
        RECT -2.235 -299.055 -2.005 -298.055 ;
        RECT -1.255 -299.055 -1.025 -298.055 ;
        RECT -0.275 -299.055 -0.045 -298.055 ;
        RECT 1.435 -298.970 1.665 -297.970 ;
        RECT 2.415 -298.970 2.645 -297.970 ;
        RECT 5.125 -298.970 5.355 -297.970 ;
        RECT 6.105 -298.970 6.335 -297.970 ;
        RECT 7.085 -298.970 7.315 -297.970 ;
        RECT 8.065 -298.970 8.295 -297.970 ;
        RECT 10.100 -298.905 10.330 -298.405 ;
        RECT 11.080 -298.905 11.310 -298.405 ;
        RECT 12.060 -298.905 12.290 -298.405 ;
        RECT 13.040 -298.905 13.270 -298.405 ;
        RECT 14.125 -298.900 14.355 -297.400 ;
        RECT 15.105 -298.900 15.335 -297.400 ;
        RECT 16.085 -298.900 16.315 -297.400 ;
        RECT 18.125 -298.895 18.355 -298.395 ;
        RECT 19.105 -298.895 19.335 -298.395 ;
        RECT 20.085 -298.895 20.315 -298.395 ;
        RECT 21.065 -298.895 21.295 -298.395 ;
        RECT 22.150 -298.890 22.380 -297.390 ;
        RECT 23.130 -298.890 23.360 -297.390 ;
        RECT 24.110 -298.890 24.340 -297.390 ;
        RECT 93.845 -297.750 94.075 -295.750 ;
        RECT 94.825 -297.750 95.055 -295.750 ;
        RECT 98.575 -297.750 98.805 -295.750 ;
        RECT 99.555 -297.750 99.785 -295.750 ;
        RECT 103.155 -297.920 103.385 -296.920 ;
        RECT 104.135 -297.920 104.365 -296.920 ;
        RECT 105.115 -297.920 105.345 -296.920 ;
        RECT 106.095 -297.920 106.325 -296.920 ;
        RECT 108.805 -297.920 109.035 -296.920 ;
        RECT 109.785 -297.920 110.015 -296.920 ;
        RECT 112.450 -297.885 112.680 -296.885 ;
        RECT 113.430 -297.885 113.660 -296.885 ;
        RECT 114.410 -297.885 114.640 -296.885 ;
        RECT 116.850 -297.530 117.080 -294.030 ;
        RECT 117.830 -297.530 118.060 -294.030 ;
        RECT 118.850 -297.530 119.080 -294.030 ;
        RECT 119.830 -297.530 120.060 -294.030 ;
        RECT 121.850 -297.530 122.080 -294.030 ;
        RECT 122.830 -297.530 123.060 -294.030 ;
        RECT 123.850 -297.530 124.080 -294.030 ;
        RECT 124.830 -297.530 125.060 -294.030 ;
        RECT 126.850 -297.530 127.080 -294.030 ;
        RECT 127.830 -297.530 128.060 -294.030 ;
        RECT 128.850 -297.530 129.080 -294.030 ;
        RECT 129.830 -297.530 130.060 -294.030 ;
        RECT 141.725 -295.530 141.955 -294.530 ;
        RECT 142.705 -295.530 142.935 -294.530 ;
        RECT 143.685 -295.530 143.915 -294.530 ;
        RECT 144.665 -295.530 144.895 -294.530 ;
        RECT 146.590 -296.175 146.820 -294.675 ;
        RECT 147.570 -296.175 147.800 -294.675 ;
        RECT 148.550 -296.175 148.780 -294.675 ;
        RECT 149.635 -296.180 149.865 -295.680 ;
        RECT 150.615 -296.180 150.845 -295.680 ;
        RECT 151.595 -296.180 151.825 -295.680 ;
        RECT 152.575 -296.180 152.805 -295.680 ;
        RECT 160.065 -295.685 160.295 -294.685 ;
        RECT 161.045 -295.685 161.275 -294.685 ;
        RECT 162.025 -295.685 162.255 -294.685 ;
        RECT 163.005 -295.685 163.235 -294.685 ;
        RECT 164.930 -296.330 165.160 -294.830 ;
        RECT 165.910 -296.330 166.140 -294.830 ;
        RECT 166.890 -296.330 167.120 -294.830 ;
        RECT 183.925 -295.585 184.155 -294.585 ;
        RECT 184.905 -295.585 185.135 -294.585 ;
        RECT 185.885 -295.585 186.115 -294.585 ;
        RECT 186.865 -295.585 187.095 -294.585 ;
        RECT 167.975 -296.335 168.205 -295.835 ;
        RECT 168.955 -296.335 169.185 -295.835 ;
        RECT 169.935 -296.335 170.165 -295.835 ;
        RECT 170.915 -296.335 171.145 -295.835 ;
        RECT 188.790 -296.230 189.020 -294.730 ;
        RECT 189.770 -296.230 190.000 -294.730 ;
        RECT 190.750 -296.230 190.980 -294.730 ;
        RECT 191.835 -296.235 192.065 -295.735 ;
        RECT 192.815 -296.235 193.045 -295.735 ;
        RECT 193.795 -296.235 194.025 -295.735 ;
        RECT 194.775 -296.235 195.005 -295.735 ;
        RECT 202.265 -295.740 202.495 -294.740 ;
        RECT 203.245 -295.740 203.475 -294.740 ;
        RECT 204.225 -295.740 204.455 -294.740 ;
        RECT 205.205 -295.740 205.435 -294.740 ;
        RECT 207.130 -296.385 207.360 -294.885 ;
        RECT 208.110 -296.385 208.340 -294.885 ;
        RECT 209.090 -296.385 209.320 -294.885 ;
        RECT 228.240 -295.780 228.470 -294.780 ;
        RECT 229.220 -295.780 229.450 -294.780 ;
        RECT 230.200 -295.780 230.430 -294.780 ;
        RECT 231.180 -295.780 231.410 -294.780 ;
        RECT 210.175 -296.390 210.405 -295.890 ;
        RECT 211.155 -296.390 211.385 -295.890 ;
        RECT 212.135 -296.390 212.365 -295.890 ;
        RECT 213.115 -296.390 213.345 -295.890 ;
        RECT 233.105 -296.425 233.335 -294.925 ;
        RECT 234.085 -296.425 234.315 -294.925 ;
        RECT 235.065 -296.425 235.295 -294.925 ;
        RECT 236.150 -296.430 236.380 -295.930 ;
        RECT 237.130 -296.430 237.360 -295.930 ;
        RECT 238.110 -296.430 238.340 -295.930 ;
        RECT 239.090 -296.430 239.320 -295.930 ;
        RECT 246.580 -295.935 246.810 -294.935 ;
        RECT 247.560 -295.935 247.790 -294.935 ;
        RECT 248.540 -295.935 248.770 -294.935 ;
        RECT 249.520 -295.935 249.750 -294.935 ;
        RECT 251.445 -296.580 251.675 -295.080 ;
        RECT 252.425 -296.580 252.655 -295.080 ;
        RECT 253.405 -296.580 253.635 -295.080 ;
        RECT 274.230 -295.610 274.460 -294.610 ;
        RECT 275.210 -295.610 275.440 -294.610 ;
        RECT 276.190 -295.610 276.420 -294.610 ;
        RECT 277.170 -295.610 277.400 -294.610 ;
        RECT 254.490 -296.585 254.720 -296.085 ;
        RECT 255.470 -296.585 255.700 -296.085 ;
        RECT 256.450 -296.585 256.680 -296.085 ;
        RECT 257.430 -296.585 257.660 -296.085 ;
        RECT 279.095 -296.255 279.325 -294.755 ;
        RECT 280.075 -296.255 280.305 -294.755 ;
        RECT 281.055 -296.255 281.285 -294.755 ;
        RECT 282.140 -296.260 282.370 -295.760 ;
        RECT 283.120 -296.260 283.350 -295.760 ;
        RECT 284.100 -296.260 284.330 -295.760 ;
        RECT 285.080 -296.260 285.310 -295.760 ;
        RECT 292.570 -295.765 292.800 -294.765 ;
        RECT 293.550 -295.765 293.780 -294.765 ;
        RECT 294.530 -295.765 294.760 -294.765 ;
        RECT 295.510 -295.765 295.740 -294.765 ;
        RECT 297.435 -296.410 297.665 -294.910 ;
        RECT 298.415 -296.410 298.645 -294.910 ;
        RECT 299.395 -296.410 299.625 -294.910 ;
        RECT 318.000 -295.280 318.230 -294.280 ;
        RECT 318.980 -295.280 319.210 -294.280 ;
        RECT 319.960 -295.280 320.190 -294.280 ;
        RECT 320.940 -295.280 321.170 -294.280 ;
        RECT 300.480 -296.415 300.710 -295.915 ;
        RECT 301.460 -296.415 301.690 -295.915 ;
        RECT 302.440 -296.415 302.670 -295.915 ;
        RECT 303.420 -296.415 303.650 -295.915 ;
        RECT 322.865 -295.925 323.095 -294.425 ;
        RECT 323.845 -295.925 324.075 -294.425 ;
        RECT 324.825 -295.925 325.055 -294.425 ;
        RECT 325.910 -295.930 326.140 -295.430 ;
        RECT 326.890 -295.930 327.120 -295.430 ;
        RECT 327.870 -295.930 328.100 -295.430 ;
        RECT 328.850 -295.930 329.080 -295.430 ;
        RECT 336.340 -295.435 336.570 -294.435 ;
        RECT 337.320 -295.435 337.550 -294.435 ;
        RECT 338.300 -295.435 338.530 -294.435 ;
        RECT 339.280 -295.435 339.510 -294.435 ;
        RECT 341.205 -296.080 341.435 -294.580 ;
        RECT 342.185 -296.080 342.415 -294.580 ;
        RECT 343.165 -296.080 343.395 -294.580 ;
        RECT 363.765 -295.195 363.995 -294.195 ;
        RECT 364.745 -295.195 364.975 -294.195 ;
        RECT 365.725 -295.195 365.955 -294.195 ;
        RECT 366.705 -295.195 366.935 -294.195 ;
        RECT 344.250 -296.085 344.480 -295.585 ;
        RECT 345.230 -296.085 345.460 -295.585 ;
        RECT 346.210 -296.085 346.440 -295.585 ;
        RECT 347.190 -296.085 347.420 -295.585 ;
        RECT 368.630 -295.840 368.860 -294.340 ;
        RECT 369.610 -295.840 369.840 -294.340 ;
        RECT 370.590 -295.840 370.820 -294.340 ;
        RECT 371.675 -295.845 371.905 -295.345 ;
        RECT 372.655 -295.845 372.885 -295.345 ;
        RECT 373.635 -295.845 373.865 -295.345 ;
        RECT 374.615 -295.845 374.845 -295.345 ;
        RECT 382.105 -295.350 382.335 -294.350 ;
        RECT 383.085 -295.350 383.315 -294.350 ;
        RECT 384.065 -295.350 384.295 -294.350 ;
        RECT 385.045 -295.350 385.275 -294.350 ;
        RECT 386.970 -295.995 387.200 -294.495 ;
        RECT 387.950 -295.995 388.180 -294.495 ;
        RECT 388.930 -295.995 389.160 -294.495 ;
        RECT 410.585 -295.005 410.815 -294.005 ;
        RECT 411.565 -295.005 411.795 -294.005 ;
        RECT 412.545 -295.005 412.775 -294.005 ;
        RECT 413.525 -295.005 413.755 -294.005 ;
        RECT 390.015 -296.000 390.245 -295.500 ;
        RECT 390.995 -296.000 391.225 -295.500 ;
        RECT 391.975 -296.000 392.205 -295.500 ;
        RECT 392.955 -296.000 393.185 -295.500 ;
        RECT 415.450 -295.650 415.680 -294.150 ;
        RECT 416.430 -295.650 416.660 -294.150 ;
        RECT 417.410 -295.650 417.640 -294.150 ;
        RECT 418.495 -295.655 418.725 -295.155 ;
        RECT 419.475 -295.655 419.705 -295.155 ;
        RECT 420.455 -295.655 420.685 -295.155 ;
        RECT 421.435 -295.655 421.665 -295.155 ;
        RECT 428.925 -295.160 429.155 -294.160 ;
        RECT 429.905 -295.160 430.135 -294.160 ;
        RECT 430.885 -295.160 431.115 -294.160 ;
        RECT 431.865 -295.160 432.095 -294.160 ;
        RECT 433.790 -295.805 434.020 -294.305 ;
        RECT 434.770 -295.805 435.000 -294.305 ;
        RECT 435.750 -295.805 435.980 -294.305 ;
        RECT 436.835 -295.810 437.065 -295.310 ;
        RECT 437.815 -295.810 438.045 -295.310 ;
        RECT 438.795 -295.810 439.025 -295.310 ;
        RECT 439.775 -295.810 440.005 -295.310 ;
        RECT 323.875 -297.300 324.790 -297.095 ;
        RECT 330.390 -297.300 330.870 -297.155 ;
        RECT 369.640 -297.215 370.555 -297.010 ;
        RECT 416.460 -297.025 417.375 -296.820 ;
        RECT 422.975 -297.025 423.455 -296.880 ;
        RECT 376.155 -297.215 376.635 -297.070 ;
        RECT 147.600 -297.550 148.515 -297.345 ;
        RECT 154.115 -297.550 154.595 -297.405 ;
        RECT 147.600 -297.960 154.595 -297.550 ;
        RECT 26.245 -299.015 26.475 -298.015 ;
        RECT 27.225 -299.015 27.455 -298.015 ;
        RECT 29.935 -299.015 30.165 -298.015 ;
        RECT 30.915 -299.015 31.145 -298.015 ;
        RECT 31.895 -299.015 32.125 -298.015 ;
        RECT 32.875 -299.015 33.105 -298.015 ;
        RECT 38.680 -298.960 38.910 -297.960 ;
        RECT 39.660 -298.960 39.890 -297.960 ;
        RECT 40.640 -298.960 40.870 -297.960 ;
        RECT 41.210 -298.960 41.440 -297.960 ;
        RECT 42.190 -298.960 42.420 -297.960 ;
        RECT 42.755 -298.960 42.985 -297.960 ;
        RECT 43.735 -298.960 43.965 -297.960 ;
        RECT 147.600 -297.995 148.515 -297.960 ;
        RECT 154.115 -298.090 154.595 -297.960 ;
        RECT 171.215 -297.660 171.670 -297.600 ;
        RECT 172.465 -297.660 173.220 -297.525 ;
        RECT 171.215 -298.355 173.220 -297.660 ;
        RECT 189.800 -297.605 190.715 -297.400 ;
        RECT 196.315 -297.605 196.795 -297.460 ;
        RECT 189.800 -298.015 196.795 -297.605 ;
        RECT 189.800 -298.050 190.715 -298.015 ;
        RECT 196.315 -298.145 196.795 -298.015 ;
        RECT 213.415 -297.715 213.870 -297.655 ;
        RECT 214.665 -297.715 215.420 -297.580 ;
        RECT 171.215 -298.415 171.670 -298.355 ;
        RECT 172.465 -298.480 173.220 -298.355 ;
        RECT 213.415 -298.410 215.420 -297.715 ;
        RECT 234.115 -297.800 235.030 -297.595 ;
        RECT 280.105 -297.630 281.020 -297.425 ;
        RECT 286.620 -297.630 287.100 -297.485 ;
        RECT 240.630 -297.800 241.110 -297.655 ;
        RECT 234.115 -298.210 241.110 -297.800 ;
        RECT 234.115 -298.245 235.030 -298.210 ;
        RECT 240.630 -298.340 241.110 -298.210 ;
        RECT 257.730 -297.910 258.185 -297.850 ;
        RECT 258.980 -297.910 259.735 -297.775 ;
        RECT 213.415 -298.470 213.870 -298.410 ;
        RECT 214.665 -298.535 215.420 -298.410 ;
        RECT 257.730 -298.605 259.735 -297.910 ;
        RECT 280.105 -298.040 287.100 -297.630 ;
        RECT 280.105 -298.075 281.020 -298.040 ;
        RECT 286.620 -298.170 287.100 -298.040 ;
        RECT 303.720 -297.740 304.175 -297.680 ;
        RECT 304.970 -297.740 305.725 -297.605 ;
        RECT 303.720 -298.435 305.725 -297.740 ;
        RECT 323.875 -297.710 330.870 -297.300 ;
        RECT 323.875 -297.745 324.790 -297.710 ;
        RECT 330.390 -297.840 330.870 -297.710 ;
        RECT 347.490 -297.410 347.945 -297.350 ;
        RECT 348.740 -297.410 349.495 -297.275 ;
        RECT 347.490 -298.105 349.495 -297.410 ;
        RECT 369.640 -297.625 376.635 -297.215 ;
        RECT 369.640 -297.660 370.555 -297.625 ;
        RECT 376.155 -297.755 376.635 -297.625 ;
        RECT 393.255 -297.325 393.710 -297.265 ;
        RECT 394.505 -297.325 395.260 -297.190 ;
        RECT 393.255 -298.020 395.260 -297.325 ;
        RECT 416.460 -297.435 423.455 -297.025 ;
        RECT 416.460 -297.470 417.375 -297.435 ;
        RECT 422.975 -297.565 423.455 -297.435 ;
        RECT 440.075 -297.135 440.530 -297.075 ;
        RECT 441.325 -297.135 442.080 -297.000 ;
        RECT 440.075 -297.830 442.080 -297.135 ;
        RECT 440.075 -297.890 440.530 -297.830 ;
        RECT 441.325 -297.955 442.080 -297.830 ;
        RECT 393.255 -298.080 393.710 -298.020 ;
        RECT 347.490 -298.165 347.945 -298.105 ;
        RECT 348.740 -298.230 349.495 -298.105 ;
        RECT 394.505 -298.145 395.260 -298.020 ;
        RECT 303.720 -298.495 304.175 -298.435 ;
        RECT 304.970 -298.560 305.725 -298.435 ;
        RECT 257.730 -298.665 258.185 -298.605 ;
        RECT 258.980 -298.730 259.735 -298.605 ;
        RECT -0.605 -299.305 0.010 -299.260 ;
        RECT 0.865 -299.305 1.480 -299.265 ;
        RECT -0.605 -299.880 1.480 -299.305 ;
        RECT 15.755 -299.270 16.370 -299.200 ;
        RECT 17.700 -299.270 18.315 -299.205 ;
        RECT 15.755 -299.805 18.315 -299.270 ;
        RECT 15.755 -299.880 16.370 -299.805 ;
        RECT -0.605 -299.940 0.010 -299.880 ;
        RECT 0.865 -299.945 1.480 -299.880 ;
        RECT 17.700 -299.885 18.315 -299.805 ;
        RECT 23.840 -299.420 24.455 -299.320 ;
        RECT 25.845 -299.420 26.460 -299.330 ;
        RECT 23.840 -299.955 26.460 -299.420 ;
        RECT 23.840 -300.000 24.455 -299.955 ;
        RECT 25.845 -300.010 26.460 -299.955 ;
        RECT 32.625 -299.395 33.240 -299.305 ;
        RECT 38.705 -299.395 39.320 -299.300 ;
        RECT 32.625 -299.920 39.320 -299.395 ;
        RECT 32.625 -299.985 33.240 -299.920 ;
        RECT 38.705 -299.980 39.320 -299.920 ;
        RECT 141.595 -300.675 141.825 -299.175 ;
        RECT 142.575 -300.675 142.805 -299.175 ;
        RECT 143.555 -300.675 143.785 -299.175 ;
        RECT 144.640 -299.670 144.870 -299.170 ;
        RECT 145.620 -299.670 145.850 -299.170 ;
        RECT 146.600 -299.670 146.830 -299.170 ;
        RECT 147.580 -299.670 147.810 -299.170 ;
        RECT 148.830 -301.730 149.060 -298.730 ;
        RECT 149.810 -301.730 150.040 -298.730 ;
        RECT 151.925 -301.730 152.155 -298.730 ;
        RECT 159.935 -300.830 160.165 -299.330 ;
        RECT 160.915 -300.830 161.145 -299.330 ;
        RECT 161.895 -300.830 162.125 -299.330 ;
        RECT 162.980 -299.825 163.210 -299.325 ;
        RECT 163.960 -299.825 164.190 -299.325 ;
        RECT 164.940 -299.825 165.170 -299.325 ;
        RECT 165.920 -299.825 166.150 -299.325 ;
        RECT -90.715 -303.335 -89.755 -302.475 ;
        RECT -19.735 -303.270 -19.120 -302.590 ;
        RECT 59.835 -302.810 60.065 -301.810 ;
        RECT 60.815 -302.810 61.045 -301.810 ;
        RECT 61.795 -302.810 62.025 -301.810 ;
        RECT 64.245 -302.810 64.475 -301.810 ;
        RECT 65.225 -302.810 65.455 -301.810 ;
        RECT 66.205 -302.810 66.435 -301.810 ;
        RECT 72.960 -302.810 73.190 -301.810 ;
        RECT 73.940 -302.810 74.170 -301.810 ;
        RECT 74.920 -302.810 75.150 -301.810 ;
        RECT 77.745 -302.810 77.975 -301.810 ;
        RECT 78.725 -302.810 78.955 -301.810 ;
        RECT 79.705 -302.810 79.935 -301.810 ;
        RECT 86.460 -302.810 86.690 -301.810 ;
        RECT 87.440 -302.810 87.670 -301.810 ;
        RECT 88.420 -302.810 88.650 -301.810 ;
        RECT 167.170 -301.885 167.400 -298.885 ;
        RECT 168.150 -301.885 168.380 -298.885 ;
        RECT 170.265 -301.885 170.495 -298.885 ;
        RECT 183.795 -300.730 184.025 -299.230 ;
        RECT 184.775 -300.730 185.005 -299.230 ;
        RECT 185.755 -300.730 185.985 -299.230 ;
        RECT 186.840 -299.725 187.070 -299.225 ;
        RECT 187.820 -299.725 188.050 -299.225 ;
        RECT 188.800 -299.725 189.030 -299.225 ;
        RECT 189.780 -299.725 190.010 -299.225 ;
        RECT 191.030 -301.785 191.260 -298.785 ;
        RECT 192.010 -301.785 192.240 -298.785 ;
        RECT 194.125 -301.785 194.355 -298.785 ;
        RECT 202.135 -300.885 202.365 -299.385 ;
        RECT 203.115 -300.885 203.345 -299.385 ;
        RECT 204.095 -300.885 204.325 -299.385 ;
        RECT 205.180 -299.880 205.410 -299.380 ;
        RECT 206.160 -299.880 206.390 -299.380 ;
        RECT 207.140 -299.880 207.370 -299.380 ;
        RECT 208.120 -299.880 208.350 -299.380 ;
        RECT 209.370 -301.940 209.600 -298.940 ;
        RECT 210.350 -301.940 210.580 -298.940 ;
        RECT 212.465 -301.940 212.695 -298.940 ;
        RECT 228.110 -300.925 228.340 -299.425 ;
        RECT 229.090 -300.925 229.320 -299.425 ;
        RECT 230.070 -300.925 230.300 -299.425 ;
        RECT 231.155 -299.920 231.385 -299.420 ;
        RECT 232.135 -299.920 232.365 -299.420 ;
        RECT 233.115 -299.920 233.345 -299.420 ;
        RECT 234.095 -299.920 234.325 -299.420 ;
        RECT 235.345 -301.980 235.575 -298.980 ;
        RECT 236.325 -301.980 236.555 -298.980 ;
        RECT 238.440 -301.980 238.670 -298.980 ;
        RECT 246.450 -301.080 246.680 -299.580 ;
        RECT 247.430 -301.080 247.660 -299.580 ;
        RECT 248.410 -301.080 248.640 -299.580 ;
        RECT 249.495 -300.075 249.725 -299.575 ;
        RECT 250.475 -300.075 250.705 -299.575 ;
        RECT 251.455 -300.075 251.685 -299.575 ;
        RECT 252.435 -300.075 252.665 -299.575 ;
        RECT 253.685 -302.135 253.915 -299.135 ;
        RECT 254.665 -302.135 254.895 -299.135 ;
        RECT 256.780 -302.135 257.010 -299.135 ;
        RECT 274.100 -300.755 274.330 -299.255 ;
        RECT 275.080 -300.755 275.310 -299.255 ;
        RECT 276.060 -300.755 276.290 -299.255 ;
        RECT 277.145 -299.750 277.375 -299.250 ;
        RECT 278.125 -299.750 278.355 -299.250 ;
        RECT 279.105 -299.750 279.335 -299.250 ;
        RECT 280.085 -299.750 280.315 -299.250 ;
        RECT 281.335 -301.810 281.565 -298.810 ;
        RECT 282.315 -301.810 282.545 -298.810 ;
        RECT 284.430 -301.810 284.660 -298.810 ;
        RECT 292.440 -300.910 292.670 -299.410 ;
        RECT 293.420 -300.910 293.650 -299.410 ;
        RECT 294.400 -300.910 294.630 -299.410 ;
        RECT 295.485 -299.905 295.715 -299.405 ;
        RECT 296.465 -299.905 296.695 -299.405 ;
        RECT 297.445 -299.905 297.675 -299.405 ;
        RECT 298.425 -299.905 298.655 -299.405 ;
        RECT 299.675 -301.965 299.905 -298.965 ;
        RECT 300.655 -301.965 300.885 -298.965 ;
        RECT 302.770 -301.965 303.000 -298.965 ;
        RECT 317.870 -300.425 318.100 -298.925 ;
        RECT 318.850 -300.425 319.080 -298.925 ;
        RECT 319.830 -300.425 320.060 -298.925 ;
        RECT 320.915 -299.420 321.145 -298.920 ;
        RECT 321.895 -299.420 322.125 -298.920 ;
        RECT 322.875 -299.420 323.105 -298.920 ;
        RECT 323.855 -299.420 324.085 -298.920 ;
        RECT 325.105 -301.480 325.335 -298.480 ;
        RECT 326.085 -301.480 326.315 -298.480 ;
        RECT 328.200 -301.480 328.430 -298.480 ;
        RECT 336.210 -300.580 336.440 -299.080 ;
        RECT 337.190 -300.580 337.420 -299.080 ;
        RECT 338.170 -300.580 338.400 -299.080 ;
        RECT 339.255 -299.575 339.485 -299.075 ;
        RECT 340.235 -299.575 340.465 -299.075 ;
        RECT 341.215 -299.575 341.445 -299.075 ;
        RECT 342.195 -299.575 342.425 -299.075 ;
        RECT 343.445 -301.635 343.675 -298.635 ;
        RECT 344.425 -301.635 344.655 -298.635 ;
        RECT 346.540 -301.635 346.770 -298.635 ;
        RECT 363.635 -300.340 363.865 -298.840 ;
        RECT 364.615 -300.340 364.845 -298.840 ;
        RECT 365.595 -300.340 365.825 -298.840 ;
        RECT 366.680 -299.335 366.910 -298.835 ;
        RECT 367.660 -299.335 367.890 -298.835 ;
        RECT 368.640 -299.335 368.870 -298.835 ;
        RECT 369.620 -299.335 369.850 -298.835 ;
        RECT 370.870 -301.395 371.100 -298.395 ;
        RECT 371.850 -301.395 372.080 -298.395 ;
        RECT 373.965 -301.395 374.195 -298.395 ;
        RECT 381.975 -300.495 382.205 -298.995 ;
        RECT 382.955 -300.495 383.185 -298.995 ;
        RECT 383.935 -300.495 384.165 -298.995 ;
        RECT 385.020 -299.490 385.250 -298.990 ;
        RECT 386.000 -299.490 386.230 -298.990 ;
        RECT 386.980 -299.490 387.210 -298.990 ;
        RECT 387.960 -299.490 388.190 -298.990 ;
        RECT 389.210 -301.550 389.440 -298.550 ;
        RECT 390.190 -301.550 390.420 -298.550 ;
        RECT 392.305 -301.550 392.535 -298.550 ;
        RECT 410.455 -300.150 410.685 -298.650 ;
        RECT 411.435 -300.150 411.665 -298.650 ;
        RECT 412.415 -300.150 412.645 -298.650 ;
        RECT 413.500 -299.145 413.730 -298.645 ;
        RECT 414.480 -299.145 414.710 -298.645 ;
        RECT 415.460 -299.145 415.690 -298.645 ;
        RECT 416.440 -299.145 416.670 -298.645 ;
        RECT 417.690 -301.205 417.920 -298.205 ;
        RECT 418.670 -301.205 418.900 -298.205 ;
        RECT 420.785 -301.205 421.015 -298.205 ;
        RECT 428.795 -300.305 429.025 -298.805 ;
        RECT 429.775 -300.305 430.005 -298.805 ;
        RECT 430.755 -300.305 430.985 -298.805 ;
        RECT 431.840 -299.300 432.070 -298.800 ;
        RECT 432.820 -299.300 433.050 -298.800 ;
        RECT 433.800 -299.300 434.030 -298.800 ;
        RECT 434.780 -299.300 435.010 -298.800 ;
        RECT 436.030 -301.360 436.260 -298.360 ;
        RECT 437.010 -301.360 437.240 -298.360 ;
        RECT 439.125 -301.360 439.355 -298.360 ;
        RECT -88.410 -305.995 -88.180 -304.995 ;
        RECT -87.430 -305.995 -87.200 -304.995 ;
        RECT -86.450 -305.995 -86.220 -304.995 ;
        RECT -85.470 -305.995 -85.240 -304.995 ;
        RECT -83.545 -305.850 -83.315 -304.350 ;
        RECT -82.565 -305.850 -82.335 -304.350 ;
        RECT -81.585 -305.850 -81.355 -304.350 ;
        RECT -80.500 -304.845 -80.270 -304.345 ;
        RECT -79.520 -304.845 -79.290 -304.345 ;
        RECT -78.540 -304.845 -78.310 -304.345 ;
        RECT -77.560 -304.845 -77.330 -304.345 ;
        RECT -19.710 -306.425 -19.140 -303.270 ;
        RECT -6.900 -303.990 -6.285 -303.310 ;
        RECT -6.875 -306.250 -6.305 -303.990 ;
        RECT 5.515 -304.160 7.045 -303.850 ;
        RECT 5.515 -304.165 6.130 -304.160 ;
        RECT 5.540 -306.250 6.110 -304.165 ;
        RECT -19.730 -307.105 -19.115 -306.425 ;
        RECT -6.895 -306.930 -6.280 -306.250 ;
        RECT 5.520 -306.930 6.135 -306.250 ;
        RECT -107.790 -310.645 -107.560 -309.645 ;
        RECT -106.810 -310.645 -106.580 -309.645 ;
        RECT -104.100 -310.645 -103.870 -309.645 ;
        RECT -103.120 -310.645 -102.890 -309.645 ;
        RECT -102.140 -310.645 -101.910 -309.645 ;
        RECT -101.160 -310.645 -100.930 -309.645 ;
        RECT -94.740 -311.465 -93.860 -308.310 ;
        RECT -26.370 -310.215 -26.140 -309.215 ;
        RECT -25.390 -310.215 -25.160 -309.215 ;
        RECT -24.410 -310.215 -24.180 -309.215 ;
        RECT -23.840 -310.215 -23.610 -309.215 ;
        RECT -22.860 -310.215 -22.630 -309.215 ;
        RECT -22.295 -310.215 -22.065 -309.215 ;
        RECT -21.315 -310.215 -21.085 -309.215 ;
        RECT -13.870 -310.215 -13.640 -309.215 ;
        RECT -12.890 -310.215 -12.660 -309.215 ;
        RECT -11.910 -310.215 -11.680 -309.215 ;
        RECT -11.340 -310.215 -11.110 -309.215 ;
        RECT -10.360 -310.215 -10.130 -309.215 ;
        RECT -9.795 -310.215 -9.565 -309.215 ;
        RECT -8.815 -310.215 -8.585 -309.215 ;
        RECT -1.370 -310.215 -1.140 -309.215 ;
        RECT -0.390 -310.215 -0.160 -309.215 ;
        RECT 0.590 -310.215 0.820 -309.215 ;
        RECT 1.160 -310.215 1.390 -309.215 ;
        RECT 2.140 -310.215 2.370 -309.215 ;
        RECT 2.705 -310.215 2.935 -309.215 ;
        RECT 3.685 -310.215 3.915 -309.215 ;
        RECT 11.130 -310.215 11.360 -309.215 ;
        RECT 12.110 -310.215 12.340 -309.215 ;
        RECT 13.090 -310.215 13.320 -309.215 ;
        RECT 13.660 -310.215 13.890 -309.215 ;
        RECT 14.640 -310.215 14.870 -309.215 ;
        RECT 15.205 -310.215 15.435 -309.215 ;
        RECT 16.185 -310.215 16.415 -309.215 ;
        RECT 23.630 -310.215 23.860 -309.215 ;
        RECT 24.610 -310.215 24.840 -309.215 ;
        RECT 25.590 -310.215 25.820 -309.215 ;
        RECT 26.160 -310.215 26.390 -309.215 ;
        RECT 27.140 -310.215 27.370 -309.215 ;
        RECT 27.705 -310.215 27.935 -309.215 ;
        RECT 28.685 -310.215 28.915 -309.215 ;
        RECT 38.630 -310.215 38.860 -309.215 ;
        RECT 39.610 -310.215 39.840 -309.215 ;
        RECT 40.590 -310.215 40.820 -309.215 ;
        RECT 41.160 -310.215 41.390 -309.215 ;
        RECT 42.140 -310.215 42.370 -309.215 ;
        RECT 42.705 -310.215 42.935 -309.215 ;
        RECT 43.685 -310.215 43.915 -309.215 ;
        RECT 69.265 -309.400 69.495 -308.400 ;
        RECT 70.245 -309.400 70.475 -308.400 ;
        RECT 71.225 -309.400 71.455 -308.400 ;
        RECT 73.450 -309.400 73.680 -308.400 ;
        RECT 74.430 -309.400 74.660 -308.400 ;
        RECT 75.410 -309.400 75.640 -308.400 ;
        RECT 82.765 -309.400 82.995 -308.400 ;
        RECT 83.745 -309.400 83.975 -308.400 ;
        RECT 84.725 -309.400 84.955 -308.400 ;
        RECT 86.950 -309.400 87.180 -308.400 ;
        RECT 87.930 -309.400 88.160 -308.400 ;
        RECT 88.910 -309.400 89.140 -308.400 ;
    END
  END VDD
  PIN VSS
    ANTENNAGATEAREA 141.000000 ;
    ANTENNADIFFAREA 1162.211548 ;
    PORT
      LAYER pwell ;
        RECT -64.340 595.535 -63.670 599.530 ;
        RECT -52.850 596.365 -52.195 599.270 ;
        RECT -60.085 591.370 -59.430 594.275 ;
        RECT -50.305 593.150 -49.740 595.655 ;
        RECT -62.540 588.155 -61.975 590.660 ;
        RECT -51.205 588.455 -50.550 591.360 ;
        RECT -46.990 586.760 -45.925 594.385 ;
        RECT -64.185 577.195 -63.515 581.190 ;
        RECT -52.695 578.025 -52.040 580.930 ;
        RECT -59.930 573.030 -59.275 575.935 ;
        RECT -50.150 574.810 -49.585 577.315 ;
        RECT -46.920 577.235 -46.250 581.230 ;
        RECT -35.430 578.065 -34.775 580.970 ;
        RECT -42.665 573.070 -42.010 575.975 ;
        RECT -32.885 574.850 -32.320 577.355 ;
        RECT -62.385 569.815 -61.820 572.320 ;
        RECT -51.050 570.115 -50.395 573.020 ;
        RECT -45.120 569.855 -44.555 572.360 ;
        RECT -33.785 570.155 -33.130 573.060 ;
        RECT -64.530 548.715 -63.860 552.710 ;
        RECT -53.040 549.545 -52.385 552.450 ;
        RECT -60.275 544.550 -59.620 547.455 ;
        RECT -50.495 546.330 -49.930 548.835 ;
        RECT -62.730 541.335 -62.165 543.840 ;
        RECT -51.395 541.635 -50.740 544.540 ;
        RECT -47.180 539.940 -46.115 547.565 ;
        RECT -64.375 530.375 -63.705 534.370 ;
        RECT -52.885 531.205 -52.230 534.110 ;
        RECT -60.120 526.210 -59.465 529.115 ;
        RECT -50.340 527.990 -49.775 530.495 ;
        RECT -47.110 530.415 -46.440 534.410 ;
        RECT -35.620 531.245 -34.965 534.150 ;
        RECT -42.855 526.250 -42.200 529.155 ;
        RECT -33.075 528.030 -32.510 530.535 ;
        RECT -62.575 522.995 -62.010 525.500 ;
        RECT -51.240 523.295 -50.585 526.200 ;
        RECT -45.310 523.035 -44.745 525.540 ;
        RECT -33.975 523.335 -33.320 526.240 ;
        RECT -64.615 502.950 -63.945 506.945 ;
        RECT -53.125 503.780 -52.470 506.685 ;
        RECT -60.360 498.785 -59.705 501.690 ;
        RECT -50.580 500.565 -50.015 503.070 ;
        RECT -62.815 495.570 -62.250 498.075 ;
        RECT -51.480 495.870 -50.825 498.775 ;
        RECT -47.265 494.175 -46.200 501.800 ;
        RECT -64.460 484.610 -63.790 488.605 ;
        RECT -52.970 485.440 -52.315 488.345 ;
        RECT -60.205 480.445 -59.550 483.350 ;
        RECT -50.425 482.225 -49.860 484.730 ;
        RECT -47.195 484.650 -46.525 488.645 ;
        RECT -35.705 485.480 -35.050 488.385 ;
        RECT -42.940 480.485 -42.285 483.390 ;
        RECT -33.160 482.265 -32.595 484.770 ;
        RECT -62.660 477.230 -62.095 479.735 ;
        RECT -51.325 477.530 -50.670 480.435 ;
        RECT -45.395 477.270 -44.830 479.775 ;
        RECT -34.060 477.570 -33.405 480.475 ;
        RECT -64.945 459.180 -64.275 463.175 ;
        RECT -53.455 460.010 -52.800 462.915 ;
        RECT -60.690 455.015 -60.035 457.920 ;
        RECT -50.910 456.795 -50.345 459.300 ;
        RECT -63.145 451.800 -62.580 454.305 ;
        RECT -51.810 452.100 -51.155 455.005 ;
        RECT -47.595 450.405 -46.530 458.030 ;
        RECT -64.790 440.840 -64.120 444.835 ;
        RECT -53.300 441.670 -52.645 444.575 ;
        RECT -60.535 436.675 -59.880 439.580 ;
        RECT -50.755 438.455 -50.190 440.960 ;
        RECT -47.525 440.880 -46.855 444.875 ;
        RECT -36.035 441.710 -35.380 444.615 ;
        RECT -43.270 436.715 -42.615 439.620 ;
        RECT -33.490 438.495 -32.925 441.000 ;
        RECT -62.990 433.460 -62.425 435.965 ;
        RECT -51.655 433.760 -51.000 436.665 ;
        RECT -45.725 433.500 -45.160 436.005 ;
        RECT -34.390 433.800 -33.735 436.705 ;
        RECT -65.115 413.190 -64.445 417.185 ;
        RECT -53.625 414.020 -52.970 416.925 ;
        RECT -60.860 409.025 -60.205 411.930 ;
        RECT -51.080 410.805 -50.515 413.310 ;
        RECT -63.315 405.810 -62.750 408.315 ;
        RECT -51.980 406.110 -51.325 409.015 ;
        RECT -47.765 404.415 -46.700 412.040 ;
        RECT -64.960 394.850 -64.290 398.845 ;
        RECT -53.470 395.680 -52.815 398.585 ;
        RECT -60.705 390.685 -60.050 393.590 ;
        RECT -50.925 392.465 -50.360 394.970 ;
        RECT -47.695 394.890 -47.025 398.885 ;
        RECT -36.205 395.720 -35.550 398.625 ;
        RECT -43.440 390.725 -42.785 393.630 ;
        RECT -33.660 392.505 -33.095 395.010 ;
        RECT -63.160 387.470 -62.595 389.975 ;
        RECT -51.825 387.770 -51.170 390.675 ;
        RECT -45.895 387.510 -45.330 390.015 ;
        RECT -34.560 387.810 -33.905 390.715 ;
        RECT -64.920 368.875 -64.250 372.870 ;
        RECT -53.430 369.705 -52.775 372.610 ;
        RECT -60.665 364.710 -60.010 367.615 ;
        RECT -50.885 366.490 -50.320 368.995 ;
        RECT -63.120 361.495 -62.555 364.000 ;
        RECT -51.785 361.795 -51.130 364.700 ;
        RECT -47.570 360.100 -46.505 367.725 ;
        RECT -64.765 350.535 -64.095 354.530 ;
        RECT -53.275 351.365 -52.620 354.270 ;
        RECT -60.510 346.370 -59.855 349.275 ;
        RECT -50.730 348.150 -50.165 350.655 ;
        RECT -47.500 350.575 -46.830 354.570 ;
        RECT -36.010 351.405 -35.355 354.310 ;
        RECT -43.245 346.410 -42.590 349.315 ;
        RECT -33.465 348.190 -32.900 350.695 ;
        RECT -62.965 343.155 -62.400 345.660 ;
        RECT -51.630 343.455 -50.975 346.360 ;
        RECT -45.700 343.195 -45.135 345.700 ;
        RECT -34.365 343.495 -33.710 346.400 ;
        RECT -64.865 326.675 -64.195 330.670 ;
        RECT -53.375 327.505 -52.720 330.410 ;
        RECT -60.610 322.510 -59.955 325.415 ;
        RECT -50.830 324.290 -50.265 326.795 ;
        RECT -63.065 319.295 -62.500 321.800 ;
        RECT -51.730 319.595 -51.075 322.500 ;
        RECT -47.515 317.900 -46.450 325.525 ;
        RECT -64.710 308.335 -64.040 312.330 ;
        RECT -53.220 309.165 -52.565 312.070 ;
        RECT -60.455 304.170 -59.800 307.075 ;
        RECT -50.675 305.950 -50.110 308.455 ;
        RECT -47.445 308.375 -46.775 312.370 ;
        RECT -35.955 309.205 -35.300 312.110 ;
        RECT -43.190 304.210 -42.535 307.115 ;
        RECT -33.410 305.990 -32.845 308.495 ;
        RECT -62.910 300.955 -62.345 303.460 ;
        RECT -51.575 301.255 -50.920 304.160 ;
        RECT -45.645 300.995 -45.080 303.500 ;
        RECT -34.310 301.295 -33.655 304.200 ;
        RECT -47.985 275.825 -47.240 289.720 ;
        RECT -42.910 286.515 -42.310 289.445 ;
        RECT -41.010 286.555 -40.410 289.485 ;
        RECT -41.010 282.370 -40.410 285.300 ;
        RECT -42.910 277.800 -42.310 280.730 ;
        RECT -54.175 271.865 -53.575 274.795 ;
        RECT -53.560 271.995 -52.895 274.650 ;
        RECT -42.910 273.015 -42.310 275.945 ;
        RECT -41.010 273.055 -40.410 275.985 ;
        RECT -51.385 262.615 -50.800 269.245 ;
        RECT -41.010 268.870 -40.410 271.800 ;
        RECT -42.910 264.300 -42.310 267.230 ;
        RECT -51.720 257.860 -51.015 261.105 ;
        RECT -42.910 259.890 -42.310 262.820 ;
        RECT -51.720 253.130 -51.015 256.375 ;
        RECT -38.600 253.275 -37.810 257.820 ;
        RECT -65.690 245.915 -65.090 248.845 ;
        RECT -63.790 245.875 -63.190 248.805 ;
        RECT -65.690 241.730 -65.090 244.660 ;
        RECT -63.790 237.160 -63.190 240.090 ;
        RECT -65.690 232.415 -65.090 235.345 ;
        RECT -63.790 232.375 -63.190 235.305 ;
        RECT -65.690 228.230 -65.090 231.160 ;
        RECT -63.790 223.660 -63.190 226.590 ;
        RECT -63.790 219.250 -63.190 222.180 ;
        RECT -64.745 200.195 -64.005 203.615 ;
        RECT -53.490 200.245 -52.750 203.665 ;
        RECT -41.660 200.245 -40.920 203.665 ;
        RECT -30.405 200.195 -29.665 203.615 ;
        RECT -64.745 185.195 -64.005 188.615 ;
        RECT -52.480 186.135 -51.895 192.765 ;
        RECT -42.515 186.135 -41.930 192.765 ;
        RECT -30.405 185.195 -29.665 188.615 ;
        RECT -53.390 181.595 -52.825 184.100 ;
        RECT -41.585 181.595 -41.020 184.100 ;
        RECT -55.935 177.980 -55.280 180.885 ;
        RECT -39.130 177.980 -38.475 180.885 ;
        RECT -64.745 172.695 -64.005 176.115 ;
        RECT -53.400 173.570 -52.835 176.075 ;
        RECT -41.575 173.570 -41.010 176.075 ;
        RECT -55.945 169.955 -55.290 172.860 ;
        RECT -39.120 169.955 -38.465 172.860 ;
        RECT -30.405 172.695 -29.665 176.115 ;
        RECT -64.745 160.195 -64.005 163.615 ;
        RECT -52.435 161.325 -51.850 167.955 ;
        RECT -42.560 161.325 -41.975 167.955 ;
        RECT -30.405 160.195 -29.665 163.615 ;
        RECT -55.345 156.730 -54.745 159.660 ;
        RECT -39.665 156.730 -39.065 159.660 ;
        RECT -55.345 152.320 -54.745 155.250 ;
        RECT -39.665 152.320 -39.065 155.250 ;
        RECT -64.745 147.695 -64.005 151.115 ;
        RECT -53.445 147.750 -52.845 150.680 ;
        RECT -41.565 147.750 -40.965 150.680 ;
        RECT -30.405 147.695 -29.665 151.115 ;
        RECT -55.345 143.605 -54.745 146.535 ;
        RECT -53.445 143.565 -52.845 146.495 ;
        RECT -41.565 143.565 -40.965 146.495 ;
        RECT -39.665 143.605 -39.065 146.535 ;
        RECT -55.345 138.820 -54.745 141.750 ;
        RECT -39.665 138.820 -39.065 141.750 ;
        RECT -64.745 135.195 -64.005 138.615 ;
        RECT -53.445 134.250 -52.845 137.180 ;
        RECT -41.565 134.250 -40.965 137.180 ;
        RECT -30.405 135.195 -29.665 138.615 ;
        RECT -55.345 130.105 -54.745 133.035 ;
        RECT -53.445 130.065 -52.845 132.995 ;
        RECT -41.565 130.065 -40.965 132.995 ;
        RECT -39.665 130.105 -39.065 133.035 ;
        RECT -30.460 131.350 -29.860 134.280 ;
        RECT -56.195 122.170 -55.525 126.165 ;
        RECT -31.525 122.035 -30.855 126.030 ;
        RECT -54.010 117.360 -53.410 120.290 ;
        RECT -29.375 117.360 -28.775 120.290 ;
        RECT -54.010 112.950 -53.410 115.880 ;
        RECT -29.375 112.950 -28.775 115.880 ;
        RECT -52.110 108.380 -51.510 111.310 ;
        RECT -27.475 108.380 -26.875 111.310 ;
        RECT -54.010 104.235 -53.410 107.165 ;
        RECT -52.110 104.195 -51.510 107.125 ;
        RECT -45.510 103.975 -44.855 106.880 ;
        RECT -54.010 99.450 -53.410 102.380 ;
        RECT -47.965 100.760 -47.400 103.265 ;
        RECT -34.035 103.145 -33.365 107.140 ;
        RECT -29.375 104.235 -28.775 107.165 ;
        RECT -27.475 104.195 -26.875 107.125 ;
        RECT -38.275 98.980 -37.620 101.885 ;
        RECT -29.375 99.450 -28.775 102.380 ;
        RECT -52.110 94.880 -51.510 97.810 ;
        RECT -47.155 96.065 -46.500 98.970 ;
        RECT -35.730 95.765 -35.165 98.270 ;
        RECT -27.475 94.880 -26.875 97.810 ;
        RECT -54.010 90.735 -53.410 93.665 ;
        RECT -52.110 90.695 -51.510 93.625 ;
        RECT -29.375 90.735 -28.775 93.665 ;
        RECT -27.475 90.695 -26.875 93.625 ;
        RECT -65.630 79.030 -64.975 81.935 ;
        RECT -68.085 75.815 -67.520 78.320 ;
        RECT -54.155 78.200 -53.485 82.195 ;
        RECT -40.630 79.030 -39.975 81.935 ;
        RECT -58.395 74.035 -57.740 76.940 ;
        RECT -43.085 75.815 -42.520 78.320 ;
        RECT -29.155 78.200 -28.485 82.195 ;
        RECT -33.395 74.035 -32.740 76.940 ;
        RECT -67.275 71.120 -66.620 74.025 ;
        RECT -55.850 70.820 -55.285 73.325 ;
        RECT -42.275 71.120 -41.620 74.025 ;
        RECT -30.850 70.820 -30.285 73.325 ;
        RECT -59.610 63.735 -58.905 66.980 ;
        RECT -59.605 59.210 -58.900 62.455 ;
        RECT -43.900 61.895 -43.315 68.525 ;
        RECT -31.320 65.855 -30.665 68.760 ;
        RECT -33.775 62.640 -33.210 65.145 ;
        RECT -64.110 52.100 -63.525 58.730 ;
        RECT -61.435 53.300 -60.645 57.845 ;
        RECT -40.865 56.145 -40.210 59.050 ;
        RECT -43.320 52.930 -42.755 55.435 ;
        RECT -34.220 52.745 -33.635 59.375 ;
        RECT 85.545 44.830 86.705 51.050 ;
        RECT 346.040 48.060 461.860 50.410 ;
        RECT 40.410 21.660 62.880 22.650 ;
        RECT 127.905 17.530 238.300 18.765 ;
        RECT 98.795 13.745 101.725 14.345 ;
        RECT 103.045 13.745 105.975 14.345 ;
        RECT 103.045 13.060 105.975 13.660 ;
        RECT 13.970 11.965 15.625 12.670 ;
        RECT 2.695 11.300 15.625 11.965 ;
        RECT 2.695 11.230 5.765 11.300 ;
        RECT 7.675 11.240 15.625 11.300 ;
        RECT 7.675 11.230 14.955 11.240 ;
        RECT 2.825 10.730 4.090 11.230 ;
        RECT 12.145 10.730 14.955 11.230 ;
        RECT 22.400 7.920 25.330 8.520 ;
        RECT 26.650 7.920 29.580 8.520 ;
        RECT 26.650 7.235 29.580 7.835 ;
        RECT 39.180 4.065 75.445 4.955 ;
        RECT 2.825 3.080 4.090 3.580 ;
        RECT 12.145 3.080 14.955 3.580 ;
        RECT 2.695 3.010 5.765 3.080 ;
        RECT 7.675 3.010 14.955 3.080 ;
        RECT 2.695 2.345 14.955 3.010 ;
        RECT 99.655 -3.005 102.585 -2.405 ;
        RECT 103.905 -3.005 106.835 -2.405 ;
        RECT 103.905 -3.690 106.835 -3.090 ;
        RECT 22.475 -5.530 25.405 -4.930 ;
        RECT 26.725 -5.530 29.655 -4.930 ;
        RECT 26.725 -6.215 29.655 -5.615 ;
        RECT 127.905 -6.015 129.140 17.530 ;
        RECT 151.395 13.140 158.335 14.025 ;
        RECT 175.070 13.250 182.010 14.135 ;
        RECT 183.675 13.035 190.615 13.920 ;
        RECT 195.755 11.530 198.685 12.130 ;
        RECT 200.165 11.530 203.095 12.130 ;
        RECT 208.880 11.530 211.810 12.130 ;
        RECT 213.665 11.530 216.595 12.130 ;
        RECT 222.380 11.530 225.310 12.130 ;
        RECT 204.735 9.630 207.665 10.230 ;
        RECT 208.920 9.630 211.850 10.230 ;
        RECT 218.235 9.630 221.165 10.230 ;
        RECT 222.420 9.630 225.350 10.230 ;
        RECT 227.720 10.080 230.650 10.680 ;
        RECT 138.690 -1.420 147.445 -0.705 ;
        RECT 162.965 -1.455 171.720 -0.740 ;
        RECT 151.395 -2.625 158.335 -1.740 ;
        RECT 175.070 -2.510 182.010 -1.625 ;
        RECT 183.675 -2.295 190.615 -1.410 ;
        RECT 237.065 -6.015 238.300 17.530 ;
        RECT 255.570 7.950 291.835 8.840 ;
        RECT 127.905 -7.250 238.300 -6.015 ;
        RECT 254.555 -6.605 290.820 -5.715 ;
        RECT 38.975 -9.715 75.240 -8.825 ;
        RECT 311.790 -17.335 314.720 -16.735 ;
        RECT 316.040 -17.335 318.970 -16.735 ;
        RECT 316.040 -18.020 318.970 -17.420 ;
        RECT 254.555 -21.840 290.820 -20.950 ;
      LAYER li1 ;
        RECT -64.360 598.500 -63.795 599.825 ;
        RECT -64.360 598.470 -63.150 598.500 ;
        RECT -64.360 598.300 -61.735 598.470 ;
        RECT -64.360 598.265 -63.150 598.300 ;
        RECT -64.360 597.290 -63.795 598.265 ;
        RECT -52.730 598.065 -52.300 600.140 ;
        RECT -53.510 597.895 -52.300 598.065 ;
        RECT -52.730 597.740 -52.300 597.895 ;
        RECT -52.730 597.435 -49.960 597.740 ;
        RECT -64.360 597.260 -63.200 597.290 ;
        RECT -64.360 597.090 -61.735 597.260 ;
        RECT -64.360 597.055 -63.200 597.090 ;
        RECT -52.730 597.085 -52.300 597.435 ;
        RECT -64.360 596.310 -63.795 597.055 ;
        RECT -53.510 596.915 -52.300 597.085 ;
        RECT -64.360 596.280 -63.205 596.310 ;
        RECT -64.360 596.110 -61.735 596.280 ;
        RECT -52.730 596.215 -52.300 596.915 ;
        RECT -64.360 596.075 -63.205 596.110 ;
        RECT -64.360 592.745 -63.795 596.075 ;
        RECT -50.265 595.890 -49.960 597.435 ;
        RECT -50.265 595.490 -49.820 595.890 ;
        RECT -59.980 593.070 -59.550 594.295 ;
        RECT -50.250 594.040 -49.820 595.490 ;
        RECT -51.975 593.870 -49.820 594.040 ;
        RECT -50.435 593.865 -49.820 593.870 ;
        RECT -59.980 592.900 -58.770 593.070 ;
        RECT -50.250 592.995 -49.820 593.865 ;
        RECT -59.980 592.745 -59.550 592.900 ;
        RECT -64.360 592.440 -59.550 592.745 ;
        RECT -62.320 590.530 -62.015 592.440 ;
        RECT -59.980 592.090 -59.550 592.440 ;
        RECT -51.085 592.565 -49.820 592.995 ;
        RECT -46.860 593.690 -46.055 594.255 ;
        RECT -46.860 593.685 -45.470 593.690 ;
        RECT -46.860 593.515 -44.025 593.685 ;
        RECT -46.860 593.505 -45.470 593.515 ;
        RECT -59.980 591.920 -58.770 592.090 ;
        RECT -59.980 591.220 -59.550 591.920 ;
        RECT -62.410 590.495 -62.015 590.530 ;
        RECT -62.410 589.045 -62.105 590.495 ;
        RECT -51.085 590.155 -50.655 592.565 ;
        RECT -52.365 589.985 -50.655 590.155 ;
        RECT -51.085 589.175 -50.655 589.985 ;
        RECT -62.410 588.875 -60.305 589.045 ;
        RECT -52.365 589.005 -50.655 589.175 ;
        RECT -62.410 588.870 -61.845 588.875 ;
        RECT -62.410 588.285 -62.105 588.870 ;
        RECT -59.645 587.960 -59.375 588.635 ;
        RECT -51.085 588.305 -50.655 589.005 ;
        RECT -46.860 592.055 -46.055 593.505 ;
        RECT -46.860 591.885 -43.025 592.055 ;
        RECT -46.860 591.870 -45.475 591.885 ;
        RECT -46.860 591.415 -46.055 591.870 ;
        RECT -46.860 591.405 -45.480 591.415 ;
        RECT -46.860 591.235 -43.025 591.405 ;
        RECT -46.860 591.230 -45.480 591.235 ;
        RECT -59.605 587.860 -59.405 587.960 ;
        RECT -59.595 586.470 -59.415 587.860 ;
        RECT -46.860 587.640 -46.055 591.230 ;
        RECT -46.860 587.455 -46.035 587.640 ;
        RECT -46.860 587.450 -45.480 587.455 ;
        RECT -46.860 587.280 -44.025 587.450 ;
        RECT -46.860 587.270 -45.480 587.280 ;
        RECT -46.860 586.890 -46.035 587.270 ;
        RECT -65.255 585.790 -59.415 586.470 ;
        RECT -65.255 568.595 -64.575 585.790 ;
        RECT -46.600 585.150 -46.035 586.890 ;
        RECT -46.940 584.585 -46.035 585.150 ;
        RECT -64.205 580.160 -63.640 581.485 ;
        RECT -64.205 580.130 -62.995 580.160 ;
        RECT -64.205 579.960 -61.580 580.130 ;
        RECT -64.205 579.925 -62.995 579.960 ;
        RECT -64.205 578.950 -63.640 579.925 ;
        RECT -52.575 579.725 -52.145 581.800 ;
        RECT -53.355 579.555 -52.145 579.725 ;
        RECT -52.575 579.400 -52.145 579.555 ;
        RECT -46.940 580.200 -46.375 584.585 ;
        RECT -46.940 580.170 -45.730 580.200 ;
        RECT -46.940 580.000 -44.315 580.170 ;
        RECT -46.940 579.965 -45.730 580.000 ;
        RECT -52.575 579.095 -49.805 579.400 ;
        RECT -64.205 578.920 -63.045 578.950 ;
        RECT -64.205 578.750 -61.580 578.920 ;
        RECT -64.205 578.715 -63.045 578.750 ;
        RECT -52.575 578.745 -52.145 579.095 ;
        RECT -64.205 577.970 -63.640 578.715 ;
        RECT -53.355 578.575 -52.145 578.745 ;
        RECT -64.205 577.940 -63.050 577.970 ;
        RECT -64.205 577.770 -61.580 577.940 ;
        RECT -52.575 577.875 -52.145 578.575 ;
        RECT -64.205 577.735 -63.050 577.770 ;
        RECT -64.205 574.405 -63.640 577.735 ;
        RECT -50.110 577.550 -49.805 579.095 ;
        RECT -46.940 578.990 -46.375 579.965 ;
        RECT -35.310 579.765 -34.880 581.840 ;
        RECT -36.090 579.595 -34.880 579.765 ;
        RECT -35.310 579.440 -34.880 579.595 ;
        RECT -35.310 579.135 -32.540 579.440 ;
        RECT -46.940 578.960 -45.780 578.990 ;
        RECT -46.940 578.790 -44.315 578.960 ;
        RECT -46.940 578.755 -45.780 578.790 ;
        RECT -35.310 578.785 -34.880 579.135 ;
        RECT -46.940 578.010 -46.375 578.755 ;
        RECT -36.090 578.615 -34.880 578.785 ;
        RECT -46.940 577.980 -45.785 578.010 ;
        RECT -46.940 577.810 -44.315 577.980 ;
        RECT -35.310 577.915 -34.880 578.615 ;
        RECT -46.940 577.775 -45.785 577.810 ;
        RECT -50.110 577.150 -49.665 577.550 ;
        RECT -59.825 574.730 -59.395 575.955 ;
        RECT -50.095 575.700 -49.665 577.150 ;
        RECT -51.820 575.530 -49.665 575.700 ;
        RECT -50.280 575.525 -49.665 575.530 ;
        RECT -59.825 574.560 -58.615 574.730 ;
        RECT -50.095 574.655 -49.665 575.525 ;
        RECT -59.825 574.405 -59.395 574.560 ;
        RECT -64.205 574.100 -59.395 574.405 ;
        RECT -62.165 572.190 -61.860 574.100 ;
        RECT -59.825 573.750 -59.395 574.100 ;
        RECT -50.930 574.225 -49.665 574.655 ;
        RECT -46.940 574.445 -46.375 577.775 ;
        RECT -32.845 577.590 -32.540 579.135 ;
        RECT -32.845 577.190 -32.400 577.590 ;
        RECT -32.830 576.515 -32.400 577.190 ;
        RECT -30.620 576.515 -28.090 584.845 ;
        RECT -42.560 574.770 -42.130 575.995 ;
        RECT -32.830 575.740 -28.090 576.515 ;
        RECT -34.555 575.570 -28.090 575.740 ;
        RECT -33.015 575.565 -28.090 575.570 ;
        RECT -32.830 575.460 -28.090 575.565 ;
        RECT -42.560 574.600 -41.350 574.770 ;
        RECT -32.830 574.695 -32.400 575.460 ;
        RECT -42.560 574.445 -42.130 574.600 ;
        RECT -59.825 573.580 -58.615 573.750 ;
        RECT -59.825 572.880 -59.395 573.580 ;
        RECT -62.255 572.155 -61.860 572.190 ;
        RECT -62.255 570.705 -61.950 572.155 ;
        RECT -50.930 571.815 -50.500 574.225 ;
        RECT -46.940 574.140 -42.130 574.445 ;
        RECT -44.900 572.230 -44.595 574.140 ;
        RECT -42.560 573.790 -42.130 574.140 ;
        RECT -33.665 574.265 -32.400 574.695 ;
        RECT -42.560 573.620 -41.350 573.790 ;
        RECT -42.560 572.920 -42.130 573.620 ;
        RECT -52.210 571.645 -50.500 571.815 ;
        RECT -50.930 570.835 -50.500 571.645 ;
        RECT -62.255 570.535 -60.150 570.705 ;
        RECT -52.210 570.665 -50.500 570.835 ;
        RECT -62.255 570.530 -61.690 570.535 ;
        RECT -62.255 569.945 -61.950 570.530 ;
        RECT -59.490 569.620 -59.220 570.295 ;
        RECT -50.930 569.965 -50.500 570.665 ;
        RECT -44.990 572.195 -44.595 572.230 ;
        RECT -44.990 570.745 -44.685 572.195 ;
        RECT -33.665 571.855 -33.235 574.265 ;
        RECT -34.945 571.685 -33.235 571.855 ;
        RECT -33.665 570.875 -33.235 571.685 ;
        RECT -44.990 570.575 -42.885 570.745 ;
        RECT -34.945 570.705 -33.235 570.875 ;
        RECT -44.990 570.570 -44.425 570.575 ;
        RECT -44.990 569.985 -44.685 570.570 ;
        RECT -33.665 570.005 -33.235 570.705 ;
        RECT -59.450 569.520 -59.250 569.620 ;
        RECT -80.800 568.475 -64.575 568.595 ;
        RECT -59.440 568.475 -59.260 569.520 ;
        RECT -80.800 567.915 -59.260 568.475 ;
        RECT -80.800 42.775 -80.120 567.915 ;
        RECT -65.255 567.795 -59.260 567.915 ;
        RECT -59.440 566.880 -59.260 567.795 ;
        RECT -64.550 551.680 -63.985 553.005 ;
        RECT -64.550 551.650 -63.340 551.680 ;
        RECT -64.550 551.480 -61.925 551.650 ;
        RECT -64.550 551.445 -63.340 551.480 ;
        RECT -64.550 550.470 -63.985 551.445 ;
        RECT -52.920 551.245 -52.490 553.320 ;
        RECT -53.700 551.075 -52.490 551.245 ;
        RECT -52.920 550.920 -52.490 551.075 ;
        RECT -52.920 550.615 -50.150 550.920 ;
        RECT -64.550 550.440 -63.390 550.470 ;
        RECT -64.550 550.270 -61.925 550.440 ;
        RECT -64.550 550.235 -63.390 550.270 ;
        RECT -52.920 550.265 -52.490 550.615 ;
        RECT -64.550 549.490 -63.985 550.235 ;
        RECT -53.700 550.095 -52.490 550.265 ;
        RECT -64.550 549.460 -63.395 549.490 ;
        RECT -64.550 549.290 -61.925 549.460 ;
        RECT -52.920 549.395 -52.490 550.095 ;
        RECT -64.550 549.255 -63.395 549.290 ;
        RECT -64.550 545.925 -63.985 549.255 ;
        RECT -50.455 549.070 -50.150 550.615 ;
        RECT -50.455 548.670 -50.010 549.070 ;
        RECT -60.170 546.250 -59.740 547.475 ;
        RECT -50.440 547.220 -50.010 548.670 ;
        RECT -52.165 547.050 -50.010 547.220 ;
        RECT -50.625 547.045 -50.010 547.050 ;
        RECT -60.170 546.080 -58.960 546.250 ;
        RECT -50.440 546.175 -50.010 547.045 ;
        RECT -60.170 545.925 -59.740 546.080 ;
        RECT -64.550 545.620 -59.740 545.925 ;
        RECT -62.510 543.710 -62.205 545.620 ;
        RECT -60.170 545.270 -59.740 545.620 ;
        RECT -51.275 545.745 -50.010 546.175 ;
        RECT -47.050 546.870 -46.245 547.435 ;
        RECT -47.050 546.865 -45.660 546.870 ;
        RECT -47.050 546.695 -44.215 546.865 ;
        RECT -47.050 546.685 -45.660 546.695 ;
        RECT -60.170 545.100 -58.960 545.270 ;
        RECT -60.170 544.400 -59.740 545.100 ;
        RECT -62.600 543.675 -62.205 543.710 ;
        RECT -62.600 542.225 -62.295 543.675 ;
        RECT -51.275 543.335 -50.845 545.745 ;
        RECT -52.555 543.165 -50.845 543.335 ;
        RECT -51.275 542.355 -50.845 543.165 ;
        RECT -62.600 542.055 -60.495 542.225 ;
        RECT -52.555 542.185 -50.845 542.355 ;
        RECT -62.600 542.050 -62.035 542.055 ;
        RECT -62.600 541.465 -62.295 542.050 ;
        RECT -59.835 541.140 -59.565 541.815 ;
        RECT -51.275 541.485 -50.845 542.185 ;
        RECT -47.050 545.235 -46.245 546.685 ;
        RECT -47.050 545.065 -43.215 545.235 ;
        RECT -47.050 545.050 -45.665 545.065 ;
        RECT -47.050 544.595 -46.245 545.050 ;
        RECT -47.050 544.585 -45.670 544.595 ;
        RECT -47.050 544.415 -43.215 544.585 ;
        RECT -47.050 544.410 -45.670 544.415 ;
        RECT -59.795 541.040 -59.595 541.140 ;
        RECT -59.785 539.650 -59.605 541.040 ;
        RECT -47.050 540.820 -46.245 544.410 ;
        RECT -47.050 540.635 -46.225 540.820 ;
        RECT -47.050 540.630 -45.670 540.635 ;
        RECT -47.050 540.460 -44.215 540.630 ;
        RECT -47.050 540.450 -45.670 540.460 ;
        RECT -47.050 540.070 -46.225 540.450 ;
        RECT -65.445 538.970 -59.605 539.650 ;
        RECT -65.445 521.655 -64.765 538.970 ;
        RECT -46.790 538.330 -46.225 540.070 ;
        RECT -47.130 537.765 -46.225 538.330 ;
        RECT -64.395 533.340 -63.830 534.665 ;
        RECT -64.395 533.310 -63.185 533.340 ;
        RECT -64.395 533.140 -61.770 533.310 ;
        RECT -64.395 533.105 -63.185 533.140 ;
        RECT -64.395 532.130 -63.830 533.105 ;
        RECT -52.765 532.905 -52.335 534.980 ;
        RECT -53.545 532.735 -52.335 532.905 ;
        RECT -52.765 532.580 -52.335 532.735 ;
        RECT -47.130 533.380 -46.565 537.765 ;
        RECT -47.130 533.350 -45.920 533.380 ;
        RECT -47.130 533.180 -44.505 533.350 ;
        RECT -47.130 533.145 -45.920 533.180 ;
        RECT -52.765 532.275 -49.995 532.580 ;
        RECT -64.395 532.100 -63.235 532.130 ;
        RECT -64.395 531.930 -61.770 532.100 ;
        RECT -64.395 531.895 -63.235 531.930 ;
        RECT -52.765 531.925 -52.335 532.275 ;
        RECT -64.395 531.150 -63.830 531.895 ;
        RECT -53.545 531.755 -52.335 531.925 ;
        RECT -64.395 531.120 -63.240 531.150 ;
        RECT -64.395 530.950 -61.770 531.120 ;
        RECT -52.765 531.055 -52.335 531.755 ;
        RECT -64.395 530.915 -63.240 530.950 ;
        RECT -64.395 527.585 -63.830 530.915 ;
        RECT -50.300 530.730 -49.995 532.275 ;
        RECT -47.130 532.170 -46.565 533.145 ;
        RECT -35.500 532.945 -35.070 535.020 ;
        RECT -36.280 532.775 -35.070 532.945 ;
        RECT -35.500 532.620 -35.070 532.775 ;
        RECT -35.500 532.315 -32.730 532.620 ;
        RECT -47.130 532.140 -45.970 532.170 ;
        RECT -47.130 531.970 -44.505 532.140 ;
        RECT -47.130 531.935 -45.970 531.970 ;
        RECT -35.500 531.965 -35.070 532.315 ;
        RECT -47.130 531.190 -46.565 531.935 ;
        RECT -36.280 531.795 -35.070 531.965 ;
        RECT -47.130 531.160 -45.975 531.190 ;
        RECT -47.130 530.990 -44.505 531.160 ;
        RECT -35.500 531.095 -35.070 531.795 ;
        RECT -47.130 530.955 -45.975 530.990 ;
        RECT -50.300 530.330 -49.855 530.730 ;
        RECT -60.015 527.910 -59.585 529.135 ;
        RECT -50.285 528.880 -49.855 530.330 ;
        RECT -52.010 528.710 -49.855 528.880 ;
        RECT -50.470 528.705 -49.855 528.710 ;
        RECT -60.015 527.740 -58.805 527.910 ;
        RECT -50.285 527.835 -49.855 528.705 ;
        RECT -60.015 527.585 -59.585 527.740 ;
        RECT -64.395 527.280 -59.585 527.585 ;
        RECT -62.355 525.370 -62.050 527.280 ;
        RECT -60.015 526.930 -59.585 527.280 ;
        RECT -51.120 527.405 -49.855 527.835 ;
        RECT -47.130 527.625 -46.565 530.955 ;
        RECT -33.035 530.770 -32.730 532.315 ;
        RECT -33.035 530.480 -32.590 530.770 ;
        RECT -30.620 530.480 -28.090 575.460 ;
        RECT -33.035 530.370 -28.090 530.480 ;
        RECT -42.750 527.950 -42.320 529.175 ;
        RECT -33.020 528.920 -28.090 530.370 ;
        RECT -34.745 528.780 -28.090 528.920 ;
        RECT -34.745 528.750 -32.590 528.780 ;
        RECT -33.205 528.745 -32.590 528.750 ;
        RECT -42.750 527.780 -41.540 527.950 ;
        RECT -33.020 527.875 -32.590 528.745 ;
        RECT -42.750 527.625 -42.320 527.780 ;
        RECT -60.015 526.760 -58.805 526.930 ;
        RECT -60.015 526.060 -59.585 526.760 ;
        RECT -62.445 525.335 -62.050 525.370 ;
        RECT -62.445 523.885 -62.140 525.335 ;
        RECT -51.120 524.995 -50.690 527.405 ;
        RECT -47.130 527.320 -42.320 527.625 ;
        RECT -45.090 525.410 -44.785 527.320 ;
        RECT -42.750 526.970 -42.320 527.320 ;
        RECT -33.855 527.445 -32.590 527.875 ;
        RECT -42.750 526.800 -41.540 526.970 ;
        RECT -42.750 526.100 -42.320 526.800 ;
        RECT -52.400 524.825 -50.690 524.995 ;
        RECT -51.120 524.015 -50.690 524.825 ;
        RECT -62.445 523.715 -60.340 523.885 ;
        RECT -52.400 523.845 -50.690 524.015 ;
        RECT -62.445 523.710 -61.880 523.715 ;
        RECT -62.445 523.125 -62.140 523.710 ;
        RECT -59.680 522.800 -59.410 523.475 ;
        RECT -51.120 523.145 -50.690 523.845 ;
        RECT -45.180 525.375 -44.785 525.410 ;
        RECT -45.180 523.925 -44.875 525.375 ;
        RECT -33.855 525.035 -33.425 527.445 ;
        RECT -35.135 524.865 -33.425 525.035 ;
        RECT -33.855 524.055 -33.425 524.865 ;
        RECT -45.180 523.755 -43.075 523.925 ;
        RECT -35.135 523.885 -33.425 524.055 ;
        RECT -45.180 523.750 -44.615 523.755 ;
        RECT -45.180 523.165 -44.875 523.750 ;
        RECT -33.855 523.185 -33.425 523.885 ;
        RECT -59.640 522.700 -59.440 522.800 ;
        RECT -59.630 521.655 -59.450 522.700 ;
        RECT -78.950 520.975 -59.450 521.655 ;
        RECT -78.950 42.775 -78.270 520.975 ;
        RECT -59.630 520.060 -59.450 520.975 ;
        RECT -64.635 505.915 -64.070 507.240 ;
        RECT -64.635 505.885 -63.425 505.915 ;
        RECT -64.635 505.715 -62.010 505.885 ;
        RECT -64.635 505.680 -63.425 505.715 ;
        RECT -64.635 504.705 -64.070 505.680 ;
        RECT -53.005 505.480 -52.575 507.555 ;
        RECT -53.785 505.310 -52.575 505.480 ;
        RECT -53.005 505.155 -52.575 505.310 ;
        RECT -53.005 504.850 -50.235 505.155 ;
        RECT -64.635 504.675 -63.475 504.705 ;
        RECT -64.635 504.505 -62.010 504.675 ;
        RECT -64.635 504.470 -63.475 504.505 ;
        RECT -53.005 504.500 -52.575 504.850 ;
        RECT -64.635 503.725 -64.070 504.470 ;
        RECT -53.785 504.330 -52.575 504.500 ;
        RECT -64.635 503.695 -63.480 503.725 ;
        RECT -64.635 503.525 -62.010 503.695 ;
        RECT -53.005 503.630 -52.575 504.330 ;
        RECT -64.635 503.490 -63.480 503.525 ;
        RECT -64.635 500.160 -64.070 503.490 ;
        RECT -50.540 503.305 -50.235 504.850 ;
        RECT -50.540 502.905 -50.095 503.305 ;
        RECT -60.255 500.485 -59.825 501.710 ;
        RECT -50.525 501.455 -50.095 502.905 ;
        RECT -52.250 501.285 -50.095 501.455 ;
        RECT -50.710 501.280 -50.095 501.285 ;
        RECT -60.255 500.315 -59.045 500.485 ;
        RECT -50.525 500.410 -50.095 501.280 ;
        RECT -60.255 500.160 -59.825 500.315 ;
        RECT -64.635 499.855 -59.825 500.160 ;
        RECT -62.595 497.945 -62.290 499.855 ;
        RECT -60.255 499.505 -59.825 499.855 ;
        RECT -51.360 499.980 -50.095 500.410 ;
        RECT -47.135 501.105 -46.330 501.670 ;
        RECT -47.135 501.100 -45.745 501.105 ;
        RECT -47.135 500.930 -44.300 501.100 ;
        RECT -47.135 500.920 -45.745 500.930 ;
        RECT -60.255 499.335 -59.045 499.505 ;
        RECT -60.255 498.635 -59.825 499.335 ;
        RECT -62.685 497.910 -62.290 497.945 ;
        RECT -62.685 496.460 -62.380 497.910 ;
        RECT -51.360 497.570 -50.930 499.980 ;
        RECT -52.640 497.400 -50.930 497.570 ;
        RECT -51.360 496.590 -50.930 497.400 ;
        RECT -62.685 496.290 -60.580 496.460 ;
        RECT -52.640 496.420 -50.930 496.590 ;
        RECT -62.685 496.285 -62.120 496.290 ;
        RECT -62.685 495.700 -62.380 496.285 ;
        RECT -59.920 495.375 -59.650 496.050 ;
        RECT -51.360 495.720 -50.930 496.420 ;
        RECT -47.135 499.470 -46.330 500.920 ;
        RECT -47.135 499.300 -43.300 499.470 ;
        RECT -47.135 499.285 -45.750 499.300 ;
        RECT -47.135 498.830 -46.330 499.285 ;
        RECT -47.135 498.820 -45.755 498.830 ;
        RECT -47.135 498.650 -43.300 498.820 ;
        RECT -47.135 498.645 -45.755 498.650 ;
        RECT -59.880 495.275 -59.680 495.375 ;
        RECT -59.870 493.885 -59.690 495.275 ;
        RECT -47.135 495.055 -46.330 498.645 ;
        RECT -47.135 494.870 -46.310 495.055 ;
        RECT -47.135 494.865 -45.755 494.870 ;
        RECT -47.135 494.695 -44.300 494.865 ;
        RECT -47.135 494.685 -45.755 494.695 ;
        RECT -47.135 494.305 -46.310 494.685 ;
        RECT -65.530 493.205 -59.690 493.885 ;
        RECT -65.530 475.890 -64.850 493.205 ;
        RECT -46.875 492.565 -46.310 494.305 ;
        RECT -47.215 492.000 -46.310 492.565 ;
        RECT -64.480 487.575 -63.915 488.900 ;
        RECT -64.480 487.545 -63.270 487.575 ;
        RECT -64.480 487.375 -61.855 487.545 ;
        RECT -64.480 487.340 -63.270 487.375 ;
        RECT -64.480 486.365 -63.915 487.340 ;
        RECT -52.850 487.140 -52.420 489.215 ;
        RECT -53.630 486.970 -52.420 487.140 ;
        RECT -52.850 486.815 -52.420 486.970 ;
        RECT -47.215 487.615 -46.650 492.000 ;
        RECT -47.215 487.585 -46.005 487.615 ;
        RECT -47.215 487.415 -44.590 487.585 ;
        RECT -47.215 487.380 -46.005 487.415 ;
        RECT -52.850 486.510 -50.080 486.815 ;
        RECT -64.480 486.335 -63.320 486.365 ;
        RECT -64.480 486.165 -61.855 486.335 ;
        RECT -64.480 486.130 -63.320 486.165 ;
        RECT -52.850 486.160 -52.420 486.510 ;
        RECT -64.480 485.385 -63.915 486.130 ;
        RECT -53.630 485.990 -52.420 486.160 ;
        RECT -64.480 485.355 -63.325 485.385 ;
        RECT -64.480 485.185 -61.855 485.355 ;
        RECT -52.850 485.290 -52.420 485.990 ;
        RECT -64.480 485.150 -63.325 485.185 ;
        RECT -64.480 481.820 -63.915 485.150 ;
        RECT -50.385 484.965 -50.080 486.510 ;
        RECT -47.215 486.405 -46.650 487.380 ;
        RECT -35.585 487.180 -35.155 489.255 ;
        RECT -36.365 487.010 -35.155 487.180 ;
        RECT -35.585 486.855 -35.155 487.010 ;
        RECT -35.585 486.550 -32.815 486.855 ;
        RECT -47.215 486.375 -46.055 486.405 ;
        RECT -47.215 486.205 -44.590 486.375 ;
        RECT -47.215 486.170 -46.055 486.205 ;
        RECT -35.585 486.200 -35.155 486.550 ;
        RECT -47.215 485.425 -46.650 486.170 ;
        RECT -36.365 486.030 -35.155 486.200 ;
        RECT -47.215 485.395 -46.060 485.425 ;
        RECT -47.215 485.225 -44.590 485.395 ;
        RECT -35.585 485.330 -35.155 486.030 ;
        RECT -47.215 485.190 -46.060 485.225 ;
        RECT -50.385 484.565 -49.940 484.965 ;
        RECT -60.100 482.145 -59.670 483.370 ;
        RECT -50.370 483.115 -49.940 484.565 ;
        RECT -52.095 482.945 -49.940 483.115 ;
        RECT -50.555 482.940 -49.940 482.945 ;
        RECT -60.100 481.975 -58.890 482.145 ;
        RECT -50.370 482.070 -49.940 482.940 ;
        RECT -60.100 481.820 -59.670 481.975 ;
        RECT -64.480 481.515 -59.670 481.820 ;
        RECT -62.440 479.605 -62.135 481.515 ;
        RECT -60.100 481.165 -59.670 481.515 ;
        RECT -51.205 481.640 -49.940 482.070 ;
        RECT -47.215 481.860 -46.650 485.190 ;
        RECT -33.120 485.005 -32.815 486.550 ;
        RECT -33.120 484.785 -32.675 485.005 ;
        RECT -30.620 484.785 -28.090 528.780 ;
        RECT -33.120 484.605 -28.090 484.785 ;
        RECT -42.835 482.185 -42.405 483.410 ;
        RECT -33.105 483.250 -28.090 484.605 ;
        RECT -33.105 483.155 -32.675 483.250 ;
        RECT -34.830 482.985 -32.675 483.155 ;
        RECT -33.290 482.980 -32.675 482.985 ;
        RECT -42.835 482.015 -41.625 482.185 ;
        RECT -33.105 482.110 -32.675 482.980 ;
        RECT -42.835 481.860 -42.405 482.015 ;
        RECT -60.100 480.995 -58.890 481.165 ;
        RECT -60.100 480.295 -59.670 480.995 ;
        RECT -62.530 479.570 -62.135 479.605 ;
        RECT -62.530 478.120 -62.225 479.570 ;
        RECT -51.205 479.230 -50.775 481.640 ;
        RECT -47.215 481.555 -42.405 481.860 ;
        RECT -45.175 479.645 -44.870 481.555 ;
        RECT -42.835 481.205 -42.405 481.555 ;
        RECT -33.940 481.680 -32.675 482.110 ;
        RECT -42.835 481.035 -41.625 481.205 ;
        RECT -42.835 480.335 -42.405 481.035 ;
        RECT -52.485 479.060 -50.775 479.230 ;
        RECT -51.205 478.250 -50.775 479.060 ;
        RECT -62.530 477.950 -60.425 478.120 ;
        RECT -52.485 478.080 -50.775 478.250 ;
        RECT -62.530 477.945 -61.965 477.950 ;
        RECT -62.530 477.360 -62.225 477.945 ;
        RECT -59.765 477.035 -59.495 477.710 ;
        RECT -51.205 477.380 -50.775 478.080 ;
        RECT -45.265 479.610 -44.870 479.645 ;
        RECT -45.265 478.160 -44.960 479.610 ;
        RECT -33.940 479.270 -33.510 481.680 ;
        RECT -35.220 479.100 -33.510 479.270 ;
        RECT -33.940 478.290 -33.510 479.100 ;
        RECT -45.265 477.990 -43.160 478.160 ;
        RECT -35.220 478.120 -33.510 478.290 ;
        RECT -45.265 477.985 -44.700 477.990 ;
        RECT -45.265 477.400 -44.960 477.985 ;
        RECT -33.940 477.420 -33.510 478.120 ;
        RECT -59.725 476.935 -59.525 477.035 ;
        RECT -59.715 475.890 -59.535 476.935 ;
        RECT -77.455 475.210 -59.535 475.890 ;
        RECT -77.455 208.690 -76.775 475.210 ;
        RECT -59.715 474.295 -59.535 475.210 ;
        RECT -64.965 462.145 -64.400 463.470 ;
        RECT -64.965 462.115 -63.755 462.145 ;
        RECT -64.965 461.945 -62.340 462.115 ;
        RECT -64.965 461.910 -63.755 461.945 ;
        RECT -64.965 460.935 -64.400 461.910 ;
        RECT -53.335 461.710 -52.905 463.785 ;
        RECT -54.115 461.540 -52.905 461.710 ;
        RECT -53.335 461.385 -52.905 461.540 ;
        RECT -53.335 461.080 -50.565 461.385 ;
        RECT -64.965 460.905 -63.805 460.935 ;
        RECT -64.965 460.735 -62.340 460.905 ;
        RECT -64.965 460.700 -63.805 460.735 ;
        RECT -53.335 460.730 -52.905 461.080 ;
        RECT -64.965 459.955 -64.400 460.700 ;
        RECT -54.115 460.560 -52.905 460.730 ;
        RECT -64.965 459.925 -63.810 459.955 ;
        RECT -64.965 459.755 -62.340 459.925 ;
        RECT -53.335 459.860 -52.905 460.560 ;
        RECT -64.965 459.720 -63.810 459.755 ;
        RECT -64.965 456.390 -64.400 459.720 ;
        RECT -50.870 459.535 -50.565 461.080 ;
        RECT -50.870 459.135 -50.425 459.535 ;
        RECT -60.585 456.715 -60.155 457.940 ;
        RECT -50.855 457.685 -50.425 459.135 ;
        RECT -52.580 457.515 -50.425 457.685 ;
        RECT -51.040 457.510 -50.425 457.515 ;
        RECT -60.585 456.545 -59.375 456.715 ;
        RECT -50.855 456.640 -50.425 457.510 ;
        RECT -60.585 456.390 -60.155 456.545 ;
        RECT -64.965 456.085 -60.155 456.390 ;
        RECT -62.925 454.175 -62.620 456.085 ;
        RECT -60.585 455.735 -60.155 456.085 ;
        RECT -51.690 456.210 -50.425 456.640 ;
        RECT -47.465 457.335 -46.660 457.900 ;
        RECT -47.465 457.330 -46.075 457.335 ;
        RECT -47.465 457.160 -44.630 457.330 ;
        RECT -47.465 457.150 -46.075 457.160 ;
        RECT -60.585 455.565 -59.375 455.735 ;
        RECT -60.585 454.865 -60.155 455.565 ;
        RECT -63.015 454.140 -62.620 454.175 ;
        RECT -63.015 452.690 -62.710 454.140 ;
        RECT -51.690 453.800 -51.260 456.210 ;
        RECT -52.970 453.630 -51.260 453.800 ;
        RECT -51.690 452.820 -51.260 453.630 ;
        RECT -63.015 452.520 -60.910 452.690 ;
        RECT -52.970 452.650 -51.260 452.820 ;
        RECT -63.015 452.515 -62.450 452.520 ;
        RECT -63.015 451.930 -62.710 452.515 ;
        RECT -51.690 451.950 -51.260 452.650 ;
        RECT -47.465 455.700 -46.660 457.150 ;
        RECT -47.465 455.530 -43.630 455.700 ;
        RECT -47.465 455.515 -46.080 455.530 ;
        RECT -47.465 455.060 -46.660 455.515 ;
        RECT -47.465 455.050 -46.085 455.060 ;
        RECT -47.465 454.880 -43.630 455.050 ;
        RECT -47.465 454.875 -46.085 454.880 ;
        RECT -47.465 451.285 -46.660 454.875 ;
        RECT -47.465 451.100 -46.640 451.285 ;
        RECT -47.465 451.095 -46.085 451.100 ;
        RECT -47.465 450.925 -44.630 451.095 ;
        RECT -47.465 450.915 -46.085 450.925 ;
        RECT -47.465 450.535 -46.640 450.915 ;
        RECT -47.205 448.795 -46.640 450.535 ;
        RECT -47.545 448.230 -46.640 448.795 ;
        RECT -64.810 443.805 -64.245 445.130 ;
        RECT -64.810 443.775 -63.600 443.805 ;
        RECT -64.810 443.605 -62.185 443.775 ;
        RECT -64.810 443.570 -63.600 443.605 ;
        RECT -64.810 442.595 -64.245 443.570 ;
        RECT -53.180 443.370 -52.750 445.445 ;
        RECT -53.960 443.200 -52.750 443.370 ;
        RECT -53.180 443.045 -52.750 443.200 ;
        RECT -47.545 443.845 -46.980 448.230 ;
        RECT -47.545 443.815 -46.335 443.845 ;
        RECT -47.545 443.645 -44.920 443.815 ;
        RECT -47.545 443.610 -46.335 443.645 ;
        RECT -53.180 442.740 -50.410 443.045 ;
        RECT -64.810 442.565 -63.650 442.595 ;
        RECT -64.810 442.395 -62.185 442.565 ;
        RECT -64.810 442.360 -63.650 442.395 ;
        RECT -53.180 442.390 -52.750 442.740 ;
        RECT -64.810 441.615 -64.245 442.360 ;
        RECT -53.960 442.220 -52.750 442.390 ;
        RECT -64.810 441.585 -63.655 441.615 ;
        RECT -64.810 441.415 -62.185 441.585 ;
        RECT -53.180 441.520 -52.750 442.220 ;
        RECT -64.810 441.380 -63.655 441.415 ;
        RECT -64.810 438.050 -64.245 441.380 ;
        RECT -50.715 441.195 -50.410 442.740 ;
        RECT -47.545 442.635 -46.980 443.610 ;
        RECT -35.915 443.410 -35.485 445.485 ;
        RECT -36.695 443.240 -35.485 443.410 ;
        RECT -35.915 443.085 -35.485 443.240 ;
        RECT -35.915 442.780 -33.145 443.085 ;
        RECT -47.545 442.605 -46.385 442.635 ;
        RECT -47.545 442.435 -44.920 442.605 ;
        RECT -47.545 442.400 -46.385 442.435 ;
        RECT -35.915 442.430 -35.485 442.780 ;
        RECT -47.545 441.655 -46.980 442.400 ;
        RECT -36.695 442.260 -35.485 442.430 ;
        RECT -47.545 441.625 -46.390 441.655 ;
        RECT -47.545 441.455 -44.920 441.625 ;
        RECT -35.915 441.560 -35.485 442.260 ;
        RECT -47.545 441.420 -46.390 441.455 ;
        RECT -50.715 440.795 -50.270 441.195 ;
        RECT -60.430 438.375 -60.000 439.600 ;
        RECT -50.700 439.345 -50.270 440.795 ;
        RECT -52.425 439.175 -50.270 439.345 ;
        RECT -50.885 439.170 -50.270 439.175 ;
        RECT -60.430 438.205 -59.220 438.375 ;
        RECT -50.700 438.300 -50.270 439.170 ;
        RECT -60.430 438.050 -60.000 438.205 ;
        RECT -64.810 437.745 -60.000 438.050 ;
        RECT -62.770 435.835 -62.465 437.745 ;
        RECT -60.430 437.395 -60.000 437.745 ;
        RECT -51.535 437.870 -50.270 438.300 ;
        RECT -47.545 438.090 -46.980 441.420 ;
        RECT -33.450 441.235 -33.145 442.780 ;
        RECT -33.450 440.835 -33.005 441.235 ;
        RECT -33.435 440.690 -33.005 440.835 ;
        RECT -30.620 440.690 -28.090 483.250 ;
        RECT -43.165 438.415 -42.735 439.640 ;
        RECT -33.435 439.385 -28.090 440.690 ;
        RECT -35.160 439.275 -28.090 439.385 ;
        RECT -35.160 439.215 -33.005 439.275 ;
        RECT -33.620 439.210 -33.005 439.215 ;
        RECT -43.165 438.245 -41.955 438.415 ;
        RECT -33.435 438.340 -33.005 439.210 ;
        RECT -43.165 438.090 -42.735 438.245 ;
        RECT -60.430 437.225 -59.220 437.395 ;
        RECT -60.430 436.525 -60.000 437.225 ;
        RECT -62.860 435.800 -62.465 435.835 ;
        RECT -62.860 434.350 -62.555 435.800 ;
        RECT -51.535 435.460 -51.105 437.870 ;
        RECT -47.545 437.785 -42.735 438.090 ;
        RECT -45.505 435.875 -45.200 437.785 ;
        RECT -43.165 437.435 -42.735 437.785 ;
        RECT -34.270 437.910 -33.005 438.340 ;
        RECT -43.165 437.265 -41.955 437.435 ;
        RECT -43.165 436.565 -42.735 437.265 ;
        RECT -52.815 435.290 -51.105 435.460 ;
        RECT -51.535 434.480 -51.105 435.290 ;
        RECT -62.860 434.180 -60.755 434.350 ;
        RECT -52.815 434.310 -51.105 434.480 ;
        RECT -62.860 434.175 -62.295 434.180 ;
        RECT -62.860 433.590 -62.555 434.175 ;
        RECT -51.535 433.610 -51.105 434.310 ;
        RECT -45.595 435.840 -45.200 435.875 ;
        RECT -45.595 434.390 -45.290 435.840 ;
        RECT -34.270 435.500 -33.840 437.910 ;
        RECT -35.550 435.330 -33.840 435.500 ;
        RECT -34.270 434.520 -33.840 435.330 ;
        RECT -45.595 434.220 -43.490 434.390 ;
        RECT -35.550 434.350 -33.840 434.520 ;
        RECT -45.595 434.215 -45.030 434.220 ;
        RECT -45.595 433.630 -45.290 434.215 ;
        RECT -34.270 433.650 -33.840 434.350 ;
        RECT -65.135 416.155 -64.570 417.480 ;
        RECT -65.135 416.125 -63.925 416.155 ;
        RECT -65.135 415.955 -62.510 416.125 ;
        RECT -65.135 415.920 -63.925 415.955 ;
        RECT -65.135 414.945 -64.570 415.920 ;
        RECT -53.505 415.720 -53.075 417.795 ;
        RECT -54.285 415.550 -53.075 415.720 ;
        RECT -53.505 415.395 -53.075 415.550 ;
        RECT -53.505 415.090 -50.735 415.395 ;
        RECT -65.135 414.915 -63.975 414.945 ;
        RECT -65.135 414.745 -62.510 414.915 ;
        RECT -65.135 414.710 -63.975 414.745 ;
        RECT -53.505 414.740 -53.075 415.090 ;
        RECT -65.135 413.965 -64.570 414.710 ;
        RECT -54.285 414.570 -53.075 414.740 ;
        RECT -65.135 413.935 -63.980 413.965 ;
        RECT -65.135 413.765 -62.510 413.935 ;
        RECT -53.505 413.870 -53.075 414.570 ;
        RECT -65.135 413.730 -63.980 413.765 ;
        RECT -65.135 410.400 -64.570 413.730 ;
        RECT -51.040 413.545 -50.735 415.090 ;
        RECT -51.040 413.145 -50.595 413.545 ;
        RECT -60.755 410.725 -60.325 411.950 ;
        RECT -51.025 411.695 -50.595 413.145 ;
        RECT -52.750 411.525 -50.595 411.695 ;
        RECT -51.210 411.520 -50.595 411.525 ;
        RECT -60.755 410.555 -59.545 410.725 ;
        RECT -51.025 410.650 -50.595 411.520 ;
        RECT -60.755 410.400 -60.325 410.555 ;
        RECT -65.135 410.095 -60.325 410.400 ;
        RECT -63.095 408.185 -62.790 410.095 ;
        RECT -60.755 409.745 -60.325 410.095 ;
        RECT -51.860 410.220 -50.595 410.650 ;
        RECT -47.635 411.345 -46.830 411.910 ;
        RECT -47.635 411.340 -46.245 411.345 ;
        RECT -47.635 411.170 -44.800 411.340 ;
        RECT -47.635 411.160 -46.245 411.170 ;
        RECT -60.755 409.575 -59.545 409.745 ;
        RECT -60.755 408.875 -60.325 409.575 ;
        RECT -63.185 408.150 -62.790 408.185 ;
        RECT -63.185 406.700 -62.880 408.150 ;
        RECT -51.860 407.810 -51.430 410.220 ;
        RECT -53.140 407.640 -51.430 407.810 ;
        RECT -51.860 406.830 -51.430 407.640 ;
        RECT -63.185 406.530 -61.080 406.700 ;
        RECT -53.140 406.660 -51.430 406.830 ;
        RECT -63.185 406.525 -62.620 406.530 ;
        RECT -63.185 405.940 -62.880 406.525 ;
        RECT -51.860 405.960 -51.430 406.660 ;
        RECT -47.635 409.710 -46.830 411.160 ;
        RECT -47.635 409.540 -43.800 409.710 ;
        RECT -47.635 409.525 -46.250 409.540 ;
        RECT -47.635 409.070 -46.830 409.525 ;
        RECT -47.635 409.060 -46.255 409.070 ;
        RECT -47.635 408.890 -43.800 409.060 ;
        RECT -47.635 408.885 -46.255 408.890 ;
        RECT -47.635 405.295 -46.830 408.885 ;
        RECT -47.635 405.110 -46.810 405.295 ;
        RECT -47.635 405.105 -46.255 405.110 ;
        RECT -47.635 404.935 -44.800 405.105 ;
        RECT -47.635 404.925 -46.255 404.935 ;
        RECT -47.635 404.545 -46.810 404.925 ;
        RECT -47.375 402.805 -46.810 404.545 ;
        RECT -47.715 402.240 -46.810 402.805 ;
        RECT -64.980 397.815 -64.415 399.140 ;
        RECT -64.980 397.785 -63.770 397.815 ;
        RECT -64.980 397.615 -62.355 397.785 ;
        RECT -64.980 397.580 -63.770 397.615 ;
        RECT -64.980 396.605 -64.415 397.580 ;
        RECT -53.350 397.380 -52.920 399.455 ;
        RECT -54.130 397.210 -52.920 397.380 ;
        RECT -53.350 397.055 -52.920 397.210 ;
        RECT -47.715 397.855 -47.150 402.240 ;
        RECT -47.715 397.825 -46.505 397.855 ;
        RECT -47.715 397.655 -45.090 397.825 ;
        RECT -47.715 397.620 -46.505 397.655 ;
        RECT -53.350 396.750 -50.580 397.055 ;
        RECT -64.980 396.575 -63.820 396.605 ;
        RECT -64.980 396.405 -62.355 396.575 ;
        RECT -64.980 396.370 -63.820 396.405 ;
        RECT -53.350 396.400 -52.920 396.750 ;
        RECT -64.980 395.625 -64.415 396.370 ;
        RECT -54.130 396.230 -52.920 396.400 ;
        RECT -64.980 395.595 -63.825 395.625 ;
        RECT -64.980 395.425 -62.355 395.595 ;
        RECT -53.350 395.530 -52.920 396.230 ;
        RECT -64.980 395.390 -63.825 395.425 ;
        RECT -64.980 392.060 -64.415 395.390 ;
        RECT -50.885 395.205 -50.580 396.750 ;
        RECT -47.715 396.645 -47.150 397.620 ;
        RECT -36.085 397.420 -35.655 399.495 ;
        RECT -36.865 397.250 -35.655 397.420 ;
        RECT -36.085 397.095 -35.655 397.250 ;
        RECT -36.085 396.790 -33.315 397.095 ;
        RECT -47.715 396.615 -46.555 396.645 ;
        RECT -47.715 396.445 -45.090 396.615 ;
        RECT -47.715 396.410 -46.555 396.445 ;
        RECT -36.085 396.440 -35.655 396.790 ;
        RECT -47.715 395.665 -47.150 396.410 ;
        RECT -36.865 396.270 -35.655 396.440 ;
        RECT -47.715 395.635 -46.560 395.665 ;
        RECT -47.715 395.465 -45.090 395.635 ;
        RECT -36.085 395.570 -35.655 396.270 ;
        RECT -47.715 395.430 -46.560 395.465 ;
        RECT -50.885 394.805 -50.440 395.205 ;
        RECT -60.600 392.385 -60.170 393.610 ;
        RECT -50.870 393.355 -50.440 394.805 ;
        RECT -52.595 393.185 -50.440 393.355 ;
        RECT -51.055 393.180 -50.440 393.185 ;
        RECT -60.600 392.215 -59.390 392.385 ;
        RECT -50.870 392.310 -50.440 393.180 ;
        RECT -60.600 392.060 -60.170 392.215 ;
        RECT -64.980 391.755 -60.170 392.060 ;
        RECT -62.940 389.845 -62.635 391.755 ;
        RECT -60.600 391.405 -60.170 391.755 ;
        RECT -51.705 391.880 -50.440 392.310 ;
        RECT -47.715 392.100 -47.150 395.430 ;
        RECT -33.620 395.245 -33.315 396.790 ;
        RECT -33.620 394.845 -33.175 395.245 ;
        RECT -33.605 394.595 -33.175 394.845 ;
        RECT -30.620 394.595 -28.090 439.275 ;
        RECT -43.335 392.425 -42.905 393.650 ;
        RECT -33.605 393.395 -28.090 394.595 ;
        RECT -35.330 393.225 -28.090 393.395 ;
        RECT -33.790 393.220 -28.090 393.225 ;
        RECT -33.605 393.180 -28.090 393.220 ;
        RECT -43.335 392.255 -42.125 392.425 ;
        RECT -33.605 392.350 -33.175 393.180 ;
        RECT -43.335 392.100 -42.905 392.255 ;
        RECT -60.600 391.235 -59.390 391.405 ;
        RECT -60.600 390.535 -60.170 391.235 ;
        RECT -63.030 389.810 -62.635 389.845 ;
        RECT -63.030 388.360 -62.725 389.810 ;
        RECT -51.705 389.470 -51.275 391.880 ;
        RECT -47.715 391.795 -42.905 392.100 ;
        RECT -45.675 389.885 -45.370 391.795 ;
        RECT -43.335 391.445 -42.905 391.795 ;
        RECT -34.440 391.920 -33.175 392.350 ;
        RECT -43.335 391.275 -42.125 391.445 ;
        RECT -43.335 390.575 -42.905 391.275 ;
        RECT -52.985 389.300 -51.275 389.470 ;
        RECT -51.705 388.490 -51.275 389.300 ;
        RECT -63.030 388.190 -60.925 388.360 ;
        RECT -52.985 388.320 -51.275 388.490 ;
        RECT -63.030 388.185 -62.465 388.190 ;
        RECT -63.030 387.600 -62.725 388.185 ;
        RECT -51.705 387.620 -51.275 388.320 ;
        RECT -45.765 389.850 -45.370 389.885 ;
        RECT -45.765 388.400 -45.460 389.850 ;
        RECT -34.440 389.510 -34.010 391.920 ;
        RECT -35.720 389.340 -34.010 389.510 ;
        RECT -34.440 388.530 -34.010 389.340 ;
        RECT -45.765 388.230 -43.660 388.400 ;
        RECT -35.720 388.360 -34.010 388.530 ;
        RECT -45.765 388.225 -45.200 388.230 ;
        RECT -45.765 387.640 -45.460 388.225 ;
        RECT -34.440 387.660 -34.010 388.360 ;
        RECT -64.940 371.840 -64.375 373.165 ;
        RECT -64.940 371.810 -63.730 371.840 ;
        RECT -64.940 371.640 -62.315 371.810 ;
        RECT -64.940 371.605 -63.730 371.640 ;
        RECT -64.940 370.630 -64.375 371.605 ;
        RECT -53.310 371.405 -52.880 373.480 ;
        RECT -54.090 371.235 -52.880 371.405 ;
        RECT -53.310 371.080 -52.880 371.235 ;
        RECT -53.310 370.775 -50.540 371.080 ;
        RECT -64.940 370.600 -63.780 370.630 ;
        RECT -64.940 370.430 -62.315 370.600 ;
        RECT -64.940 370.395 -63.780 370.430 ;
        RECT -53.310 370.425 -52.880 370.775 ;
        RECT -64.940 369.650 -64.375 370.395 ;
        RECT -54.090 370.255 -52.880 370.425 ;
        RECT -64.940 369.620 -63.785 369.650 ;
        RECT -64.940 369.450 -62.315 369.620 ;
        RECT -53.310 369.555 -52.880 370.255 ;
        RECT -64.940 369.415 -63.785 369.450 ;
        RECT -64.940 366.085 -64.375 369.415 ;
        RECT -50.845 369.230 -50.540 370.775 ;
        RECT -50.845 368.830 -50.400 369.230 ;
        RECT -60.560 366.410 -60.130 367.635 ;
        RECT -50.830 367.380 -50.400 368.830 ;
        RECT -52.555 367.210 -50.400 367.380 ;
        RECT -51.015 367.205 -50.400 367.210 ;
        RECT -60.560 366.240 -59.350 366.410 ;
        RECT -50.830 366.335 -50.400 367.205 ;
        RECT -60.560 366.085 -60.130 366.240 ;
        RECT -64.940 365.780 -60.130 366.085 ;
        RECT -62.900 363.870 -62.595 365.780 ;
        RECT -60.560 365.430 -60.130 365.780 ;
        RECT -51.665 365.905 -50.400 366.335 ;
        RECT -47.440 367.030 -46.635 367.595 ;
        RECT -47.440 367.025 -46.050 367.030 ;
        RECT -47.440 366.855 -44.605 367.025 ;
        RECT -47.440 366.845 -46.050 366.855 ;
        RECT -60.560 365.260 -59.350 365.430 ;
        RECT -60.560 364.560 -60.130 365.260 ;
        RECT -62.990 363.835 -62.595 363.870 ;
        RECT -62.990 362.385 -62.685 363.835 ;
        RECT -51.665 363.495 -51.235 365.905 ;
        RECT -52.945 363.325 -51.235 363.495 ;
        RECT -51.665 362.515 -51.235 363.325 ;
        RECT -62.990 362.215 -60.885 362.385 ;
        RECT -52.945 362.345 -51.235 362.515 ;
        RECT -62.990 362.210 -62.425 362.215 ;
        RECT -62.990 361.625 -62.685 362.210 ;
        RECT -51.665 361.645 -51.235 362.345 ;
        RECT -47.440 365.395 -46.635 366.845 ;
        RECT -47.440 365.225 -43.605 365.395 ;
        RECT -47.440 365.210 -46.055 365.225 ;
        RECT -47.440 364.755 -46.635 365.210 ;
        RECT -47.440 364.745 -46.060 364.755 ;
        RECT -47.440 364.575 -43.605 364.745 ;
        RECT -47.440 364.570 -46.060 364.575 ;
        RECT -47.440 360.980 -46.635 364.570 ;
        RECT -47.440 360.795 -46.615 360.980 ;
        RECT -47.440 360.790 -46.060 360.795 ;
        RECT -47.440 360.620 -44.605 360.790 ;
        RECT -47.440 360.610 -46.060 360.620 ;
        RECT -47.440 360.230 -46.615 360.610 ;
        RECT -47.180 358.490 -46.615 360.230 ;
        RECT -47.520 357.925 -46.615 358.490 ;
        RECT -64.785 353.500 -64.220 354.825 ;
        RECT -64.785 353.470 -63.575 353.500 ;
        RECT -64.785 353.300 -62.160 353.470 ;
        RECT -64.785 353.265 -63.575 353.300 ;
        RECT -64.785 352.290 -64.220 353.265 ;
        RECT -53.155 353.065 -52.725 355.140 ;
        RECT -53.935 352.895 -52.725 353.065 ;
        RECT -53.155 352.740 -52.725 352.895 ;
        RECT -47.520 353.540 -46.955 357.925 ;
        RECT -47.520 353.510 -46.310 353.540 ;
        RECT -47.520 353.340 -44.895 353.510 ;
        RECT -47.520 353.305 -46.310 353.340 ;
        RECT -53.155 352.435 -50.385 352.740 ;
        RECT -64.785 352.260 -63.625 352.290 ;
        RECT -64.785 352.090 -62.160 352.260 ;
        RECT -64.785 352.055 -63.625 352.090 ;
        RECT -53.155 352.085 -52.725 352.435 ;
        RECT -64.785 351.310 -64.220 352.055 ;
        RECT -53.935 351.915 -52.725 352.085 ;
        RECT -64.785 351.280 -63.630 351.310 ;
        RECT -64.785 351.110 -62.160 351.280 ;
        RECT -53.155 351.215 -52.725 351.915 ;
        RECT -64.785 351.075 -63.630 351.110 ;
        RECT -64.785 347.745 -64.220 351.075 ;
        RECT -50.690 350.890 -50.385 352.435 ;
        RECT -47.520 352.330 -46.955 353.305 ;
        RECT -35.890 353.105 -35.460 355.180 ;
        RECT -36.670 352.935 -35.460 353.105 ;
        RECT -35.890 352.780 -35.460 352.935 ;
        RECT -35.890 352.475 -33.120 352.780 ;
        RECT -47.520 352.300 -46.360 352.330 ;
        RECT -47.520 352.130 -44.895 352.300 ;
        RECT -47.520 352.095 -46.360 352.130 ;
        RECT -35.890 352.125 -35.460 352.475 ;
        RECT -47.520 351.350 -46.955 352.095 ;
        RECT -36.670 351.955 -35.460 352.125 ;
        RECT -47.520 351.320 -46.365 351.350 ;
        RECT -47.520 351.150 -44.895 351.320 ;
        RECT -35.890 351.255 -35.460 351.955 ;
        RECT -47.520 351.115 -46.365 351.150 ;
        RECT -50.690 350.490 -50.245 350.890 ;
        RECT -60.405 348.070 -59.975 349.295 ;
        RECT -50.675 349.040 -50.245 350.490 ;
        RECT -52.400 348.870 -50.245 349.040 ;
        RECT -50.860 348.865 -50.245 348.870 ;
        RECT -60.405 347.900 -59.195 348.070 ;
        RECT -50.675 347.995 -50.245 348.865 ;
        RECT -60.405 347.745 -59.975 347.900 ;
        RECT -64.785 347.440 -59.975 347.745 ;
        RECT -62.745 345.530 -62.440 347.440 ;
        RECT -60.405 347.090 -59.975 347.440 ;
        RECT -51.510 347.565 -50.245 347.995 ;
        RECT -47.520 347.785 -46.955 351.115 ;
        RECT -33.425 350.930 -33.120 352.475 ;
        RECT -33.425 350.530 -32.980 350.930 ;
        RECT -33.410 350.035 -32.980 350.530 ;
        RECT -30.620 350.035 -28.090 393.180 ;
        RECT -43.140 348.110 -42.710 349.335 ;
        RECT -33.410 349.080 -28.090 350.035 ;
        RECT -35.135 348.910 -28.090 349.080 ;
        RECT -33.595 348.905 -28.090 348.910 ;
        RECT -33.410 348.620 -28.090 348.905 ;
        RECT -43.140 347.940 -41.930 348.110 ;
        RECT -33.410 348.035 -32.980 348.620 ;
        RECT -43.140 347.785 -42.710 347.940 ;
        RECT -60.405 346.920 -59.195 347.090 ;
        RECT -60.405 346.220 -59.975 346.920 ;
        RECT -62.835 345.495 -62.440 345.530 ;
        RECT -62.835 344.045 -62.530 345.495 ;
        RECT -51.510 345.155 -51.080 347.565 ;
        RECT -47.520 347.480 -42.710 347.785 ;
        RECT -45.480 345.570 -45.175 347.480 ;
        RECT -43.140 347.130 -42.710 347.480 ;
        RECT -34.245 347.605 -32.980 348.035 ;
        RECT -43.140 346.960 -41.930 347.130 ;
        RECT -43.140 346.260 -42.710 346.960 ;
        RECT -52.790 344.985 -51.080 345.155 ;
        RECT -51.510 344.175 -51.080 344.985 ;
        RECT -62.835 343.875 -60.730 344.045 ;
        RECT -52.790 344.005 -51.080 344.175 ;
        RECT -62.835 343.870 -62.270 343.875 ;
        RECT -62.835 343.285 -62.530 343.870 ;
        RECT -51.510 343.305 -51.080 344.005 ;
        RECT -45.570 345.535 -45.175 345.570 ;
        RECT -45.570 344.085 -45.265 345.535 ;
        RECT -34.245 345.195 -33.815 347.605 ;
        RECT -35.525 345.025 -33.815 345.195 ;
        RECT -34.245 344.215 -33.815 345.025 ;
        RECT -45.570 343.915 -43.465 344.085 ;
        RECT -35.525 344.045 -33.815 344.215 ;
        RECT -45.570 343.910 -45.005 343.915 ;
        RECT -45.570 343.325 -45.265 343.910 ;
        RECT -34.245 343.345 -33.815 344.045 ;
        RECT -64.885 329.640 -64.320 330.965 ;
        RECT -64.885 329.610 -63.675 329.640 ;
        RECT -64.885 329.440 -62.260 329.610 ;
        RECT -64.885 329.405 -63.675 329.440 ;
        RECT -64.885 328.430 -64.320 329.405 ;
        RECT -53.255 329.205 -52.825 331.280 ;
        RECT -54.035 329.035 -52.825 329.205 ;
        RECT -53.255 328.880 -52.825 329.035 ;
        RECT -53.255 328.575 -50.485 328.880 ;
        RECT -64.885 328.400 -63.725 328.430 ;
        RECT -64.885 328.230 -62.260 328.400 ;
        RECT -64.885 328.195 -63.725 328.230 ;
        RECT -53.255 328.225 -52.825 328.575 ;
        RECT -64.885 327.450 -64.320 328.195 ;
        RECT -54.035 328.055 -52.825 328.225 ;
        RECT -64.885 327.420 -63.730 327.450 ;
        RECT -64.885 327.250 -62.260 327.420 ;
        RECT -53.255 327.355 -52.825 328.055 ;
        RECT -64.885 327.215 -63.730 327.250 ;
        RECT -64.885 323.885 -64.320 327.215 ;
        RECT -50.790 327.030 -50.485 328.575 ;
        RECT -50.790 326.630 -50.345 327.030 ;
        RECT -60.505 324.210 -60.075 325.435 ;
        RECT -50.775 325.180 -50.345 326.630 ;
        RECT -52.500 325.010 -50.345 325.180 ;
        RECT -50.960 325.005 -50.345 325.010 ;
        RECT -60.505 324.040 -59.295 324.210 ;
        RECT -50.775 324.135 -50.345 325.005 ;
        RECT -60.505 323.885 -60.075 324.040 ;
        RECT -64.885 323.580 -60.075 323.885 ;
        RECT -62.845 321.670 -62.540 323.580 ;
        RECT -60.505 323.230 -60.075 323.580 ;
        RECT -51.610 323.705 -50.345 324.135 ;
        RECT -47.385 324.830 -46.580 325.395 ;
        RECT -47.385 324.825 -45.995 324.830 ;
        RECT -47.385 324.655 -44.550 324.825 ;
        RECT -47.385 324.645 -45.995 324.655 ;
        RECT -60.505 323.060 -59.295 323.230 ;
        RECT -60.505 322.360 -60.075 323.060 ;
        RECT -62.935 321.635 -62.540 321.670 ;
        RECT -62.935 320.185 -62.630 321.635 ;
        RECT -51.610 321.295 -51.180 323.705 ;
        RECT -52.890 321.125 -51.180 321.295 ;
        RECT -51.610 320.315 -51.180 321.125 ;
        RECT -62.935 320.015 -60.830 320.185 ;
        RECT -52.890 320.145 -51.180 320.315 ;
        RECT -62.935 320.010 -62.370 320.015 ;
        RECT -62.935 319.425 -62.630 320.010 ;
        RECT -51.610 319.445 -51.180 320.145 ;
        RECT -47.385 323.195 -46.580 324.645 ;
        RECT -47.385 323.025 -43.550 323.195 ;
        RECT -47.385 323.010 -46.000 323.025 ;
        RECT -47.385 322.555 -46.580 323.010 ;
        RECT -47.385 322.545 -46.005 322.555 ;
        RECT -47.385 322.375 -43.550 322.545 ;
        RECT -47.385 322.370 -46.005 322.375 ;
        RECT -47.385 318.780 -46.580 322.370 ;
        RECT -47.385 318.595 -46.560 318.780 ;
        RECT -47.385 318.590 -46.005 318.595 ;
        RECT -47.385 318.420 -44.550 318.590 ;
        RECT -47.385 318.410 -46.005 318.420 ;
        RECT -47.385 318.030 -46.560 318.410 ;
        RECT -47.125 316.290 -46.560 318.030 ;
        RECT -47.465 315.725 -46.560 316.290 ;
        RECT -64.730 311.300 -64.165 312.625 ;
        RECT -64.730 311.270 -63.520 311.300 ;
        RECT -64.730 311.100 -62.105 311.270 ;
        RECT -64.730 311.065 -63.520 311.100 ;
        RECT -64.730 310.090 -64.165 311.065 ;
        RECT -53.100 310.865 -52.670 312.940 ;
        RECT -53.880 310.695 -52.670 310.865 ;
        RECT -53.100 310.540 -52.670 310.695 ;
        RECT -47.465 311.340 -46.900 315.725 ;
        RECT -47.465 311.310 -46.255 311.340 ;
        RECT -47.465 311.140 -44.840 311.310 ;
        RECT -47.465 311.105 -46.255 311.140 ;
        RECT -53.100 310.235 -50.330 310.540 ;
        RECT -64.730 310.060 -63.570 310.090 ;
        RECT -64.730 309.890 -62.105 310.060 ;
        RECT -64.730 309.855 -63.570 309.890 ;
        RECT -53.100 309.885 -52.670 310.235 ;
        RECT -64.730 309.110 -64.165 309.855 ;
        RECT -53.880 309.715 -52.670 309.885 ;
        RECT -64.730 309.080 -63.575 309.110 ;
        RECT -64.730 308.910 -62.105 309.080 ;
        RECT -53.100 309.015 -52.670 309.715 ;
        RECT -64.730 308.875 -63.575 308.910 ;
        RECT -64.730 305.545 -64.165 308.875 ;
        RECT -50.635 308.690 -50.330 310.235 ;
        RECT -47.465 310.130 -46.900 311.105 ;
        RECT -35.835 310.905 -35.405 312.980 ;
        RECT -36.615 310.735 -35.405 310.905 ;
        RECT -35.835 310.580 -35.405 310.735 ;
        RECT -35.835 310.275 -33.065 310.580 ;
        RECT -47.465 310.100 -46.305 310.130 ;
        RECT -47.465 309.930 -44.840 310.100 ;
        RECT -47.465 309.895 -46.305 309.930 ;
        RECT -35.835 309.925 -35.405 310.275 ;
        RECT -47.465 309.150 -46.900 309.895 ;
        RECT -36.615 309.755 -35.405 309.925 ;
        RECT -47.465 309.120 -46.310 309.150 ;
        RECT -47.465 308.950 -44.840 309.120 ;
        RECT -35.835 309.055 -35.405 309.755 ;
        RECT -47.465 308.915 -46.310 308.950 ;
        RECT -50.635 308.290 -50.190 308.690 ;
        RECT -60.350 305.870 -59.920 307.095 ;
        RECT -50.620 306.840 -50.190 308.290 ;
        RECT -52.345 306.670 -50.190 306.840 ;
        RECT -50.805 306.665 -50.190 306.670 ;
        RECT -60.350 305.700 -59.140 305.870 ;
        RECT -50.620 305.795 -50.190 306.665 ;
        RECT -60.350 305.545 -59.920 305.700 ;
        RECT -64.730 305.240 -59.920 305.545 ;
        RECT -62.690 303.330 -62.385 305.240 ;
        RECT -60.350 304.890 -59.920 305.240 ;
        RECT -51.455 305.365 -50.190 305.795 ;
        RECT -47.465 305.585 -46.900 308.915 ;
        RECT -33.370 308.730 -33.065 310.275 ;
        RECT -33.370 308.330 -32.925 308.730 ;
        RECT -33.355 308.040 -32.925 308.330 ;
        RECT -30.620 308.040 -28.090 348.620 ;
        RECT -43.085 305.910 -42.655 307.135 ;
        RECT -33.355 306.880 -28.090 308.040 ;
        RECT -35.080 306.710 -28.090 306.880 ;
        RECT -33.540 306.705 -28.090 306.710 ;
        RECT -33.355 306.625 -28.090 306.705 ;
        RECT -43.085 305.740 -41.875 305.910 ;
        RECT -33.355 305.835 -32.925 306.625 ;
        RECT -43.085 305.585 -42.655 305.740 ;
        RECT -60.350 304.720 -59.140 304.890 ;
        RECT -60.350 304.020 -59.920 304.720 ;
        RECT -62.780 303.295 -62.385 303.330 ;
        RECT -62.780 301.845 -62.475 303.295 ;
        RECT -51.455 302.955 -51.025 305.365 ;
        RECT -47.465 305.280 -42.655 305.585 ;
        RECT -45.425 303.370 -45.120 305.280 ;
        RECT -43.085 304.930 -42.655 305.280 ;
        RECT -34.190 305.405 -32.925 305.835 ;
        RECT -43.085 304.760 -41.875 304.930 ;
        RECT -43.085 304.060 -42.655 304.760 ;
        RECT -52.735 302.785 -51.025 302.955 ;
        RECT -51.455 301.975 -51.025 302.785 ;
        RECT -62.780 301.675 -60.675 301.845 ;
        RECT -52.735 301.805 -51.025 301.975 ;
        RECT -62.780 301.670 -62.215 301.675 ;
        RECT -62.780 301.085 -62.475 301.670 ;
        RECT -51.455 301.105 -51.025 301.805 ;
        RECT -45.515 303.335 -45.120 303.370 ;
        RECT -45.515 301.885 -45.210 303.335 ;
        RECT -34.190 302.995 -33.760 305.405 ;
        RECT -35.470 302.825 -33.760 302.995 ;
        RECT -34.190 302.015 -33.760 302.825 ;
        RECT -45.515 301.715 -43.410 301.885 ;
        RECT -35.470 301.845 -33.760 302.015 ;
        RECT -45.515 301.710 -44.950 301.715 ;
        RECT -45.515 301.125 -45.210 301.710 ;
        RECT -34.190 301.145 -33.760 301.845 ;
        RECT -47.855 288.610 -47.370 289.590 ;
        RECT -42.780 288.820 -42.440 289.315 ;
        RECT -43.575 288.650 -42.440 288.820 ;
        RECT -51.960 288.440 -47.370 288.610 ;
        RECT -47.855 286.610 -47.370 288.440 ;
        RECT -42.780 287.840 -42.440 288.650 ;
        RECT -40.880 289.310 -40.540 289.355 ;
        RECT -40.880 289.140 -39.745 289.310 ;
        RECT -40.880 288.330 -40.540 289.140 ;
        RECT -41.315 288.170 -41.120 288.255 ;
        RECT -43.575 287.670 -42.440 287.840 ;
        RECT -42.780 286.860 -42.440 287.670 ;
        RECT -41.380 288.115 -41.080 288.170 ;
        RECT -40.880 288.160 -39.745 288.330 ;
        RECT -40.880 288.115 -40.540 288.160 ;
        RECT -41.380 287.560 -40.540 288.115 ;
        RECT -41.380 287.485 -41.080 287.560 ;
        RECT -43.575 286.690 -42.440 286.860 ;
        RECT -42.780 286.645 -42.440 286.690 ;
        RECT -51.960 286.440 -47.370 286.610 ;
        RECT -47.855 283.610 -47.370 286.440 ;
        RECT -51.960 283.440 -47.370 283.610 ;
        RECT -47.855 281.610 -47.370 283.440 ;
        RECT -51.960 281.440 -47.370 281.610 ;
        RECT -47.855 278.610 -47.370 281.440 ;
        RECT -41.315 284.060 -41.120 287.485 ;
        RECT -40.880 287.350 -40.540 287.560 ;
        RECT -40.880 287.180 -39.745 287.350 ;
        RECT -40.880 285.125 -40.540 287.180 ;
        RECT -40.880 284.955 -39.745 285.125 ;
        RECT -40.880 284.145 -40.540 284.955 ;
        RECT -40.880 284.060 -39.745 284.145 ;
        RECT -41.315 283.975 -39.745 284.060 ;
        RECT -41.315 283.505 -40.540 283.975 ;
        RECT -42.780 280.105 -42.440 280.600 ;
        RECT -43.575 279.935 -42.440 280.105 ;
        RECT -42.780 279.125 -42.440 279.935 ;
        RECT -43.575 278.955 -42.440 279.125 ;
        RECT -51.960 278.440 -47.370 278.610 ;
        RECT -47.855 276.610 -47.370 278.440 ;
        RECT -42.780 278.145 -42.440 278.955 ;
        RECT -43.575 277.975 -42.440 278.145 ;
        RECT -51.960 276.440 -47.370 276.610 ;
        RECT -47.855 275.320 -47.370 276.440 ;
        RECT -42.780 275.320 -42.440 277.975 ;
        RECT -54.045 274.970 -47.370 275.320 ;
        RECT -43.575 275.150 -42.440 275.320 ;
        RECT -41.315 275.185 -41.120 283.505 ;
        RECT -40.880 283.165 -40.540 283.505 ;
        RECT -40.880 282.995 -39.745 283.165 ;
        RECT -40.880 282.500 -40.540 282.995 ;
        RECT -40.880 275.810 -40.540 275.855 ;
        RECT -40.880 275.640 -39.745 275.810 ;
        RECT -54.045 274.520 -53.040 274.970 ;
        RECT -54.045 274.170 -53.025 274.520 ;
        RECT -42.780 274.340 -42.440 275.150 ;
        RECT -41.410 275.070 -41.110 275.185 ;
        RECT -40.880 275.070 -40.540 275.640 ;
        RECT -41.410 274.830 -40.540 275.070 ;
        RECT -41.410 274.660 -39.745 274.830 ;
        RECT -41.410 274.515 -40.540 274.660 ;
        RECT -41.410 274.500 -41.110 274.515 ;
        RECT -43.575 274.170 -42.440 274.340 ;
        RECT -54.840 274.000 -53.025 274.170 ;
        RECT -54.045 273.190 -53.025 274.000 ;
        RECT -42.780 273.360 -42.440 274.170 ;
        RECT -43.575 273.190 -42.440 273.360 ;
        RECT -54.840 273.020 -53.025 273.190 ;
        RECT -42.780 273.145 -42.440 273.190 ;
        RECT -54.045 272.460 -53.025 273.020 ;
        RECT -54.045 272.290 -51.465 272.460 ;
        RECT -54.045 272.210 -53.025 272.290 ;
        RECT -54.840 272.125 -53.025 272.210 ;
        RECT -54.840 272.040 -53.040 272.125 ;
        RECT -54.045 271.995 -53.040 272.040 ;
        RECT -53.830 270.480 -53.040 271.995 ;
        RECT -41.315 270.680 -41.120 274.500 ;
        RECT -40.880 274.155 -40.540 274.515 ;
        RECT -40.890 273.850 -40.540 274.155 ;
        RECT -40.890 273.680 -39.745 273.850 ;
        RECT -40.890 273.185 -40.540 273.680 ;
        RECT -40.890 271.670 -40.550 273.185 ;
        RECT -40.890 271.625 -40.540 271.670 ;
        RECT -40.890 271.555 -39.745 271.625 ;
        RECT -40.880 271.455 -39.745 271.555 ;
        RECT -40.880 270.680 -40.540 271.455 ;
        RECT -41.315 270.645 -40.540 270.680 ;
        RECT -51.335 270.480 -50.930 270.485 ;
        RECT -53.830 270.075 -50.930 270.480 ;
        RECT -51.510 268.905 -50.930 270.075 ;
        RECT -51.255 268.565 -50.930 268.905 ;
        RECT -53.235 268.395 -50.930 268.565 ;
        RECT -51.255 263.405 -50.930 268.395 ;
        RECT -41.315 270.475 -39.745 270.645 ;
        RECT -41.315 270.125 -40.540 270.475 ;
        RECT -42.780 266.605 -42.440 267.100 ;
        RECT -43.575 266.435 -42.440 266.605 ;
        RECT -42.780 265.625 -42.440 266.435 ;
        RECT -43.575 265.455 -42.440 265.625 ;
        RECT -42.780 264.645 -42.440 265.455 ;
        RECT -43.575 264.475 -42.440 264.645 ;
        RECT -53.740 263.235 -50.930 263.405 ;
        RECT -51.590 262.505 -50.930 263.235 ;
        RECT -51.590 259.825 -51.145 262.505 ;
        RECT -42.780 262.195 -42.440 264.475 ;
        RECT -43.575 262.025 -42.440 262.195 ;
        RECT -42.780 261.215 -42.440 262.025 ;
        RECT -41.315 262.255 -41.120 270.125 ;
        RECT -40.880 269.665 -40.540 270.125 ;
        RECT -40.880 269.495 -39.745 269.665 ;
        RECT -40.880 269.000 -40.540 269.495 ;
        RECT -41.315 261.995 -37.940 262.255 ;
        RECT -41.410 261.335 -37.940 261.995 ;
        RECT -41.315 261.330 -41.120 261.335 ;
        RECT -43.575 261.045 -42.440 261.215 ;
        RECT -42.780 260.235 -42.440 261.045 ;
        RECT -43.575 260.065 -42.440 260.235 ;
        RECT -42.780 260.020 -42.440 260.065 ;
        RECT -38.470 260.620 -37.940 261.335 ;
        RECT -30.620 260.620 -28.090 306.625 ;
        RECT -52.345 259.805 -51.145 259.825 ;
        RECT -53.145 259.635 -51.145 259.805 ;
        RECT -52.345 259.605 -51.145 259.635 ;
        RECT -51.590 259.275 -51.145 259.605 ;
        RECT -38.470 259.275 -18.735 260.620 ;
        RECT -51.590 258.855 -18.735 259.275 ;
        RECT -52.350 258.825 -18.735 258.855 ;
        RECT -53.145 258.655 -18.735 258.825 ;
        RECT -52.350 258.635 -18.735 258.655 ;
        RECT -51.590 258.530 -18.735 258.635 ;
        RECT -51.590 255.095 -51.145 258.530 ;
        RECT -38.470 257.895 -18.735 258.530 ;
        RECT -38.470 255.135 -37.940 257.895 ;
        RECT -39.215 255.100 -37.940 255.135 ;
        RECT -52.345 255.075 -51.145 255.095 ;
        RECT -53.145 254.905 -51.145 255.075 ;
        RECT -40.055 254.930 -37.940 255.100 ;
        RECT -30.620 254.980 -28.090 257.895 ;
        RECT -52.345 254.875 -51.145 254.905 ;
        RECT -39.215 254.895 -37.940 254.930 ;
        RECT -51.590 254.125 -51.145 254.875 ;
        RECT -38.470 254.165 -37.940 254.895 ;
        RECT -52.350 254.095 -51.145 254.125 ;
        RECT -39.200 254.120 -37.940 254.165 ;
        RECT -53.145 253.925 -51.145 254.095 ;
        RECT -40.055 253.950 -37.940 254.120 ;
        RECT -39.200 253.925 -37.940 253.950 ;
        RECT -52.350 253.905 -51.145 253.925 ;
        RECT -51.590 253.260 -51.145 253.905 ;
        RECT -38.470 253.405 -37.940 253.925 ;
        RECT -65.560 248.670 -65.220 248.715 ;
        RECT -66.355 248.500 -65.220 248.670 ;
        RECT -65.560 247.690 -65.220 248.500 ;
        RECT -66.355 247.520 -65.220 247.690 ;
        RECT -63.660 248.180 -63.320 248.675 ;
        RECT -63.660 248.010 -62.525 248.180 ;
        RECT -64.980 247.530 -64.785 247.615 ;
        RECT -65.560 247.475 -65.220 247.520 ;
        RECT -65.020 247.475 -64.720 247.530 ;
        RECT -65.560 246.920 -64.720 247.475 ;
        RECT -65.560 246.710 -65.220 246.920 ;
        RECT -65.020 246.845 -64.720 246.920 ;
        RECT -63.660 247.200 -63.320 248.010 ;
        RECT -63.660 247.030 -62.525 247.200 ;
        RECT -66.355 246.540 -65.220 246.710 ;
        RECT -65.560 244.485 -65.220 246.540 ;
        RECT -66.355 244.315 -65.220 244.485 ;
        RECT -65.560 243.505 -65.220 244.315 ;
        RECT -66.355 243.420 -65.220 243.505 ;
        RECT -64.980 243.420 -64.785 246.845 ;
        RECT -63.660 246.220 -63.320 247.030 ;
        RECT -63.660 246.050 -62.525 246.220 ;
        RECT -63.660 246.005 -63.320 246.050 ;
        RECT -66.355 243.335 -64.785 243.420 ;
        RECT -65.560 242.865 -64.785 243.335 ;
        RECT -65.560 242.525 -65.220 242.865 ;
        RECT -66.355 242.355 -65.220 242.525 ;
        RECT -65.560 241.860 -65.220 242.355 ;
        RECT -65.560 235.170 -65.220 235.215 ;
        RECT -66.355 235.000 -65.220 235.170 ;
        RECT -65.560 234.430 -65.220 235.000 ;
        RECT -64.980 234.545 -64.785 242.865 ;
        RECT -63.660 239.465 -63.320 239.960 ;
        RECT -63.660 239.295 -62.525 239.465 ;
        RECT -63.660 238.485 -63.320 239.295 ;
        RECT -63.660 238.315 -62.525 238.485 ;
        RECT -63.660 237.505 -63.320 238.315 ;
        RECT -63.660 237.335 -62.525 237.505 ;
        RECT -63.660 234.680 -63.320 237.335 ;
        RECT -64.990 234.430 -64.690 234.545 ;
        RECT -65.560 234.190 -64.690 234.430 ;
        RECT -66.355 234.020 -64.690 234.190 ;
        RECT -65.560 233.875 -64.690 234.020 ;
        RECT -65.560 233.515 -65.220 233.875 ;
        RECT -64.990 233.860 -64.690 233.875 ;
        RECT -63.660 234.510 -62.525 234.680 ;
        RECT -65.560 233.210 -65.210 233.515 ;
        RECT -66.355 233.040 -65.210 233.210 ;
        RECT -65.560 232.545 -65.210 233.040 ;
        RECT -65.550 231.030 -65.210 232.545 ;
        RECT -65.560 230.985 -65.210 231.030 ;
        RECT -66.355 230.915 -65.210 230.985 ;
        RECT -66.355 230.815 -65.220 230.915 ;
        RECT -65.560 230.040 -65.220 230.815 ;
        RECT -64.980 230.040 -64.785 233.860 ;
        RECT -63.660 233.700 -63.320 234.510 ;
        RECT -63.660 233.530 -62.525 233.700 ;
        RECT -63.660 232.720 -63.320 233.530 ;
        RECT -63.660 232.550 -62.525 232.720 ;
        RECT -63.660 232.505 -63.320 232.550 ;
        RECT -65.560 230.005 -64.785 230.040 ;
        RECT -66.355 229.835 -64.785 230.005 ;
        RECT -65.560 229.485 -64.785 229.835 ;
        RECT -65.560 229.025 -65.220 229.485 ;
        RECT -66.355 228.855 -65.220 229.025 ;
        RECT -65.560 228.360 -65.220 228.855 ;
        RECT -64.980 222.520 -64.785 229.485 ;
        RECT -69.575 221.355 -64.785 222.520 ;
        RECT -63.660 225.965 -63.320 226.460 ;
        RECT -63.660 225.795 -62.525 225.965 ;
        RECT -63.660 224.985 -63.320 225.795 ;
        RECT -63.660 224.815 -62.525 224.985 ;
        RECT -63.660 224.005 -63.320 224.815 ;
        RECT -63.660 223.835 -62.525 224.005 ;
        RECT -63.660 221.555 -63.320 223.835 ;
        RECT -63.660 221.385 -62.525 221.555 ;
        RECT -69.575 221.215 -64.690 221.355 ;
        RECT -69.575 213.600 -68.270 221.215 ;
        RECT -64.990 220.695 -64.690 221.215 ;
        RECT -64.980 220.690 -64.785 220.695 ;
        RECT -63.660 220.575 -63.320 221.385 ;
        RECT -63.660 220.405 -62.525 220.575 ;
        RECT -20.400 220.510 -18.735 257.895 ;
        RECT -63.660 219.595 -63.320 220.405 ;
        RECT -63.660 219.425 -62.525 219.595 ;
        RECT -63.660 219.380 -63.320 219.425 ;
        RECT -69.575 212.295 -58.065 213.600 ;
        RECT -24.100 212.350 -18.735 220.510 ;
        RECT -61.585 209.970 -61.345 210.230 ;
        RECT -70.345 209.700 -61.345 209.970 ;
        RECT -70.345 209.480 -70.075 209.700 ;
        RECT -61.585 209.490 -61.345 209.700 ;
        RECT -59.370 210.055 -58.065 212.295 ;
        RECT -70.550 209.210 -69.925 209.480 ;
        RECT -62.260 209.255 -62.040 209.325 ;
        RECT -64.685 208.985 -62.040 209.255 ;
        RECT -64.685 208.760 -64.415 208.985 ;
        RECT -77.455 208.010 -76.765 208.690 ;
        RECT -70.550 208.490 -64.415 208.760 ;
        RECT -62.260 208.710 -62.040 208.985 ;
        RECT -59.370 208.750 -52.790 210.055 ;
        RECT -62.895 208.185 -62.695 208.700 ;
        RECT -77.455 51.860 -76.775 208.010 ;
        RECT -70.550 207.915 -62.695 208.185 ;
        RECT -54.095 205.585 -52.790 208.750 ;
        RECT -20.400 205.585 -18.735 212.350 ;
        RECT -64.705 204.280 -18.735 205.585 ;
        RECT -64.705 203.465 -64.070 204.280 ;
        RECT -53.360 203.515 -52.880 203.535 ;
        RECT -53.790 203.495 -52.880 203.515 ;
        RECT -65.045 203.445 -64.070 203.465 ;
        RECT -66.040 203.275 -64.070 203.445 ;
        RECT -54.785 203.325 -52.880 203.495 ;
        RECT -53.790 203.300 -52.880 203.325 ;
        RECT -65.045 203.250 -64.070 203.275 ;
        RECT -64.705 201.920 -64.070 203.250 ;
        RECT -53.360 203.290 -52.880 203.300 ;
        RECT -50.655 203.290 -49.350 204.280 ;
        RECT -53.360 202.305 -49.350 203.290 ;
        RECT -53.360 201.970 -52.880 202.305 ;
        RECT -53.780 201.950 -52.880 201.970 ;
        RECT -65.035 201.900 -64.070 201.920 ;
        RECT -66.040 201.730 -64.070 201.900 ;
        RECT -54.785 201.780 -52.880 201.950 ;
        RECT -53.780 201.755 -52.880 201.780 ;
        RECT -65.035 201.705 -64.070 201.730 ;
        RECT -64.705 200.245 -64.070 201.705 ;
        RECT -53.360 200.775 -52.880 201.755 ;
        RECT -50.655 200.775 -49.350 202.305 ;
        RECT -53.360 200.375 -49.350 200.775 ;
        RECT -66.300 196.410 -65.000 196.580 ;
        RECT -66.300 196.395 -66.010 196.410 ;
        RECT -66.300 195.985 -66.115 196.395 ;
        RECT -66.605 195.800 -66.115 195.985 ;
        RECT -66.605 194.515 -66.420 195.800 ;
        RECT -64.445 194.515 -64.180 200.245 ;
        RECT -53.190 199.790 -49.350 200.375 ;
        RECT -53.190 198.210 -52.925 199.790 ;
        RECT -50.655 198.210 -49.350 199.790 ;
        RECT -53.190 198.115 -49.350 198.210 ;
        RECT -45.060 203.290 -43.755 204.280 ;
        RECT -41.530 203.515 -41.050 203.535 ;
        RECT -41.530 203.495 -40.620 203.515 ;
        RECT -41.530 203.325 -39.625 203.495 ;
        RECT -30.340 203.465 -29.705 204.280 ;
        RECT -30.340 203.445 -29.365 203.465 ;
        RECT -41.530 203.300 -40.620 203.325 ;
        RECT -41.530 203.290 -41.050 203.300 ;
        RECT -45.060 202.305 -41.050 203.290 ;
        RECT -45.060 200.775 -43.755 202.305 ;
        RECT -41.530 201.970 -41.050 202.305 ;
        RECT -30.340 203.275 -28.370 203.445 ;
        RECT -30.340 203.250 -29.365 203.275 ;
        RECT -41.530 201.950 -40.630 201.970 ;
        RECT -41.530 201.780 -39.625 201.950 ;
        RECT -30.340 201.920 -29.705 203.250 ;
        RECT -30.340 201.900 -29.375 201.920 ;
        RECT -41.530 201.755 -40.630 201.780 ;
        RECT -41.530 200.775 -41.050 201.755 ;
        RECT -45.060 200.375 -41.050 200.775 ;
        RECT -30.340 201.730 -28.370 201.900 ;
        RECT -30.340 201.705 -29.375 201.730 ;
        RECT -45.060 199.790 -41.220 200.375 ;
        RECT -30.340 200.245 -29.705 201.705 ;
        RECT -45.060 198.210 -43.755 199.790 ;
        RECT -41.485 198.210 -41.220 199.790 ;
        RECT -45.060 198.115 -41.220 198.210 ;
        RECT -53.190 197.225 -41.220 198.115 ;
        RECT -55.045 196.460 -53.745 196.630 ;
        RECT -55.045 196.445 -54.755 196.460 ;
        RECT -55.045 196.035 -54.860 196.445 ;
        RECT -66.605 194.510 -66.005 194.515 ;
        RECT -65.060 194.510 -64.180 194.515 ;
        RECT -66.605 194.340 -64.180 194.510 ;
        RECT -55.350 195.850 -54.860 196.035 ;
        RECT -55.350 194.565 -55.165 195.850 ;
        RECT -53.190 195.545 -52.925 197.225 ;
        RECT -50.655 196.810 -43.755 197.225 ;
        RECT -50.655 195.545 -49.350 196.810 ;
        RECT -53.190 194.565 -49.350 195.545 ;
        RECT -55.350 194.560 -54.750 194.565 ;
        RECT -53.805 194.560 -49.350 194.565 ;
        RECT -55.350 194.390 -52.925 194.560 ;
        RECT -55.350 194.380 -54.750 194.390 ;
        RECT -53.805 194.370 -52.925 194.390 ;
        RECT -66.605 194.330 -66.005 194.340 ;
        RECT -65.060 194.320 -64.180 194.340 ;
        RECT -64.445 188.485 -64.180 194.320 ;
        RECT -52.350 192.470 -52.025 192.635 ;
        RECT -50.655 192.470 -49.350 194.560 ;
        RECT -52.350 192.145 -49.350 192.470 ;
        RECT -54.835 191.975 -49.350 192.145 ;
        RECT -52.350 191.740 -49.350 191.975 ;
        RECT -52.350 190.670 -52.025 191.740 ;
        RECT -50.655 190.670 -49.350 191.740 ;
        RECT -52.350 189.940 -49.350 190.670 ;
        RECT -52.350 189.340 -52.025 189.940 ;
        RECT -50.655 189.340 -49.350 189.940 ;
        RECT -52.350 188.610 -49.350 189.340 ;
        RECT -64.615 188.465 -64.135 188.485 ;
        RECT -65.045 188.445 -64.135 188.465 ;
        RECT -66.040 188.275 -64.135 188.445 ;
        RECT -65.045 188.250 -64.135 188.275 ;
        RECT -64.615 186.920 -64.135 188.250 ;
        RECT -52.350 187.115 -52.025 188.610 ;
        RECT -50.655 188.385 -49.350 188.610 ;
        RECT -45.060 195.545 -43.755 196.810 ;
        RECT -41.485 195.545 -41.220 197.225 ;
        RECT -40.665 196.460 -39.365 196.630 ;
        RECT -39.655 196.445 -39.365 196.460 ;
        RECT -39.550 196.035 -39.365 196.445 ;
        RECT -39.550 195.850 -39.060 196.035 ;
        RECT -45.060 194.565 -41.220 195.545 ;
        RECT -39.245 194.565 -39.060 195.850 ;
        RECT -45.060 194.560 -40.605 194.565 ;
        RECT -39.660 194.560 -39.060 194.565 ;
        RECT -45.060 192.470 -43.755 194.560 ;
        RECT -41.485 194.390 -39.060 194.560 ;
        RECT -41.485 194.370 -40.605 194.390 ;
        RECT -39.660 194.380 -39.060 194.390 ;
        RECT -30.230 194.515 -29.965 200.245 ;
        RECT -29.410 196.410 -28.110 196.580 ;
        RECT -28.400 196.395 -28.110 196.410 ;
        RECT -28.295 195.985 -28.110 196.395 ;
        RECT -28.295 195.800 -27.805 195.985 ;
        RECT -27.990 194.515 -27.805 195.800 ;
        RECT -30.230 194.510 -29.350 194.515 ;
        RECT -28.405 194.510 -27.805 194.515 ;
        RECT -30.230 194.340 -27.805 194.510 ;
        RECT -30.230 194.320 -29.350 194.340 ;
        RECT -28.405 194.330 -27.805 194.340 ;
        RECT -42.385 192.470 -42.060 192.635 ;
        RECT -45.060 192.145 -42.060 192.470 ;
        RECT -45.060 191.975 -39.575 192.145 ;
        RECT -45.060 191.740 -42.060 191.975 ;
        RECT -45.060 190.670 -43.755 191.740 ;
        RECT -42.385 190.670 -42.060 191.740 ;
        RECT -45.060 189.940 -42.060 190.670 ;
        RECT -45.060 189.340 -43.755 189.940 ;
        RECT -42.385 189.340 -42.060 189.940 ;
        RECT -45.060 188.610 -42.060 189.340 ;
        RECT -45.060 188.385 -43.755 188.610 ;
        RECT -50.655 187.115 -43.755 188.385 ;
        RECT -42.385 187.115 -42.060 188.610 ;
        RECT -30.230 188.485 -29.965 194.320 ;
        RECT -52.350 187.080 -42.060 187.115 ;
        RECT -52.350 186.985 -49.350 187.080 ;
        RECT -65.035 186.900 -64.135 186.920 ;
        RECT -66.040 186.730 -64.135 186.900 ;
        RECT -54.330 186.815 -49.350 186.985 ;
        RECT -65.035 186.705 -64.135 186.730 ;
        RECT -64.615 185.325 -64.135 186.705 ;
        RECT -52.350 186.385 -49.350 186.815 ;
        RECT -52.350 186.265 -52.025 186.385 ;
        RECT -66.300 181.410 -65.000 181.580 ;
        RECT -66.300 181.395 -66.010 181.410 ;
        RECT -66.300 180.985 -66.115 181.395 ;
        RECT -66.605 180.800 -66.115 180.985 ;
        RECT -66.605 179.515 -66.420 180.800 ;
        RECT -64.445 179.515 -64.180 185.325 ;
        RECT -53.260 183.940 -52.955 183.970 ;
        RECT -50.655 183.940 -49.350 186.385 ;
        RECT -53.260 183.385 -49.350 183.940 ;
        RECT -53.520 183.380 -49.350 183.385 ;
        RECT -55.060 183.210 -49.350 183.380 ;
        RECT -53.260 183.185 -49.350 183.210 ;
        RECT -53.260 182.475 -52.955 183.185 ;
        RECT -50.655 182.475 -49.350 183.185 ;
        RECT -53.260 182.315 -49.350 182.475 ;
        RECT -45.060 186.985 -42.060 187.080 ;
        RECT -30.275 188.465 -29.795 188.485 ;
        RECT -30.275 188.445 -29.365 188.465 ;
        RECT -30.275 188.275 -28.370 188.445 ;
        RECT -30.275 188.250 -29.365 188.275 ;
        RECT -45.060 186.815 -40.080 186.985 ;
        RECT -30.275 186.920 -29.795 188.250 ;
        RECT -30.275 186.900 -29.375 186.920 ;
        RECT -45.060 186.385 -42.060 186.815 ;
        RECT -45.060 183.940 -43.755 186.385 ;
        RECT -42.385 186.265 -42.060 186.385 ;
        RECT -30.275 186.730 -28.370 186.900 ;
        RECT -30.275 186.705 -29.375 186.730 ;
        RECT -30.275 185.325 -29.795 186.705 ;
        RECT -41.455 183.940 -41.150 183.970 ;
        RECT -45.060 183.385 -41.150 183.940 ;
        RECT -45.060 183.380 -40.890 183.385 ;
        RECT -45.060 183.210 -39.350 183.380 ;
        RECT -45.060 183.185 -41.150 183.210 ;
        RECT -45.060 182.475 -43.755 183.185 ;
        RECT -41.455 182.475 -41.150 183.185 ;
        RECT -45.060 182.315 -41.150 182.475 ;
        RECT -53.260 181.760 -41.150 182.315 ;
        RECT -53.350 181.720 -41.060 181.760 ;
        RECT -55.815 180.335 -55.385 181.035 ;
        RECT -56.595 180.165 -55.385 180.335 ;
        RECT -66.605 179.510 -66.005 179.515 ;
        RECT -65.060 179.510 -64.180 179.515 ;
        RECT -66.605 179.340 -64.180 179.510 ;
        RECT -55.815 179.815 -55.385 180.165 ;
        RECT -53.350 180.265 -53.045 181.720 ;
        RECT -50.655 181.010 -43.755 181.720 ;
        RECT -50.655 180.265 -49.350 181.010 ;
        RECT -53.350 179.815 -49.350 180.265 ;
        RECT -55.815 179.510 -49.350 179.815 ;
        RECT -55.815 179.355 -55.385 179.510 ;
        RECT -66.605 179.330 -66.005 179.340 ;
        RECT -65.060 179.320 -64.180 179.340 ;
        RECT -64.445 175.985 -64.180 179.320 ;
        RECT -56.595 179.185 -55.385 179.355 ;
        RECT -55.815 177.960 -55.385 179.185 ;
        RECT -64.615 175.965 -64.135 175.985 ;
        RECT -65.045 175.945 -64.135 175.965 ;
        RECT -66.040 175.775 -64.135 175.945 ;
        RECT -65.045 175.750 -64.135 175.775 ;
        RECT -66.730 174.135 -66.460 174.830 ;
        RECT -64.615 174.420 -64.135 175.750 ;
        RECT -53.270 175.640 -52.965 175.945 ;
        RECT -50.655 175.640 -49.350 179.510 ;
        RECT -53.270 175.360 -49.350 175.640 ;
        RECT -53.530 175.355 -49.350 175.360 ;
        RECT -55.070 175.185 -49.350 175.355 ;
        RECT -65.035 174.400 -64.135 174.420 ;
        RECT -66.040 174.230 -64.135 174.400 ;
        RECT -65.035 174.205 -64.135 174.230 ;
        RECT -64.615 172.825 -64.135 174.205 ;
        RECT -53.270 175.025 -49.350 175.185 ;
        RECT -45.060 180.265 -43.755 181.010 ;
        RECT -41.365 180.265 -41.060 181.720 ;
        RECT -45.060 179.815 -41.060 180.265 ;
        RECT -39.025 180.335 -38.595 181.035 ;
        RECT -39.025 180.165 -37.815 180.335 ;
        RECT -39.025 179.815 -38.595 180.165 ;
        RECT -45.060 179.510 -38.595 179.815 ;
        RECT -45.060 175.640 -43.755 179.510 ;
        RECT -39.025 179.355 -38.595 179.510 ;
        RECT -30.230 179.515 -29.965 185.325 ;
        RECT -29.410 181.410 -28.110 181.580 ;
        RECT -28.400 181.395 -28.110 181.410 ;
        RECT -28.295 180.985 -28.110 181.395 ;
        RECT -28.295 180.800 -27.805 180.985 ;
        RECT -27.990 179.515 -27.805 180.800 ;
        RECT -30.230 179.510 -29.350 179.515 ;
        RECT -28.405 179.510 -27.805 179.515 ;
        RECT -39.025 179.185 -37.815 179.355 ;
        RECT -30.230 179.340 -27.805 179.510 ;
        RECT -30.230 179.320 -29.350 179.340 ;
        RECT -28.405 179.330 -27.805 179.340 ;
        RECT -39.025 177.960 -38.595 179.185 ;
        RECT -30.230 175.985 -29.965 179.320 ;
        RECT -30.275 175.965 -29.795 175.985 ;
        RECT -30.275 175.945 -29.365 175.965 ;
        RECT -41.445 175.640 -41.140 175.945 ;
        RECT -45.060 175.360 -41.140 175.640 ;
        RECT -30.275 175.775 -28.370 175.945 ;
        RECT -30.275 175.750 -29.365 175.775 ;
        RECT -45.060 175.355 -40.880 175.360 ;
        RECT -45.060 175.185 -39.340 175.355 ;
        RECT -45.060 175.025 -41.140 175.185 ;
        RECT -53.270 175.020 -41.140 175.025 ;
        RECT -53.270 173.990 -52.965 175.020 ;
        RECT -50.655 173.990 -43.755 175.020 ;
        RECT -41.445 173.990 -41.140 175.020 ;
        RECT -53.270 173.735 -41.140 173.990 ;
        RECT -30.275 174.420 -29.795 175.750 ;
        RECT -30.275 174.400 -29.375 174.420 ;
        RECT -30.275 174.230 -28.370 174.400 ;
        RECT -30.275 174.205 -29.375 174.230 ;
        RECT -53.360 173.720 -41.050 173.735 ;
        RECT -53.360 173.370 -49.350 173.720 ;
        RECT -66.760 168.745 -66.490 169.440 ;
        RECT -66.300 168.910 -65.000 169.080 ;
        RECT -66.300 168.895 -66.010 168.910 ;
        RECT -66.300 168.485 -66.115 168.895 ;
        RECT -66.605 168.300 -66.115 168.485 ;
        RECT -66.605 167.015 -66.420 168.300 ;
        RECT -64.445 167.015 -64.180 172.825 ;
        RECT -55.825 172.310 -55.395 173.010 ;
        RECT -56.605 172.140 -55.395 172.310 ;
        RECT -55.825 171.790 -55.395 172.140 ;
        RECT -53.360 172.240 -53.055 173.370 ;
        RECT -50.655 172.240 -49.350 173.370 ;
        RECT -53.360 171.790 -49.350 172.240 ;
        RECT -55.825 171.485 -49.350 171.790 ;
        RECT -55.825 171.330 -55.395 171.485 ;
        RECT -56.605 171.160 -55.395 171.330 ;
        RECT -55.825 169.935 -55.395 171.160 ;
        RECT -50.655 169.825 -49.350 171.485 ;
        RECT -45.060 173.370 -41.050 173.720 ;
        RECT -45.060 172.240 -43.755 173.370 ;
        RECT -41.355 172.240 -41.050 173.370 ;
        RECT -45.060 171.790 -41.050 172.240 ;
        RECT -39.015 172.310 -38.585 173.010 ;
        RECT -30.275 172.825 -29.795 174.205 ;
        RECT -27.950 174.135 -27.680 174.830 ;
        RECT -39.015 172.140 -37.805 172.310 ;
        RECT -39.015 171.790 -38.585 172.140 ;
        RECT -45.060 171.485 -38.585 171.790 ;
        RECT -45.060 169.825 -43.755 171.485 ;
        RECT -39.015 171.330 -38.585 171.485 ;
        RECT -39.015 171.160 -37.805 171.330 ;
        RECT -39.015 169.935 -38.585 171.160 ;
        RECT -50.655 168.520 -43.755 169.825 ;
        RECT -52.305 167.515 -51.980 167.825 ;
        RECT -50.655 167.515 -49.350 168.520 ;
        RECT -52.305 167.335 -49.350 167.515 ;
        RECT -54.790 167.165 -49.350 167.335 ;
        RECT -66.605 167.010 -66.005 167.015 ;
        RECT -65.060 167.010 -64.180 167.015 ;
        RECT -66.605 166.840 -64.180 167.010 ;
        RECT -66.605 166.830 -66.005 166.840 ;
        RECT -65.060 166.820 -64.180 166.840 ;
        RECT -64.445 163.485 -64.180 166.820 ;
        RECT -52.305 166.865 -49.350 167.165 ;
        RECT -52.305 165.285 -51.980 166.865 ;
        RECT -50.655 165.640 -49.350 166.865 ;
        RECT -45.060 167.515 -43.755 168.520 ;
        RECT -42.430 167.515 -42.105 167.825 ;
        RECT -45.060 167.335 -42.105 167.515 ;
        RECT -45.060 167.165 -39.620 167.335 ;
        RECT -45.060 166.865 -42.105 167.165 ;
        RECT -45.060 165.640 -43.755 166.865 ;
        RECT -50.655 165.285 -43.755 165.640 ;
        RECT -42.430 165.285 -42.105 166.865 ;
        RECT -52.305 164.635 -42.105 165.285 ;
        RECT -52.305 163.700 -51.980 164.635 ;
        RECT -50.655 164.335 -43.755 164.635 ;
        RECT -50.655 163.700 -49.350 164.335 ;
        RECT -64.615 163.465 -64.135 163.485 ;
        RECT -65.045 163.445 -64.135 163.465 ;
        RECT -66.040 163.275 -64.135 163.445 ;
        RECT -65.045 163.250 -64.135 163.275 ;
        RECT -66.730 161.635 -66.460 162.330 ;
        RECT -64.615 161.920 -64.135 163.250 ;
        RECT -52.305 163.050 -49.350 163.700 ;
        RECT -52.305 162.175 -51.980 163.050 ;
        RECT -54.285 162.170 -51.980 162.175 ;
        RECT -50.655 162.170 -49.350 163.050 ;
        RECT -54.285 162.005 -49.350 162.170 ;
        RECT -65.035 161.900 -64.135 161.920 ;
        RECT -66.040 161.730 -64.135 161.900 ;
        RECT -65.035 161.705 -64.135 161.730 ;
        RECT -64.615 160.325 -64.135 161.705 ;
        RECT -52.305 161.520 -49.350 162.005 ;
        RECT -52.305 161.455 -51.980 161.520 ;
        RECT -66.760 156.245 -66.490 156.940 ;
        RECT -66.300 156.410 -65.000 156.580 ;
        RECT -66.300 156.395 -66.010 156.410 ;
        RECT -66.300 155.985 -66.115 156.395 ;
        RECT -66.605 155.800 -66.115 155.985 ;
        RECT -66.605 154.515 -66.420 155.800 ;
        RECT -64.445 154.515 -64.180 160.325 ;
        RECT -55.215 159.485 -54.875 159.530 ;
        RECT -56.010 159.315 -54.875 159.485 ;
        RECT -55.215 158.505 -54.875 159.315 ;
        RECT -56.010 158.335 -54.875 158.505 ;
        RECT -55.215 157.525 -54.875 158.335 ;
        RECT -53.750 158.215 -53.555 158.220 ;
        RECT -53.845 157.780 -53.545 158.215 ;
        RECT -50.655 157.780 -49.350 161.520 ;
        RECT -45.060 163.700 -43.755 164.335 ;
        RECT -42.430 163.700 -42.105 164.635 ;
        RECT -45.060 163.050 -42.105 163.700 ;
        RECT -30.230 167.015 -29.965 172.825 ;
        RECT -29.410 168.910 -28.110 169.080 ;
        RECT -28.400 168.895 -28.110 168.910 ;
        RECT -28.295 168.485 -28.110 168.895 ;
        RECT -27.920 168.745 -27.650 169.440 ;
        RECT -28.295 168.300 -27.805 168.485 ;
        RECT -27.990 167.015 -27.805 168.300 ;
        RECT -30.230 167.010 -29.350 167.015 ;
        RECT -28.405 167.010 -27.805 167.015 ;
        RECT -30.230 166.840 -27.805 167.010 ;
        RECT -30.230 166.820 -29.350 166.840 ;
        RECT -28.405 166.830 -27.805 166.840 ;
        RECT -30.230 163.485 -29.965 166.820 ;
        RECT -45.060 162.170 -43.755 163.050 ;
        RECT -42.430 162.175 -42.105 163.050 ;
        RECT -30.275 163.465 -29.795 163.485 ;
        RECT -30.275 163.445 -29.365 163.465 ;
        RECT -30.275 163.275 -28.370 163.445 ;
        RECT -30.275 163.250 -29.365 163.275 ;
        RECT -42.430 162.170 -40.125 162.175 ;
        RECT -45.060 162.005 -40.125 162.170 ;
        RECT -45.060 161.520 -42.105 162.005 ;
        RECT -45.060 157.780 -43.755 161.520 ;
        RECT -42.430 161.455 -42.105 161.520 ;
        RECT -30.275 161.920 -29.795 163.250 ;
        RECT -30.275 161.900 -29.375 161.920 ;
        RECT -30.275 161.730 -28.370 161.900 ;
        RECT -30.275 161.705 -29.375 161.730 ;
        RECT -30.275 160.325 -29.795 161.705 ;
        RECT -27.950 161.635 -27.680 162.330 ;
        RECT -39.535 159.485 -39.195 159.530 ;
        RECT -39.535 159.315 -38.400 159.485 ;
        RECT -40.855 158.865 -40.660 158.870 ;
        RECT -40.865 158.205 -40.565 158.865 ;
        RECT -39.535 158.505 -39.195 159.315 ;
        RECT -39.535 158.335 -38.400 158.505 ;
        RECT -40.855 157.780 -40.660 158.205 ;
        RECT -53.845 157.555 -40.660 157.780 ;
        RECT -56.010 157.355 -54.875 157.525 ;
        RECT -55.215 155.075 -54.875 157.355 ;
        RECT -56.010 154.905 -54.875 155.075 ;
        RECT -66.605 154.510 -66.005 154.515 ;
        RECT -65.060 154.510 -64.180 154.515 ;
        RECT -66.605 154.340 -64.180 154.510 ;
        RECT -66.605 154.330 -66.005 154.340 ;
        RECT -65.060 154.320 -64.180 154.340 ;
        RECT -64.445 150.985 -64.180 154.320 ;
        RECT -55.215 154.095 -54.875 154.905 ;
        RECT -56.010 153.925 -54.875 154.095 ;
        RECT -55.215 153.115 -54.875 153.925 ;
        RECT -56.010 152.945 -54.875 153.115 ;
        RECT -55.215 152.450 -54.875 152.945 ;
        RECT -53.750 156.290 -40.660 157.555 ;
        RECT -64.615 150.965 -64.135 150.985 ;
        RECT -65.045 150.945 -64.135 150.965 ;
        RECT -66.040 150.775 -64.135 150.945 ;
        RECT -65.045 150.750 -64.135 150.775 ;
        RECT -66.730 149.135 -66.460 149.830 ;
        RECT -64.615 149.420 -64.135 150.750 ;
        RECT -65.035 149.400 -64.135 149.420 ;
        RECT -66.040 149.230 -64.135 149.400 ;
        RECT -65.035 149.205 -64.135 149.230 ;
        RECT -64.615 147.825 -64.135 149.205 ;
        RECT -53.750 149.425 -53.555 156.290 ;
        RECT -53.315 150.055 -52.975 150.550 ;
        RECT -41.435 150.055 -41.095 150.550 ;
        RECT -53.315 149.885 -52.180 150.055 ;
        RECT -42.230 149.885 -41.095 150.055 ;
        RECT -53.315 149.425 -52.975 149.885 ;
        RECT -53.750 149.075 -52.975 149.425 ;
        RECT -41.435 149.425 -41.095 149.885 ;
        RECT -40.855 149.425 -40.660 156.290 ;
        RECT -39.535 157.525 -39.195 158.335 ;
        RECT -39.535 157.355 -38.400 157.525 ;
        RECT -39.535 155.075 -39.195 157.355 ;
        RECT -39.535 154.905 -38.400 155.075 ;
        RECT -39.535 154.095 -39.195 154.905 ;
        RECT -30.230 154.515 -29.965 160.325 ;
        RECT -29.410 156.410 -28.110 156.580 ;
        RECT -28.400 156.395 -28.110 156.410 ;
        RECT -28.295 155.985 -28.110 156.395 ;
        RECT -27.920 156.245 -27.650 156.940 ;
        RECT -28.295 155.800 -27.805 155.985 ;
        RECT -27.990 154.515 -27.805 155.800 ;
        RECT -30.230 154.510 -29.350 154.515 ;
        RECT -28.405 154.510 -27.805 154.515 ;
        RECT -30.230 154.340 -27.805 154.510 ;
        RECT -30.230 154.320 -29.350 154.340 ;
        RECT -28.405 154.330 -27.805 154.340 ;
        RECT -39.535 153.925 -38.400 154.095 ;
        RECT -39.535 153.115 -39.195 153.925 ;
        RECT -39.535 152.945 -38.400 153.115 ;
        RECT -39.535 152.450 -39.195 152.945 ;
        RECT -30.230 150.985 -29.965 154.320 ;
        RECT -41.435 149.075 -40.660 149.425 ;
        RECT -53.750 148.905 -52.180 149.075 ;
        RECT -42.230 148.905 -40.660 149.075 ;
        RECT -53.750 148.870 -52.975 148.905 ;
        RECT -66.760 143.745 -66.490 144.440 ;
        RECT -66.300 143.910 -65.000 144.080 ;
        RECT -66.300 143.895 -66.010 143.910 ;
        RECT -66.300 143.485 -66.115 143.895 ;
        RECT -66.605 143.300 -66.115 143.485 ;
        RECT -66.605 142.015 -66.420 143.300 ;
        RECT -64.445 142.015 -64.180 147.825 ;
        RECT -55.215 146.360 -54.875 146.405 ;
        RECT -56.010 146.190 -54.875 146.360 ;
        RECT -55.215 145.380 -54.875 146.190 ;
        RECT -56.010 145.210 -54.875 145.380 ;
        RECT -55.215 144.400 -54.875 145.210 ;
        RECT -53.750 145.050 -53.555 148.870 ;
        RECT -53.315 148.095 -52.975 148.870 ;
        RECT -41.435 148.870 -40.660 148.905 ;
        RECT -41.435 148.095 -41.095 148.870 ;
        RECT -53.315 147.995 -52.180 148.095 ;
        RECT -53.325 147.925 -52.180 147.995 ;
        RECT -42.230 147.995 -41.095 148.095 ;
        RECT -42.230 147.925 -41.085 147.995 ;
        RECT -53.325 147.880 -52.975 147.925 ;
        RECT -41.435 147.880 -41.085 147.925 ;
        RECT -53.325 146.365 -52.985 147.880 ;
        RECT -41.425 146.365 -41.085 147.880 ;
        RECT -53.325 145.870 -52.975 146.365 ;
        RECT -41.435 145.870 -41.085 146.365 ;
        RECT -53.325 145.700 -52.180 145.870 ;
        RECT -42.230 145.700 -41.085 145.870 ;
        RECT -53.325 145.395 -52.975 145.700 ;
        RECT -56.010 144.230 -54.875 144.400 ;
        RECT -53.845 145.035 -53.545 145.050 ;
        RECT -53.315 145.035 -52.975 145.395 ;
        RECT -53.845 144.890 -52.975 145.035 ;
        RECT -41.435 145.395 -41.085 145.700 ;
        RECT -41.435 145.035 -41.095 145.395 ;
        RECT -40.855 145.050 -40.660 148.870 ;
        RECT -30.275 150.965 -29.795 150.985 ;
        RECT -30.275 150.945 -29.365 150.965 ;
        RECT -30.275 150.775 -28.370 150.945 ;
        RECT -30.275 150.750 -29.365 150.775 ;
        RECT -30.275 149.420 -29.795 150.750 ;
        RECT -30.275 149.400 -29.375 149.420 ;
        RECT -30.275 149.230 -28.370 149.400 ;
        RECT -30.275 149.205 -29.375 149.230 ;
        RECT -30.275 147.825 -29.795 149.205 ;
        RECT -27.950 149.135 -27.680 149.830 ;
        RECT -39.535 146.360 -39.195 146.405 ;
        RECT -39.535 146.190 -38.400 146.360 ;
        RECT -39.535 145.380 -39.195 146.190 ;
        RECT -39.535 145.210 -38.400 145.380 ;
        RECT -40.865 145.035 -40.565 145.050 ;
        RECT -41.435 144.890 -40.565 145.035 ;
        RECT -53.845 144.720 -52.180 144.890 ;
        RECT -42.230 144.720 -40.565 144.890 ;
        RECT -53.845 144.480 -52.975 144.720 ;
        RECT -53.845 144.365 -53.545 144.480 ;
        RECT -66.605 142.010 -66.005 142.015 ;
        RECT -65.060 142.010 -64.180 142.015 ;
        RECT -66.605 141.840 -64.180 142.010 ;
        RECT -66.605 141.830 -66.005 141.840 ;
        RECT -65.060 141.820 -64.180 141.840 ;
        RECT -64.620 138.485 -64.185 141.820 ;
        RECT -55.215 141.575 -54.875 144.230 ;
        RECT -56.010 141.405 -54.875 141.575 ;
        RECT -55.215 140.595 -54.875 141.405 ;
        RECT -56.010 140.425 -54.875 140.595 ;
        RECT -55.215 139.615 -54.875 140.425 ;
        RECT -56.010 139.445 -54.875 139.615 ;
        RECT -55.215 138.950 -54.875 139.445 ;
        RECT -64.620 138.465 -64.135 138.485 ;
        RECT -65.045 138.445 -64.135 138.465 ;
        RECT -66.040 138.275 -64.135 138.445 ;
        RECT -65.045 138.250 -64.135 138.275 ;
        RECT -64.620 137.880 -64.135 138.250 ;
        RECT -64.615 136.920 -64.135 137.880 ;
        RECT -65.035 136.900 -64.135 136.920 ;
        RECT -66.040 136.730 -64.135 136.900 ;
        RECT -65.035 136.705 -64.135 136.730 ;
        RECT -64.615 135.325 -64.135 136.705 ;
        RECT -53.750 136.045 -53.555 144.365 ;
        RECT -53.315 143.910 -52.975 144.480 ;
        RECT -41.435 144.480 -40.565 144.720 ;
        RECT -41.435 143.910 -41.095 144.480 ;
        RECT -40.865 144.365 -40.565 144.480 ;
        RECT -39.535 144.400 -39.195 145.210 ;
        RECT -53.315 143.740 -52.180 143.910 ;
        RECT -42.230 143.740 -41.095 143.910 ;
        RECT -53.315 143.695 -52.975 143.740 ;
        RECT -41.435 143.695 -41.095 143.740 ;
        RECT -53.315 136.555 -52.975 137.050 ;
        RECT -41.435 136.555 -41.095 137.050 ;
        RECT -53.315 136.385 -52.180 136.555 ;
        RECT -42.230 136.385 -41.095 136.555 ;
        RECT -53.315 136.045 -52.975 136.385 ;
        RECT -53.750 135.575 -52.975 136.045 ;
        RECT -41.435 136.045 -41.095 136.385 ;
        RECT -40.855 136.045 -40.660 144.365 ;
        RECT -39.535 144.230 -38.400 144.400 ;
        RECT -39.535 141.575 -39.195 144.230 ;
        RECT -30.230 142.015 -29.965 147.825 ;
        RECT -29.410 143.910 -28.110 144.080 ;
        RECT -28.400 143.895 -28.110 143.910 ;
        RECT -28.295 143.485 -28.110 143.895 ;
        RECT -27.920 143.745 -27.650 144.440 ;
        RECT -28.295 143.300 -27.805 143.485 ;
        RECT -27.990 142.015 -27.805 143.300 ;
        RECT -30.230 142.010 -29.350 142.015 ;
        RECT -28.405 142.010 -27.805 142.015 ;
        RECT -30.230 141.840 -27.805 142.010 ;
        RECT -30.230 141.820 -29.350 141.840 ;
        RECT -28.405 141.830 -27.805 141.840 ;
        RECT -39.535 141.405 -38.400 141.575 ;
        RECT -39.535 140.595 -39.195 141.405 ;
        RECT -39.535 140.425 -38.400 140.595 ;
        RECT -39.535 139.615 -39.195 140.425 ;
        RECT -39.535 139.445 -38.400 139.615 ;
        RECT -39.535 138.950 -39.195 139.445 ;
        RECT -30.225 138.485 -29.790 141.820 ;
        RECT -41.435 135.575 -40.660 136.045 ;
        RECT -53.750 135.490 -52.180 135.575 ;
        RECT -66.300 131.410 -65.000 131.580 ;
        RECT -66.300 131.395 -66.010 131.410 ;
        RECT -66.300 130.985 -66.115 131.395 ;
        RECT -66.605 130.800 -66.115 130.985 ;
        RECT -66.605 129.515 -66.420 130.800 ;
        RECT -64.445 129.515 -64.180 135.325 ;
        RECT -55.215 132.860 -54.875 132.905 ;
        RECT -56.010 132.690 -54.875 132.860 ;
        RECT -55.215 131.880 -54.875 132.690 ;
        RECT -53.750 132.065 -53.555 135.490 ;
        RECT -53.315 135.405 -52.180 135.490 ;
        RECT -42.230 135.490 -40.660 135.575 ;
        RECT -42.230 135.405 -41.095 135.490 ;
        RECT -53.315 134.595 -52.975 135.405 ;
        RECT -41.435 134.595 -41.095 135.405 ;
        RECT -53.315 134.425 -52.180 134.595 ;
        RECT -42.230 134.425 -41.095 134.595 ;
        RECT -53.315 132.370 -52.975 134.425 ;
        RECT -41.435 132.370 -41.095 134.425 ;
        RECT -53.315 132.200 -52.180 132.370 ;
        RECT -42.230 132.200 -41.095 132.370 ;
        RECT -56.010 131.710 -54.875 131.880 ;
        RECT -55.215 130.900 -54.875 131.710 ;
        RECT -53.815 131.990 -53.515 132.065 ;
        RECT -53.315 131.990 -52.975 132.200 ;
        RECT -53.815 131.435 -52.975 131.990 ;
        RECT -53.815 131.380 -53.515 131.435 ;
        RECT -53.315 131.390 -52.975 131.435 ;
        RECT -41.435 131.990 -41.095 132.200 ;
        RECT -40.855 132.065 -40.660 135.490 ;
        RECT -30.275 138.465 -29.790 138.485 ;
        RECT -30.275 138.445 -29.365 138.465 ;
        RECT -30.275 138.275 -28.370 138.445 ;
        RECT -30.275 138.250 -29.365 138.275 ;
        RECT -30.275 137.880 -29.790 138.250 ;
        RECT -30.275 136.920 -29.795 137.880 ;
        RECT -30.275 136.900 -29.375 136.920 ;
        RECT -30.275 136.730 -28.370 136.900 ;
        RECT -30.275 136.705 -29.375 136.730 ;
        RECT -30.275 135.325 -29.795 136.705 ;
        RECT -30.230 134.150 -29.965 135.325 ;
        RECT -30.330 133.655 -29.965 134.150 ;
        RECT -31.125 133.485 -29.965 133.655 ;
        RECT -39.535 132.860 -39.195 132.905 ;
        RECT -39.535 132.690 -38.400 132.860 ;
        RECT -40.895 131.990 -40.595 132.065 ;
        RECT -41.435 131.435 -40.595 131.990 ;
        RECT -41.435 131.390 -41.095 131.435 ;
        RECT -53.750 131.295 -53.555 131.380 ;
        RECT -56.010 130.730 -54.875 130.900 ;
        RECT -55.215 130.235 -54.875 130.730 ;
        RECT -53.315 131.220 -52.180 131.390 ;
        RECT -42.230 131.220 -41.095 131.390 ;
        RECT -40.895 131.380 -40.595 131.435 ;
        RECT -39.535 131.880 -39.195 132.690 ;
        RECT -30.330 132.675 -29.965 133.485 ;
        RECT -31.125 132.505 -29.965 132.675 ;
        RECT -39.535 131.710 -38.400 131.880 ;
        RECT -40.855 131.295 -40.660 131.380 ;
        RECT -53.315 130.410 -52.975 131.220 ;
        RECT -41.435 130.410 -41.095 131.220 ;
        RECT -53.315 130.240 -52.180 130.410 ;
        RECT -42.230 130.240 -41.095 130.410 ;
        RECT -53.315 130.195 -52.975 130.240 ;
        RECT -41.435 130.195 -41.095 130.240 ;
        RECT -39.535 130.900 -39.195 131.710 ;
        RECT -30.330 131.695 -29.965 132.505 ;
        RECT -31.125 131.525 -29.965 131.695 ;
        RECT -30.330 131.480 -29.965 131.525 ;
        RECT -39.535 130.730 -38.400 130.900 ;
        RECT -39.535 130.235 -39.195 130.730 ;
        RECT -66.605 129.510 -66.005 129.515 ;
        RECT -65.060 129.510 -64.180 129.515 ;
        RECT -66.605 129.340 -64.180 129.510 ;
        RECT -66.605 129.330 -66.005 129.340 ;
        RECT -65.060 129.320 -64.180 129.340 ;
        RECT -30.230 129.515 -29.965 131.480 ;
        RECT -29.410 131.410 -28.110 131.580 ;
        RECT -28.400 131.395 -28.110 131.410 ;
        RECT -28.295 130.985 -28.110 131.395 ;
        RECT -28.295 130.800 -27.805 130.985 ;
        RECT -27.990 129.515 -27.805 130.800 ;
        RECT -30.230 129.510 -29.350 129.515 ;
        RECT -28.405 129.510 -27.805 129.515 ;
        RECT -30.230 129.340 -27.805 129.510 ;
        RECT -30.230 129.320 -29.350 129.340 ;
        RECT -28.405 129.330 -27.805 129.340 ;
        RECT -56.100 127.945 -55.625 128.470 ;
        RECT -56.065 125.625 -55.655 127.945 ;
        RECT -56.065 125.590 -55.060 125.625 ;
        RECT -56.065 125.420 -53.590 125.590 ;
        RECT -31.395 125.490 -30.985 125.900 ;
        RECT -31.395 125.455 -30.390 125.490 ;
        RECT -56.065 125.390 -55.060 125.420 ;
        RECT -56.065 124.645 -55.655 125.390 ;
        RECT -31.395 125.285 -28.920 125.455 ;
        RECT -31.395 125.255 -30.390 125.285 ;
        RECT -56.065 124.610 -55.055 124.645 ;
        RECT -56.065 124.440 -53.590 124.610 ;
        RECT -31.395 124.510 -30.985 125.255 ;
        RECT -31.395 124.475 -30.385 124.510 ;
        RECT -56.065 124.410 -55.055 124.440 ;
        RECT -56.065 123.435 -55.655 124.410 ;
        RECT -31.395 124.305 -28.920 124.475 ;
        RECT -31.395 124.275 -30.385 124.305 ;
        RECT -56.065 123.400 -55.005 123.435 ;
        RECT -56.065 123.230 -53.590 123.400 ;
        RECT -31.395 123.300 -30.985 124.275 ;
        RECT -31.395 123.265 -30.335 123.300 ;
        RECT -56.065 123.200 -55.005 123.230 ;
        RECT -56.065 122.300 -55.655 123.200 ;
        RECT -31.395 123.095 -28.920 123.265 ;
        RECT -31.395 123.065 -30.335 123.095 ;
        RECT -31.395 122.335 -30.985 123.065 ;
        RECT -31.395 120.945 -30.980 122.335 ;
        RECT -53.880 120.115 -53.540 120.160 ;
        RECT -29.245 120.115 -28.905 120.160 ;
        RECT -54.675 119.945 -53.540 120.115 ;
        RECT -30.040 119.945 -28.905 120.115 ;
        RECT -53.880 119.135 -53.540 119.945 ;
        RECT -29.245 119.135 -28.905 119.945 ;
        RECT -54.675 118.965 -53.540 119.135 ;
        RECT -30.040 118.965 -28.905 119.135 ;
        RECT -53.880 118.155 -53.540 118.965 ;
        RECT -52.415 118.845 -52.220 118.850 ;
        RECT -52.510 118.185 -52.210 118.845 ;
        RECT -54.675 117.985 -53.540 118.155 ;
        RECT -53.880 115.705 -53.540 117.985 ;
        RECT -54.675 115.535 -53.540 115.705 ;
        RECT -53.880 114.725 -53.540 115.535 ;
        RECT -54.675 114.555 -53.540 114.725 ;
        RECT -53.880 113.745 -53.540 114.555 ;
        RECT -54.675 113.575 -53.540 113.745 ;
        RECT -53.880 113.080 -53.540 113.575 ;
        RECT -52.415 110.055 -52.220 118.185 ;
        RECT -29.245 118.155 -28.905 118.965 ;
        RECT -27.780 118.845 -27.585 118.850 ;
        RECT -27.875 118.185 -27.575 118.845 ;
        RECT -30.040 117.985 -28.905 118.155 ;
        RECT -29.245 115.705 -28.905 117.985 ;
        RECT -30.040 115.535 -28.905 115.705 ;
        RECT -29.245 114.725 -28.905 115.535 ;
        RECT -30.040 114.555 -28.905 114.725 ;
        RECT -29.245 113.745 -28.905 114.555 ;
        RECT -30.040 113.575 -28.905 113.745 ;
        RECT -29.245 113.080 -28.905 113.575 ;
        RECT -51.980 110.685 -51.640 111.180 ;
        RECT -51.980 110.515 -50.845 110.685 ;
        RECT -51.980 110.055 -51.640 110.515 ;
        RECT -52.415 109.705 -51.640 110.055 ;
        RECT -27.780 110.055 -27.585 118.185 ;
        RECT -27.345 110.685 -27.005 111.180 ;
        RECT -27.345 110.515 -26.210 110.685 ;
        RECT -27.345 110.055 -27.005 110.515 ;
        RECT -27.780 109.705 -27.005 110.055 ;
        RECT -52.415 109.535 -50.845 109.705 ;
        RECT -27.780 109.535 -26.210 109.705 ;
        RECT -52.415 109.500 -51.640 109.535 ;
        RECT -53.880 106.990 -53.540 107.035 ;
        RECT -54.675 106.820 -53.540 106.990 ;
        RECT -53.880 106.010 -53.540 106.820 ;
        RECT -54.675 105.840 -53.540 106.010 ;
        RECT -53.880 105.030 -53.540 105.840 ;
        RECT -52.415 105.680 -52.220 109.500 ;
        RECT -51.980 108.725 -51.640 109.500 ;
        RECT -27.780 109.500 -27.005 109.535 ;
        RECT -51.980 108.625 -50.845 108.725 ;
        RECT -51.990 108.555 -50.845 108.625 ;
        RECT -51.990 108.510 -51.640 108.555 ;
        RECT -51.990 106.995 -51.650 108.510 ;
        RECT -51.990 106.500 -51.640 106.995 ;
        RECT -51.990 106.330 -50.845 106.500 ;
        RECT -51.990 106.025 -51.640 106.330 ;
        RECT -54.675 104.860 -53.540 105.030 ;
        RECT -52.510 105.665 -52.210 105.680 ;
        RECT -51.980 105.665 -51.640 106.025 ;
        RECT -52.510 105.520 -51.640 105.665 ;
        RECT -45.405 105.675 -44.975 107.750 ;
        RECT -33.910 106.110 -33.345 107.435 ;
        RECT -29.245 106.990 -28.905 107.035 ;
        RECT -30.040 106.820 -28.905 106.990 ;
        RECT -34.555 106.080 -33.345 106.110 ;
        RECT -35.970 105.910 -33.345 106.080 ;
        RECT -29.245 106.010 -28.905 106.820 ;
        RECT -34.555 105.875 -33.345 105.910 ;
        RECT -52.510 105.350 -50.845 105.520 ;
        RECT -45.405 105.505 -44.195 105.675 ;
        RECT -45.405 105.350 -44.975 105.505 ;
        RECT -52.510 105.110 -51.640 105.350 ;
        RECT -52.510 104.995 -52.210 105.110 ;
        RECT -53.880 102.205 -53.540 104.860 ;
        RECT -54.675 102.035 -53.540 102.205 ;
        RECT -53.880 101.225 -53.540 102.035 ;
        RECT -54.675 101.055 -53.540 101.225 ;
        RECT -53.880 100.245 -53.540 101.055 ;
        RECT -54.675 100.075 -53.540 100.245 ;
        RECT -53.880 99.580 -53.540 100.075 ;
        RECT -52.415 96.675 -52.220 104.995 ;
        RECT -51.980 104.540 -51.640 105.110 ;
        RECT -47.745 105.045 -44.975 105.350 ;
        RECT -51.980 104.370 -50.845 104.540 ;
        RECT -51.980 104.325 -51.640 104.370 ;
        RECT -47.745 103.500 -47.440 105.045 ;
        RECT -45.405 104.695 -44.975 105.045 ;
        RECT -33.910 104.900 -33.345 105.875 ;
        RECT -30.040 105.840 -28.905 106.010 ;
        RECT -29.245 105.030 -28.905 105.840 ;
        RECT -27.780 105.680 -27.585 109.500 ;
        RECT -27.345 108.725 -27.005 109.500 ;
        RECT -27.345 108.625 -26.210 108.725 ;
        RECT -27.355 108.555 -26.210 108.625 ;
        RECT -27.355 108.510 -27.005 108.555 ;
        RECT -27.355 106.995 -27.015 108.510 ;
        RECT -27.355 106.500 -27.005 106.995 ;
        RECT -27.355 106.330 -26.210 106.500 ;
        RECT -27.355 106.025 -27.005 106.330 ;
        RECT -34.505 104.870 -33.345 104.900 ;
        RECT -35.970 104.700 -33.345 104.870 ;
        RECT -30.040 104.860 -28.905 105.030 ;
        RECT -27.875 105.665 -27.575 105.680 ;
        RECT -27.345 105.665 -27.005 106.025 ;
        RECT -27.875 105.520 -27.005 105.665 ;
        RECT -27.875 105.350 -26.210 105.520 ;
        RECT -27.875 105.110 -27.005 105.350 ;
        RECT -27.875 104.995 -27.575 105.110 ;
        RECT -45.405 104.525 -44.195 104.695 ;
        RECT -34.505 104.665 -33.345 104.700 ;
        RECT -45.405 103.825 -44.975 104.525 ;
        RECT -33.910 103.920 -33.345 104.665 ;
        RECT -34.500 103.890 -33.345 103.920 ;
        RECT -35.970 103.720 -33.345 103.890 ;
        RECT -34.500 103.685 -33.345 103.720 ;
        RECT -47.885 103.100 -47.440 103.500 ;
        RECT -47.885 101.650 -47.455 103.100 ;
        RECT -47.885 101.480 -45.730 101.650 ;
        RECT -47.885 101.475 -47.270 101.480 ;
        RECT -47.885 100.605 -47.455 101.475 ;
        RECT -38.155 100.680 -37.725 101.905 ;
        RECT -47.885 100.175 -46.620 100.605 ;
        RECT -38.935 100.510 -37.725 100.680 ;
        RECT -47.050 97.765 -46.620 100.175 ;
        RECT -38.155 100.355 -37.725 100.510 ;
        RECT -33.910 100.355 -33.345 103.685 ;
        RECT -29.245 102.205 -28.905 104.860 ;
        RECT -30.040 102.035 -28.905 102.205 ;
        RECT -29.245 101.225 -28.905 102.035 ;
        RECT -30.040 101.055 -28.905 101.225 ;
        RECT -38.155 100.050 -33.345 100.355 ;
        RECT -29.245 100.245 -28.905 101.055 ;
        RECT -30.040 100.075 -28.905 100.245 ;
        RECT -38.155 99.700 -37.725 100.050 ;
        RECT -38.935 99.530 -37.725 99.700 ;
        RECT -38.155 98.830 -37.725 99.530 ;
        RECT -35.690 98.140 -35.385 100.050 ;
        RECT -29.245 99.580 -28.905 100.075 ;
        RECT -35.690 98.105 -35.295 98.140 ;
        RECT -51.980 97.185 -51.640 97.680 ;
        RECT -47.050 97.595 -45.340 97.765 ;
        RECT -51.980 97.015 -50.845 97.185 ;
        RECT -51.980 96.675 -51.640 97.015 ;
        RECT -52.415 96.205 -51.640 96.675 ;
        RECT -47.050 96.785 -46.620 97.595 ;
        RECT -47.050 96.615 -45.340 96.785 ;
        RECT -35.600 96.655 -35.295 98.105 ;
        RECT -52.415 96.120 -50.845 96.205 ;
        RECT -53.880 93.490 -53.540 93.535 ;
        RECT -54.675 93.320 -53.540 93.490 ;
        RECT -53.880 92.510 -53.540 93.320 ;
        RECT -52.415 92.695 -52.220 96.120 ;
        RECT -51.980 96.035 -50.845 96.120 ;
        RECT -51.980 95.225 -51.640 96.035 ;
        RECT -47.050 95.915 -46.620 96.615 ;
        RECT -37.400 96.485 -35.295 96.655 ;
        RECT -35.860 96.480 -35.295 96.485 ;
        RECT -35.600 95.895 -35.295 96.480 ;
        RECT -27.780 96.675 -27.585 104.995 ;
        RECT -27.345 104.540 -27.005 105.110 ;
        RECT -27.345 104.370 -26.210 104.540 ;
        RECT -27.345 104.325 -27.005 104.370 ;
        RECT -27.345 97.185 -27.005 97.680 ;
        RECT -27.345 97.015 -26.210 97.185 ;
        RECT -27.345 96.675 -27.005 97.015 ;
        RECT -27.780 96.205 -27.005 96.675 ;
        RECT -27.780 96.120 -26.210 96.205 ;
        RECT -51.980 95.055 -50.845 95.225 ;
        RECT -51.980 93.000 -51.640 95.055 ;
        RECT -29.245 93.490 -28.905 93.535 ;
        RECT -30.040 93.320 -28.905 93.490 ;
        RECT -51.980 92.830 -50.845 93.000 ;
        RECT -54.675 92.340 -53.540 92.510 ;
        RECT -53.880 91.530 -53.540 92.340 ;
        RECT -52.480 92.620 -52.180 92.695 ;
        RECT -51.980 92.620 -51.640 92.830 ;
        RECT -52.480 92.065 -51.640 92.620 ;
        RECT -29.245 92.510 -28.905 93.320 ;
        RECT -27.780 92.695 -27.585 96.120 ;
        RECT -27.345 96.035 -26.210 96.120 ;
        RECT -27.345 95.225 -27.005 96.035 ;
        RECT -27.345 95.055 -26.210 95.225 ;
        RECT -27.345 93.000 -27.005 95.055 ;
        RECT -27.345 92.830 -26.210 93.000 ;
        RECT -30.040 92.340 -28.905 92.510 ;
        RECT -52.480 92.010 -52.180 92.065 ;
        RECT -51.980 92.020 -51.640 92.065 ;
        RECT -52.415 91.925 -52.220 92.010 ;
        RECT -54.675 91.360 -53.540 91.530 ;
        RECT -53.880 90.865 -53.540 91.360 ;
        RECT -51.980 91.850 -50.845 92.020 ;
        RECT -51.980 91.040 -51.640 91.850 ;
        RECT -29.245 91.530 -28.905 92.340 ;
        RECT -27.845 92.620 -27.545 92.695 ;
        RECT -27.345 92.620 -27.005 92.830 ;
        RECT -27.845 92.065 -27.005 92.620 ;
        RECT -27.845 92.010 -27.545 92.065 ;
        RECT -27.345 92.020 -27.005 92.065 ;
        RECT -27.780 91.925 -27.585 92.010 ;
        RECT -30.040 91.360 -28.905 91.530 ;
        RECT -51.980 90.870 -50.845 91.040 ;
        RECT -51.980 90.825 -51.640 90.870 ;
        RECT -29.245 90.865 -28.905 91.360 ;
        RECT -27.345 91.850 -26.210 92.020 ;
        RECT -27.345 91.040 -27.005 91.850 ;
        RECT -27.345 90.870 -26.210 91.040 ;
        RECT -27.345 90.825 -27.005 90.870 ;
        RECT -65.525 80.730 -65.095 82.805 ;
        RECT -54.030 81.165 -53.465 82.490 ;
        RECT -54.675 81.135 -53.465 81.165 ;
        RECT -56.090 80.965 -53.465 81.135 ;
        RECT -54.675 80.930 -53.465 80.965 ;
        RECT -65.525 80.560 -64.315 80.730 ;
        RECT -65.525 80.405 -65.095 80.560 ;
        RECT -67.865 80.100 -65.095 80.405 ;
        RECT -67.865 78.555 -67.560 80.100 ;
        RECT -65.525 79.750 -65.095 80.100 ;
        RECT -54.030 79.955 -53.465 80.930 ;
        RECT -40.525 80.730 -40.095 82.805 ;
        RECT -29.030 81.165 -28.465 82.490 ;
        RECT -29.675 81.135 -28.465 81.165 ;
        RECT -31.090 80.965 -28.465 81.135 ;
        RECT -29.675 80.930 -28.465 80.965 ;
        RECT -40.525 80.560 -39.315 80.730 ;
        RECT -40.525 80.405 -40.095 80.560 ;
        RECT -54.625 79.925 -53.465 79.955 ;
        RECT -56.090 79.755 -53.465 79.925 ;
        RECT -65.525 79.580 -64.315 79.750 ;
        RECT -54.625 79.720 -53.465 79.755 ;
        RECT -65.525 78.880 -65.095 79.580 ;
        RECT -54.030 78.975 -53.465 79.720 ;
        RECT -54.620 78.945 -53.465 78.975 ;
        RECT -56.090 78.775 -53.465 78.945 ;
        RECT -54.620 78.740 -53.465 78.775 ;
        RECT -68.005 78.155 -67.560 78.555 ;
        RECT -68.005 76.705 -67.575 78.155 ;
        RECT -68.005 76.535 -65.850 76.705 ;
        RECT -68.005 76.530 -67.390 76.535 ;
        RECT -68.005 75.660 -67.575 76.530 ;
        RECT -58.275 75.735 -57.845 76.960 ;
        RECT -68.005 75.230 -66.740 75.660 ;
        RECT -59.055 75.565 -57.845 75.735 ;
        RECT -67.170 72.820 -66.740 75.230 ;
        RECT -58.275 75.410 -57.845 75.565 ;
        RECT -54.030 75.410 -53.465 78.740 ;
        RECT -42.865 80.100 -40.095 80.405 ;
        RECT -42.865 78.555 -42.560 80.100 ;
        RECT -40.525 79.750 -40.095 80.100 ;
        RECT -29.030 79.955 -28.465 80.930 ;
        RECT -29.625 79.925 -28.465 79.955 ;
        RECT -31.090 79.755 -28.465 79.925 ;
        RECT -40.525 79.580 -39.315 79.750 ;
        RECT -29.625 79.720 -28.465 79.755 ;
        RECT -40.525 78.880 -40.095 79.580 ;
        RECT -29.030 78.975 -28.465 79.720 ;
        RECT -29.620 78.945 -28.465 78.975 ;
        RECT -31.090 78.775 -28.465 78.945 ;
        RECT -29.620 78.740 -28.465 78.775 ;
        RECT -43.005 78.155 -42.560 78.555 ;
        RECT -43.005 76.705 -42.575 78.155 ;
        RECT -43.005 76.535 -40.850 76.705 ;
        RECT -43.005 76.530 -42.390 76.535 ;
        RECT -43.005 76.460 -42.575 76.530 ;
        RECT -58.275 75.105 -53.465 75.410 ;
        RECT -44.085 75.660 -42.575 76.460 ;
        RECT -33.275 75.735 -32.845 76.960 ;
        RECT -44.085 75.410 -41.740 75.660 ;
        RECT -34.055 75.565 -32.845 75.735 ;
        RECT -58.275 74.755 -57.845 75.105 ;
        RECT -59.055 74.585 -57.845 74.755 ;
        RECT -58.275 73.885 -57.845 74.585 ;
        RECT -55.810 73.195 -55.505 75.105 ;
        RECT -67.170 72.650 -65.460 72.820 ;
        RECT -67.170 71.840 -66.740 72.650 ;
        RECT -67.170 71.670 -65.460 71.840 ;
        RECT -55.810 71.710 -55.415 73.195 ;
        RECT -67.170 70.970 -66.740 71.670 ;
        RECT -57.520 71.540 -55.415 71.710 ;
        RECT -55.980 71.535 -55.415 71.540 ;
        RECT -55.810 70.950 -55.415 71.535 ;
        RECT -55.810 68.695 -55.505 70.950 ;
        RECT -57.905 68.390 -55.505 68.695 ;
        RECT -59.480 66.760 -59.035 66.850 ;
        RECT -57.905 66.760 -57.600 68.390 ;
        RECT -59.480 66.455 -57.600 66.760 ;
        RECT -44.085 67.845 -43.310 75.410 ;
        RECT -43.005 75.230 -41.740 75.410 ;
        RECT -42.170 72.820 -41.740 75.230 ;
        RECT -33.275 75.410 -32.845 75.565 ;
        RECT -29.030 75.410 -28.465 78.740 ;
        RECT -33.275 75.105 -28.465 75.410 ;
        RECT -33.275 74.755 -32.845 75.105 ;
        RECT -34.055 74.585 -32.845 74.755 ;
        RECT -33.275 73.885 -32.845 74.585 ;
        RECT -30.810 73.195 -30.505 75.105 ;
        RECT -42.170 72.650 -40.460 72.820 ;
        RECT -42.170 71.840 -41.740 72.650 ;
        RECT -42.170 71.670 -40.460 71.840 ;
        RECT -30.810 71.710 -30.415 73.195 ;
        RECT -42.170 70.970 -41.740 71.670 ;
        RECT -32.520 71.540 -30.415 71.710 ;
        RECT -30.980 71.535 -30.415 71.540 ;
        RECT -30.810 70.950 -30.415 71.535 ;
        RECT -30.810 68.875 -30.505 70.950 ;
        RECT -31.225 68.570 -30.505 68.875 ;
        RECT -44.085 67.675 -41.465 67.845 ;
        RECT -44.085 66.670 -43.310 67.675 ;
        RECT -31.215 67.555 -30.785 68.570 ;
        RECT -31.215 67.385 -30.005 67.555 ;
        RECT -34.080 67.230 -33.320 67.380 ;
        RECT -31.215 67.230 -30.785 67.385 ;
        RECT -34.080 66.925 -30.785 67.230 ;
        RECT -59.480 65.770 -59.035 66.455 ;
        RECT -59.785 65.700 -59.035 65.770 ;
        RECT -59.785 65.680 -58.280 65.700 ;
        RECT -59.785 65.510 -57.480 65.680 ;
        RECT -59.785 65.480 -58.280 65.510 ;
        RECT -59.785 64.730 -59.035 65.480 ;
        RECT -56.905 65.175 -56.605 65.890 ;
        RECT -59.785 64.700 -58.275 64.730 ;
        RECT -59.785 64.530 -57.480 64.700 ;
        RECT -59.785 64.510 -58.275 64.530 ;
        RECT -59.785 63.865 -59.035 64.510 ;
        RECT -57.305 64.060 -57.005 64.790 ;
        RECT -57.265 63.870 -57.085 64.060 ;
        RECT -63.250 63.550 -62.565 63.840 ;
        RECT -63.980 58.110 -63.655 58.600 ;
        RECT -66.465 57.940 -63.655 58.110 ;
        RECT -63.980 57.125 -63.655 57.940 ;
        RECT -64.075 52.950 -63.500 57.125 ;
        RECT -65.960 52.780 -63.500 52.950 ;
        RECT -64.075 52.210 -63.500 52.780 ;
        RECT -77.480 42.775 -76.775 51.860 ;
        RECT -63.250 51.290 -63.045 63.550 ;
        RECT -63.730 51.000 -63.045 51.290 ;
        RECT -62.865 63.085 -62.180 63.375 ;
        RECT -62.865 50.565 -62.660 63.085 ;
        RECT -59.785 62.325 -59.205 63.865 ;
        RECT -57.710 63.580 -57.025 63.870 ;
        RECT -56.820 63.485 -56.640 65.175 ;
        RECT -56.850 63.195 -56.165 63.485 ;
        RECT -44.085 62.685 -43.445 66.670 ;
        RECT -34.080 64.980 -33.250 66.925 ;
        RECT -31.215 66.575 -30.785 66.925 ;
        RECT -31.215 66.405 -30.005 66.575 ;
        RECT -31.215 65.705 -30.785 66.405 ;
        RECT -34.080 63.530 -33.320 64.980 ;
        RECT -34.080 63.360 -31.540 63.530 ;
        RECT -34.080 63.355 -33.080 63.360 ;
        RECT -44.085 62.515 -40.960 62.685 ;
        RECT -59.785 61.175 -59.030 62.325 ;
        RECT -44.085 62.025 -43.445 62.515 ;
        RECT -59.785 61.155 -58.275 61.175 ;
        RECT -59.785 60.985 -57.475 61.155 ;
        RECT -44.085 61.115 -43.460 62.025 ;
        RECT -35.065 61.145 -34.405 61.410 ;
        RECT -59.785 60.955 -58.275 60.985 ;
        RECT -59.785 60.205 -59.030 60.955 ;
        RECT -44.085 60.540 -42.795 61.115 ;
        RECT -59.785 60.175 -58.270 60.205 ;
        RECT -59.785 60.005 -57.475 60.175 ;
        RECT -59.785 59.985 -58.270 60.005 ;
        RECT -59.785 59.340 -59.030 59.985 ;
        RECT -57.300 59.535 -57.000 60.265 ;
        RECT -62.470 58.980 -61.785 59.270 ;
        RECT -63.340 50.275 -62.655 50.565 ;
        RECT -62.470 49.995 -62.265 58.980 ;
        RECT -61.305 57.295 -60.775 57.715 ;
        RECT -61.440 57.145 -60.690 57.295 ;
        RECT -59.785 57.145 -59.205 59.340 ;
        RECT -57.260 59.280 -57.080 59.535 ;
        RECT -57.700 58.990 -57.015 59.280 ;
        RECT -61.440 56.565 -59.205 57.145 ;
        RECT -43.370 57.520 -42.795 60.540 ;
        RECT -40.760 57.845 -40.330 59.070 ;
        RECT -40.760 57.675 -39.550 57.845 ;
        RECT -40.760 57.520 -40.330 57.675 ;
        RECT -43.370 57.215 -40.330 57.520 ;
        RECT -61.440 55.160 -60.690 56.565 ;
        RECT -43.370 55.270 -42.795 57.215 ;
        RECT -40.760 56.865 -40.330 57.215 ;
        RECT -40.760 56.695 -39.550 56.865 ;
        RECT -40.760 55.995 -40.330 56.695 ;
        RECT -43.370 55.265 -42.885 55.270 ;
        RECT -61.440 55.125 -60.030 55.160 ;
        RECT -61.440 54.955 -59.190 55.125 ;
        RECT -61.440 54.920 -60.030 54.955 ;
        RECT -61.440 54.190 -60.690 54.920 ;
        RECT -61.440 54.145 -60.045 54.190 ;
        RECT -61.440 53.975 -59.190 54.145 ;
        RECT -61.440 53.950 -60.045 53.975 ;
        RECT -61.440 53.275 -60.690 53.950 ;
        RECT -43.190 53.820 -42.885 55.265 ;
        RECT -40.900 55.060 -40.545 55.430 ;
        RECT -43.190 53.650 -41.085 53.820 ;
        RECT -43.190 53.645 -42.625 53.650 ;
        RECT -43.190 53.060 -42.885 53.645 ;
        RECT -40.870 53.355 -40.675 55.060 ;
        RECT -40.875 53.005 -40.675 53.355 ;
        RECT -40.875 53.000 -40.665 53.005 ;
        RECT -42.575 50.570 -41.390 50.585 ;
        RECT -40.865 50.570 -40.665 53.000 ;
        RECT -40.425 52.735 -40.155 53.410 ;
        RECT -40.385 52.635 -40.185 52.735 ;
        RECT -40.375 51.300 -40.195 52.635 ;
        RECT -40.385 51.000 -39.200 51.300 ;
        RECT -42.575 50.370 -40.665 50.570 ;
        RECT -42.575 50.285 -41.390 50.370 ;
        RECT -35.065 50.010 -34.885 61.145 ;
        RECT -34.080 59.245 -33.320 63.355 ;
        RECT -30.880 62.445 -30.610 63.120 ;
        RECT -30.840 62.345 -30.640 62.445 ;
        RECT -30.830 61.980 -30.650 62.345 ;
        RECT -30.855 61.295 -30.565 61.980 ;
        RECT -34.090 58.695 -33.320 59.245 ;
        RECT -34.090 58.525 -31.785 58.695 ;
        RECT -34.090 57.600 -33.320 58.525 ;
        RECT -34.090 53.535 -33.765 57.600 ;
        RECT -34.090 53.365 -31.280 53.535 ;
        RECT -34.090 52.875 -33.765 53.365 ;
        RECT -62.935 49.705 -62.250 49.995 ;
        RECT -35.075 49.705 -33.995 50.010 ;
        RECT -80.910 41.050 -76.775 42.775 ;
        RECT -10.525 42.720 -3.730 221.290 ;
        RECT 84.745 65.025 86.410 84.195 ;
        RECT 84.745 56.750 86.575 65.025 ;
        RECT 85.625 51.250 86.575 56.750 ;
        RECT 85.590 50.860 86.685 51.250 ;
        RECT 80.070 50.690 81.110 50.860 ;
        RECT 84.070 50.690 86.685 50.860 ;
        RECT 85.590 48.280 86.685 50.690 ;
        RECT 346.220 50.060 461.680 50.230 ;
        RECT 346.220 48.410 346.390 50.060 ;
        RECT 461.510 48.410 461.680 50.060 ;
        RECT 346.220 48.340 461.680 48.410 ;
        RECT 80.070 48.110 81.110 48.280 ;
        RECT 84.070 48.110 86.685 48.280 ;
        RECT 85.590 45.700 86.685 48.110 ;
        RECT 80.070 45.530 81.110 45.700 ;
        RECT 84.070 45.530 86.685 45.700 ;
        RECT 80.145 44.860 80.605 45.030 ;
        RECT 85.590 44.540 86.685 45.530 ;
        RECT 346.215 48.240 461.680 48.340 ;
        RECT -80.910 40.220 -76.835 41.050 ;
        RECT -33.235 35.925 -3.725 42.720 ;
        RECT 85.625 41.705 86.575 44.540 ;
        RECT 346.215 44.390 461.555 48.240 ;
        RECT 88.355 41.705 461.555 44.390 ;
        RECT 85.625 40.755 461.555 41.705 ;
        RECT 88.355 38.230 461.555 40.755 ;
        RECT 133.765 38.115 190.365 38.230 ;
        RECT -10.525 22.755 -3.730 35.925 ;
        RECT 14.330 22.755 16.250 22.800 ;
        RECT 40.900 22.755 41.070 32.235 ;
        RECT 49.480 22.755 49.650 32.235 ;
        RECT 58.060 23.215 58.230 32.235 ;
        RECT 58.060 22.755 58.235 23.215 ;
        RECT -10.985 20.425 63.270 22.755 ;
        RECT 127.865 18.890 131.960 18.895 ;
        RECT 132.915 18.890 194.330 19.430 ;
        RECT 127.865 17.420 238.370 18.890 ;
        RECT 97.835 14.385 98.160 14.390 ;
        RECT 97.815 14.000 98.180 14.385 ;
        RECT 98.970 14.220 99.140 15.010 ;
        RECT 99.950 14.220 100.120 15.010 ;
        RECT 100.930 14.220 101.100 15.010 ;
        RECT 98.970 14.215 101.505 14.220 ;
        RECT 103.220 14.215 103.390 15.010 ;
        RECT 104.200 14.215 104.370 15.010 ;
        RECT 105.180 14.215 105.350 15.010 ;
        RECT 14.100 11.835 15.495 12.540 ;
        RECT 2.825 11.370 15.495 11.835 ;
        RECT 2.825 11.360 14.825 11.370 ;
        RECT 2.955 10.860 3.960 11.360 ;
        RECT 3.565 9.985 3.735 10.860 ;
        RECT 6.125 9.930 6.295 11.360 ;
        RECT 7.575 9.955 7.745 11.360 ;
        RECT 12.275 10.860 14.825 11.360 ;
        RECT 9.735 9.990 9.905 10.630 ;
        RECT 10.915 9.990 11.085 10.630 ;
        RECT 12.500 9.985 12.670 10.860 ;
        RECT 14.045 9.985 14.215 10.860 ;
        RECT 22.575 8.390 22.745 9.185 ;
        RECT 23.555 8.390 23.725 9.185 ;
        RECT 24.535 8.390 24.705 9.185 ;
        RECT 26.825 8.390 26.995 9.185 ;
        RECT 27.805 8.390 27.975 9.185 ;
        RECT 28.785 8.390 28.955 9.185 ;
        RECT 22.530 8.050 29.450 8.390 ;
        RECT 23.130 7.585 23.840 8.050 ;
        RECT 3.565 3.450 3.735 4.325 ;
        RECT 2.955 2.950 3.960 3.450 ;
        RECT 6.125 2.950 6.295 4.380 ;
        RECT 7.575 2.950 7.745 4.355 ;
        RECT 9.735 3.680 9.905 4.320 ;
        RECT 10.915 3.680 11.085 4.320 ;
        RECT 12.500 3.450 12.670 4.325 ;
        RECT 14.045 3.450 14.215 4.325 ;
        RECT 12.275 2.965 14.825 3.450 ;
        RECT 20.980 2.975 21.630 7.520 ;
        RECT 23.000 6.960 24.085 7.585 ;
        RECT 26.780 7.365 29.450 8.050 ;
        RECT 57.840 7.585 75.250 7.725 ;
        RECT 26.825 6.570 26.995 7.365 ;
        RECT 27.805 6.570 27.975 7.365 ;
        RECT 28.785 6.570 28.955 7.365 ;
        RECT 57.100 7.265 75.250 7.585 ;
        RECT 39.550 4.800 39.720 7.265 ;
        RECT 40.730 4.800 40.900 7.265 ;
        RECT 41.910 4.800 42.080 7.265 ;
        RECT 43.090 4.800 43.260 7.265 ;
        RECT 44.270 4.800 44.440 7.265 ;
        RECT 45.450 4.800 45.620 7.265 ;
        RECT 46.630 4.800 46.800 7.265 ;
        RECT 47.810 4.855 47.980 7.265 ;
        RECT 46.970 4.800 48.810 4.855 ;
        RECT 48.990 4.800 49.160 7.265 ;
        RECT 50.170 4.800 50.340 7.265 ;
        RECT 51.350 4.800 51.520 7.265 ;
        RECT 52.530 4.800 52.700 7.265 ;
        RECT 53.710 4.800 53.880 7.265 ;
        RECT 54.890 4.800 55.060 7.265 ;
        RECT 56.070 4.800 56.240 7.265 ;
        RECT 57.250 4.800 57.420 7.265 ;
        RECT 57.840 5.225 58.010 7.265 ;
        RECT 58.430 5.225 58.600 7.265 ;
        RECT 59.020 5.225 59.190 7.265 ;
        RECT 59.610 5.225 59.780 7.265 ;
        RECT 60.200 5.225 60.370 7.265 ;
        RECT 60.790 5.225 60.960 7.265 ;
        RECT 61.380 5.225 61.550 7.265 ;
        RECT 61.970 5.225 62.140 7.265 ;
        RECT 62.560 5.225 62.730 7.265 ;
        RECT 63.150 5.225 63.320 7.265 ;
        RECT 63.740 5.225 63.910 7.265 ;
        RECT 64.330 5.225 64.500 7.265 ;
        RECT 64.920 5.225 65.090 7.265 ;
        RECT 65.510 5.225 65.680 7.265 ;
        RECT 66.100 5.225 66.270 7.265 ;
        RECT 66.690 5.225 66.860 7.265 ;
        RECT 67.280 5.225 67.450 7.265 ;
        RECT 67.870 5.225 68.040 7.265 ;
        RECT 68.460 5.225 68.630 7.265 ;
        RECT 69.050 5.225 69.220 7.265 ;
        RECT 69.640 5.225 69.810 7.265 ;
        RECT 70.230 5.225 70.400 7.265 ;
        RECT 70.820 5.225 70.990 7.265 ;
        RECT 71.410 5.225 71.580 7.265 ;
        RECT 72.000 5.225 72.170 7.265 ;
        RECT 72.590 5.225 72.760 7.265 ;
        RECT 73.180 5.225 73.350 7.265 ;
        RECT 73.770 5.225 73.940 7.265 ;
        RECT 74.360 5.225 74.530 7.265 ;
        RECT 74.950 5.225 75.120 7.265 ;
        RECT 97.835 6.210 98.160 14.000 ;
        RECT 98.925 13.875 105.845 14.215 ;
        RECT 103.175 13.190 105.845 13.875 ;
        RECT 103.220 12.395 103.390 13.190 ;
        RECT 104.200 12.395 104.370 13.190 ;
        RECT 105.180 12.395 105.350 13.190 ;
        RECT 127.865 6.780 129.340 17.420 ;
        RECT 131.445 17.415 238.370 17.420 ;
        RECT 151.525 13.445 158.205 13.895 ;
        RECT 166.495 13.445 168.525 17.415 ;
        RECT 175.200 13.445 181.880 14.005 ;
        RECT 151.525 13.380 181.880 13.445 ;
        RECT 151.525 13.270 175.495 13.380 ;
        RECT 151.650 10.460 151.820 13.270 ;
        RECT 153.230 10.460 153.400 13.270 ;
        RECT 154.810 10.460 154.980 13.270 ;
        RECT 155.600 10.370 155.770 12.500 ;
        RECT 156.390 10.370 156.560 13.270 ;
        RECT 157.970 12.820 175.495 13.270 ;
        RECT 157.180 10.370 157.350 12.500 ;
        RECT 157.970 10.370 158.140 12.820 ;
        RECT 175.325 10.570 175.495 12.820 ;
        RECT 176.905 10.570 177.075 13.380 ;
        RECT 178.485 10.570 178.655 13.380 ;
        RECT 155.600 10.200 158.140 10.370 ;
        RECT 179.275 10.480 179.445 12.610 ;
        RECT 180.065 10.480 180.235 13.380 ;
        RECT 181.645 13.205 181.815 13.380 ;
        RECT 183.805 13.220 190.485 13.790 ;
        RECT 183.805 13.205 194.690 13.220 ;
        RECT 181.645 13.165 194.690 13.205 ;
        RECT 181.645 12.740 184.100 13.165 ;
        RECT 180.855 10.480 181.025 12.610 ;
        RECT 181.645 10.480 181.815 12.740 ;
        RECT 179.275 10.310 181.815 10.480 ;
        RECT 183.930 10.355 184.100 12.740 ;
        RECT 185.510 10.355 185.680 13.165 ;
        RECT 187.090 10.355 187.260 13.165 ;
        RECT 155.845 9.935 157.860 10.200 ;
        RECT 179.520 10.045 181.535 10.310 ;
        RECT 187.880 10.265 188.050 12.395 ;
        RECT 188.670 10.265 188.840 13.165 ;
        RECT 190.250 12.740 194.690 13.165 ;
        RECT 189.460 10.265 189.630 12.395 ;
        RECT 190.250 10.265 190.420 12.740 ;
        RECT 194.370 12.035 194.690 12.740 ;
        RECT 193.900 10.745 194.860 12.035 ;
        RECT 195.930 12.000 196.100 12.795 ;
        RECT 196.910 12.000 197.080 12.795 ;
        RECT 197.890 12.000 198.060 12.795 ;
        RECT 200.340 12.000 200.510 12.795 ;
        RECT 201.320 12.000 201.490 12.795 ;
        RECT 202.300 12.000 202.470 12.795 ;
        RECT 209.055 12.000 209.225 12.795 ;
        RECT 210.035 12.000 210.205 12.795 ;
        RECT 211.015 12.000 211.185 12.795 ;
        RECT 213.840 12.000 214.010 12.795 ;
        RECT 214.820 12.000 214.990 12.795 ;
        RECT 215.800 12.000 215.970 12.795 ;
        RECT 222.555 12.000 222.725 12.795 ;
        RECT 223.535 12.000 223.705 12.795 ;
        RECT 224.515 12.000 224.685 12.795 ;
        RECT 195.885 11.660 202.965 12.000 ;
        RECT 209.010 11.660 216.465 12.000 ;
        RECT 222.510 11.660 225.180 12.000 ;
        RECT 229.020 11.275 229.750 12.205 ;
        RECT 197.200 10.535 197.860 10.630 ;
        RECT 210.365 10.535 211.050 10.630 ;
        RECT 223.350 10.535 224.035 10.600 ;
        RECT 229.265 10.550 229.485 11.275 ;
        RECT 197.195 10.340 224.120 10.535 ;
        RECT 197.200 10.330 197.860 10.340 ;
        RECT 187.880 10.095 190.420 10.265 ;
        RECT 205.990 10.100 206.545 10.340 ;
        RECT 210.365 10.330 211.050 10.340 ;
        RECT 207.420 10.100 210.020 10.110 ;
        RECT 210.380 10.100 210.935 10.330 ;
        RECT 219.370 10.100 219.925 10.340 ;
        RECT 223.350 10.300 224.035 10.340 ;
        RECT 223.425 10.100 223.980 10.300 ;
        RECT 227.850 10.210 230.520 10.550 ;
        RECT 188.125 9.830 190.140 10.095 ;
        RECT 204.865 9.770 211.720 10.100 ;
        RECT 204.865 9.760 207.535 9.770 ;
        RECT 209.050 9.760 211.720 9.770 ;
        RECT 218.365 9.760 225.220 10.100 ;
        RECT 205.360 8.965 205.530 9.760 ;
        RECT 206.340 8.965 206.510 9.760 ;
        RECT 207.320 8.965 207.490 9.760 ;
        RECT 209.545 8.965 209.715 9.760 ;
        RECT 210.525 8.965 210.695 9.760 ;
        RECT 211.505 8.965 211.675 9.760 ;
        RECT 218.860 8.965 219.030 9.760 ;
        RECT 219.840 8.965 220.010 9.760 ;
        RECT 220.820 8.965 220.990 9.760 ;
        RECT 223.045 8.965 223.215 9.760 ;
        RECT 224.025 8.965 224.195 9.760 ;
        RECT 225.005 8.965 225.175 9.760 ;
        RECT 227.895 9.415 228.065 10.210 ;
        RECT 228.875 9.415 229.045 10.210 ;
        RECT 229.855 9.415 230.025 10.210 ;
        RECT 97.020 6.205 98.680 6.210 ;
        RECT 39.340 4.200 75.275 4.800 ;
        RECT 97.020 4.715 98.850 6.205 ;
        RECT 41.015 3.720 42.855 4.200 ;
        RECT 46.970 3.720 48.810 4.200 ;
        RECT 53.200 3.720 55.040 4.200 ;
        RECT 61.020 3.720 62.860 4.200 ;
        RECT 66.645 3.720 68.485 4.200 ;
        RECT 72.490 3.720 74.330 4.200 ;
        RECT 97.020 3.720 98.710 4.715 ;
        RECT 112.095 4.380 129.340 6.780 ;
        RECT 139.080 4.685 139.250 5.725 ;
        RECT 139.870 4.685 140.040 5.725 ;
        RECT 40.445 2.975 98.710 3.720 ;
        RECT 15.150 2.965 98.710 2.975 ;
        RECT 12.275 2.950 98.710 2.965 ;
        RECT 2.825 2.475 98.710 2.950 ;
        RECT 13.820 1.910 98.710 2.475 ;
        RECT 13.820 1.680 15.495 1.910 ;
        RECT 99.830 -2.535 100.000 -1.740 ;
        RECT 100.810 -2.535 100.980 -1.740 ;
        RECT 101.790 -2.535 101.960 -1.740 ;
        RECT 104.080 -2.535 104.250 -1.740 ;
        RECT 105.060 -2.535 105.230 -1.740 ;
        RECT 106.040 -2.535 106.210 -1.740 ;
        RECT 99.785 -2.875 106.705 -2.535 ;
        RECT 104.035 -3.560 106.705 -2.875 ;
        RECT 22.650 -5.060 22.820 -4.265 ;
        RECT 23.630 -5.060 23.800 -4.265 ;
        RECT 24.610 -5.060 24.780 -4.265 ;
        RECT 26.900 -5.060 27.070 -4.265 ;
        RECT 27.880 -5.060 28.050 -4.265 ;
        RECT 28.860 -5.060 29.030 -4.265 ;
        RECT 104.080 -4.355 104.250 -3.560 ;
        RECT 105.060 -4.355 105.230 -3.560 ;
        RECT 106.040 -4.355 106.210 -3.560 ;
        RECT 22.605 -5.400 29.525 -5.060 ;
        RECT 26.855 -6.085 29.525 -5.400 ;
        RECT 127.865 -5.775 129.340 4.380 ;
        RECT 145.610 4.290 145.780 5.705 ;
        RECT 146.400 4.290 146.570 5.705 ;
        RECT 163.355 4.650 163.525 5.690 ;
        RECT 164.145 4.650 164.315 5.690 ;
        RECT 145.505 3.885 146.680 4.290 ;
        RECT 169.885 4.255 170.055 5.670 ;
        RECT 170.675 4.255 170.845 5.670 ;
        RECT 139.080 2.430 139.250 3.465 ;
        RECT 139.870 2.430 140.040 3.465 ;
        RECT 139.080 2.015 140.040 2.430 ;
        RECT 145.605 2.425 145.775 3.885 ;
        RECT 146.395 2.425 146.565 3.885 ;
        RECT 169.780 3.850 170.955 4.255 ;
        RECT 236.895 4.120 238.370 17.415 ;
        RECT 274.230 11.470 291.640 11.610 ;
        RECT 273.490 11.150 291.640 11.470 ;
        RECT 255.940 8.685 256.110 11.150 ;
        RECT 257.120 8.685 257.290 11.150 ;
        RECT 258.300 8.685 258.470 11.150 ;
        RECT 259.480 8.685 259.650 11.150 ;
        RECT 260.660 8.685 260.830 11.150 ;
        RECT 261.840 8.685 262.010 11.150 ;
        RECT 263.020 8.685 263.190 11.150 ;
        RECT 264.200 8.685 264.370 11.150 ;
        RECT 265.380 8.685 265.550 11.150 ;
        RECT 266.560 8.685 266.730 11.150 ;
        RECT 267.740 8.685 267.910 11.150 ;
        RECT 268.920 8.685 269.090 11.150 ;
        RECT 270.100 8.685 270.270 11.150 ;
        RECT 271.280 8.685 271.450 11.150 ;
        RECT 272.460 8.685 272.630 11.150 ;
        RECT 273.640 8.685 273.810 11.150 ;
        RECT 274.230 9.110 274.400 11.150 ;
        RECT 274.820 9.110 274.990 11.150 ;
        RECT 275.410 9.110 275.580 11.150 ;
        RECT 276.000 9.110 276.170 11.150 ;
        RECT 276.590 9.110 276.760 11.150 ;
        RECT 277.180 9.110 277.350 11.150 ;
        RECT 277.770 9.110 277.940 11.150 ;
        RECT 278.360 9.110 278.530 11.150 ;
        RECT 278.950 9.110 279.120 11.150 ;
        RECT 279.540 9.110 279.710 11.150 ;
        RECT 280.130 9.110 280.300 11.150 ;
        RECT 280.720 9.110 280.890 11.150 ;
        RECT 281.310 9.110 281.480 11.150 ;
        RECT 281.900 9.110 282.070 11.150 ;
        RECT 282.490 9.110 282.660 11.150 ;
        RECT 283.080 9.110 283.250 11.150 ;
        RECT 283.670 9.110 283.840 11.150 ;
        RECT 284.260 9.110 284.430 11.150 ;
        RECT 284.850 9.110 285.020 11.150 ;
        RECT 285.440 9.110 285.610 11.150 ;
        RECT 286.030 9.110 286.200 11.150 ;
        RECT 286.620 9.110 286.790 11.150 ;
        RECT 287.210 9.110 287.380 11.150 ;
        RECT 287.800 9.110 287.970 11.150 ;
        RECT 288.390 9.110 288.560 11.150 ;
        RECT 288.980 9.110 289.150 11.150 ;
        RECT 289.570 9.110 289.740 11.150 ;
        RECT 290.160 9.110 290.330 11.150 ;
        RECT 290.750 9.110 290.920 11.150 ;
        RECT 291.340 9.110 291.510 11.150 ;
        RECT 255.730 8.085 291.665 8.685 ;
        RECT 259.350 4.120 260.785 8.085 ;
        RECT 163.355 2.395 163.525 3.430 ;
        RECT 164.145 2.395 164.315 3.430 ;
        RECT 163.355 1.980 164.315 2.395 ;
        RECT 169.880 2.390 170.050 3.850 ;
        RECT 170.670 2.390 170.840 3.850 ;
        RECT 236.895 2.685 260.785 4.120 ;
        RECT 137.685 1.010 138.645 1.370 ;
        RECT 155.845 1.200 157.860 1.465 ;
        RECT 137.685 -0.955 137.855 1.010 ;
        RECT 138.475 -0.135 138.645 1.010 ;
        RECT 155.600 1.030 158.140 1.200 ;
        RECT 139.835 -0.910 140.005 0.915 ;
        RECT 141.415 -0.910 141.585 0.915 ;
        RECT 142.995 -0.910 143.165 0.915 ;
        RECT 144.575 -0.910 144.745 0.915 ;
        RECT 146.155 -0.910 146.325 0.915 ;
        RECT 147.530 -0.205 147.700 0.915 ;
        RECT 148.320 -0.205 148.490 0.915 ;
        RECT 147.530 -0.660 148.490 -0.205 ;
        RECT 147.945 -0.910 148.235 -0.660 ;
        RECT 151.650 -0.910 151.820 0.940 ;
        RECT 138.905 -0.955 151.820 -0.910 ;
        RECT 137.685 -1.125 151.820 -0.955 ;
        RECT 137.685 -5.775 138.630 -1.125 ;
        RECT 138.905 -1.200 151.820 -1.125 ;
        RECT 147.915 -1.455 151.820 -1.200 ;
        RECT 151.650 -1.870 151.820 -1.455 ;
        RECT 153.230 -1.870 153.400 0.940 ;
        RECT 154.810 -1.870 154.980 0.940 ;
        RECT 155.600 -1.100 155.770 1.030 ;
        RECT 156.390 -1.870 156.560 1.030 ;
        RECT 157.180 -1.100 157.350 1.030 ;
        RECT 157.970 -1.085 158.140 1.030 ;
        RECT 161.960 0.975 162.920 1.335 ;
        RECT 179.520 1.315 181.535 1.580 ;
        RECT 188.125 1.530 190.140 1.795 ;
        RECT 187.880 1.360 190.420 1.530 ;
        RECT 179.275 1.145 181.815 1.315 ;
        RECT 161.960 -0.990 162.130 0.975 ;
        RECT 162.750 -0.170 162.920 0.975 ;
        RECT 164.110 -0.945 164.280 0.880 ;
        RECT 165.690 -0.945 165.860 0.880 ;
        RECT 167.270 -0.945 167.440 0.880 ;
        RECT 168.850 -0.945 169.020 0.880 ;
        RECT 170.430 -0.945 170.600 0.880 ;
        RECT 171.805 -0.240 171.975 0.880 ;
        RECT 172.595 -0.240 172.765 0.880 ;
        RECT 171.805 -0.695 172.765 -0.240 ;
        RECT 172.220 -0.945 172.510 -0.695 ;
        RECT 163.180 -0.990 172.510 -0.945 ;
        RECT 161.960 -1.085 172.510 -0.990 ;
        RECT 157.970 -1.160 172.510 -1.085 ;
        RECT 157.970 -1.535 162.495 -1.160 ;
        RECT 163.180 -1.235 172.510 -1.160 ;
        RECT 172.100 -1.300 172.510 -1.235 ;
        RECT 175.325 -1.300 175.495 1.055 ;
        RECT 172.100 -1.470 175.495 -1.300 ;
        RECT 157.970 -1.870 158.140 -1.535 ;
        RECT 175.325 -1.755 175.495 -1.470 ;
        RECT 176.905 -1.755 177.075 1.055 ;
        RECT 178.485 -1.755 178.655 1.055 ;
        RECT 179.275 -0.985 179.445 1.145 ;
        RECT 180.065 -1.755 180.235 1.145 ;
        RECT 180.855 -0.985 181.025 1.145 ;
        RECT 181.645 -1.050 181.815 1.145 ;
        RECT 183.930 -1.050 184.100 1.270 ;
        RECT 181.645 -1.325 184.100 -1.050 ;
        RECT 181.645 -1.755 181.815 -1.325 ;
        RECT 183.930 -1.540 184.100 -1.325 ;
        RECT 185.510 -1.540 185.680 1.270 ;
        RECT 187.090 -1.540 187.260 1.270 ;
        RECT 187.880 -0.770 188.050 1.360 ;
        RECT 188.670 -1.540 188.840 1.360 ;
        RECT 189.460 -0.770 189.630 1.360 ;
        RECT 190.250 -1.540 190.420 1.360 ;
        RECT 151.525 -2.495 158.205 -1.870 ;
        RECT 175.200 -2.380 181.880 -1.755 ;
        RECT 183.805 -2.165 190.485 -1.540 ;
        RECT 236.895 -5.775 238.370 2.685 ;
        RECT 273.215 -3.085 290.625 -2.945 ;
        RECT 272.475 -3.405 290.625 -3.085 ;
        RECT 26.900 -6.880 27.070 -6.085 ;
        RECT 27.880 -6.880 28.050 -6.085 ;
        RECT 28.860 -6.880 29.030 -6.085 ;
        RECT 57.635 -6.195 75.045 -6.055 ;
        RECT 56.895 -6.515 75.045 -6.195 ;
        RECT 39.345 -8.980 39.515 -6.515 ;
        RECT 40.525 -8.980 40.695 -6.515 ;
        RECT 41.705 -8.980 41.875 -6.515 ;
        RECT 42.885 -8.980 43.055 -6.515 ;
        RECT 44.065 -8.980 44.235 -6.515 ;
        RECT 45.245 -8.980 45.415 -6.515 ;
        RECT 46.425 -8.980 46.595 -6.515 ;
        RECT 47.605 -8.980 47.775 -6.515 ;
        RECT 48.785 -8.980 48.955 -6.515 ;
        RECT 49.965 -8.980 50.135 -6.515 ;
        RECT 51.145 -8.980 51.315 -6.515 ;
        RECT 52.325 -8.980 52.495 -6.515 ;
        RECT 53.505 -8.980 53.675 -6.515 ;
        RECT 54.685 -8.980 54.855 -6.515 ;
        RECT 55.865 -8.980 56.035 -6.515 ;
        RECT 57.045 -8.980 57.215 -6.515 ;
        RECT 57.635 -8.555 57.805 -6.515 ;
        RECT 58.225 -8.555 58.395 -6.515 ;
        RECT 58.815 -8.555 58.985 -6.515 ;
        RECT 59.405 -8.555 59.575 -6.515 ;
        RECT 59.995 -8.555 60.165 -6.515 ;
        RECT 60.585 -8.555 60.755 -6.515 ;
        RECT 61.175 -8.555 61.345 -6.515 ;
        RECT 61.765 -8.555 61.935 -6.515 ;
        RECT 62.355 -8.555 62.525 -6.515 ;
        RECT 62.945 -8.555 63.115 -6.515 ;
        RECT 63.535 -8.555 63.705 -6.515 ;
        RECT 64.125 -8.555 64.295 -6.515 ;
        RECT 64.715 -8.555 64.885 -6.515 ;
        RECT 65.305 -8.555 65.475 -6.515 ;
        RECT 65.895 -8.555 66.065 -6.515 ;
        RECT 66.485 -8.555 66.655 -6.515 ;
        RECT 67.075 -8.555 67.245 -6.515 ;
        RECT 67.665 -8.555 67.835 -6.515 ;
        RECT 68.255 -8.555 68.425 -6.515 ;
        RECT 68.845 -8.555 69.015 -6.515 ;
        RECT 69.435 -8.555 69.605 -6.515 ;
        RECT 70.025 -8.555 70.195 -6.515 ;
        RECT 70.615 -8.555 70.785 -6.515 ;
        RECT 71.205 -8.555 71.375 -6.515 ;
        RECT 71.795 -8.555 71.965 -6.515 ;
        RECT 72.385 -8.555 72.555 -6.515 ;
        RECT 72.975 -8.555 73.145 -6.515 ;
        RECT 73.565 -8.555 73.735 -6.515 ;
        RECT 74.155 -8.555 74.325 -6.515 ;
        RECT 74.745 -8.555 74.915 -6.515 ;
        RECT 127.865 -7.250 238.370 -5.775 ;
        RECT 254.925 -5.870 255.095 -3.405 ;
        RECT 256.105 -5.870 256.275 -3.405 ;
        RECT 257.285 -5.870 257.455 -3.405 ;
        RECT 258.465 -5.870 258.635 -3.405 ;
        RECT 259.645 -5.870 259.815 -3.405 ;
        RECT 260.825 -5.870 260.995 -3.405 ;
        RECT 262.005 -5.870 262.175 -3.405 ;
        RECT 263.185 -5.870 263.355 -3.405 ;
        RECT 264.365 -5.870 264.535 -3.405 ;
        RECT 265.545 -5.870 265.715 -3.405 ;
        RECT 266.725 -5.870 266.895 -3.405 ;
        RECT 267.905 -5.870 268.075 -3.405 ;
        RECT 269.085 -5.870 269.255 -3.405 ;
        RECT 270.265 -5.870 270.435 -3.405 ;
        RECT 271.445 -5.870 271.615 -3.405 ;
        RECT 272.625 -5.870 272.795 -3.405 ;
        RECT 273.215 -5.445 273.385 -3.405 ;
        RECT 273.805 -5.445 273.975 -3.405 ;
        RECT 274.395 -5.445 274.565 -3.405 ;
        RECT 274.985 -5.445 275.155 -3.405 ;
        RECT 275.575 -5.445 275.745 -3.405 ;
        RECT 276.165 -5.445 276.335 -3.405 ;
        RECT 276.755 -5.445 276.925 -3.405 ;
        RECT 277.345 -5.445 277.515 -3.405 ;
        RECT 277.935 -5.445 278.105 -3.405 ;
        RECT 278.525 -5.445 278.695 -3.405 ;
        RECT 279.115 -5.445 279.285 -3.405 ;
        RECT 279.705 -5.445 279.875 -3.405 ;
        RECT 280.295 -5.445 280.465 -3.405 ;
        RECT 280.885 -5.445 281.055 -3.405 ;
        RECT 281.475 -5.445 281.645 -3.405 ;
        RECT 282.065 -5.445 282.235 -3.405 ;
        RECT 282.655 -5.445 282.825 -3.405 ;
        RECT 283.245 -5.445 283.415 -3.405 ;
        RECT 283.835 -5.445 284.005 -3.405 ;
        RECT 284.425 -5.445 284.595 -3.405 ;
        RECT 285.015 -5.445 285.185 -3.405 ;
        RECT 285.605 -5.445 285.775 -3.405 ;
        RECT 286.195 -5.445 286.365 -3.405 ;
        RECT 286.785 -5.445 286.955 -3.405 ;
        RECT 287.375 -5.445 287.545 -3.405 ;
        RECT 287.965 -5.445 288.135 -3.405 ;
        RECT 288.555 -5.445 288.725 -3.405 ;
        RECT 289.145 -5.445 289.315 -3.405 ;
        RECT 289.735 -5.445 289.905 -3.405 ;
        RECT 290.325 -5.445 290.495 -3.405 ;
        RECT 254.715 -6.470 290.650 -5.870 ;
        RECT 39.135 -9.580 75.070 -8.980 ;
        RECT 41.680 -9.830 42.785 -9.580 ;
        RECT 46.370 -9.830 47.735 -9.580 ;
        RECT 51.275 -9.830 52.640 -9.580 ;
        RECT 57.285 -9.830 58.650 -9.580 ;
        RECT 62.060 -9.830 63.425 -9.580 ;
        RECT 66.030 -9.830 67.395 -9.580 ;
        RECT 69.655 -9.830 71.020 -9.580 ;
        RECT 131.405 -9.830 133.190 -7.250 ;
        RECT 40.840 -11.615 133.190 -9.830 ;
        RECT 234.320 -8.685 236.845 -7.250 ;
        RECT 262.315 -8.685 264.840 -6.470 ;
        RECT 234.320 -11.210 264.840 -8.685 ;
        RECT 234.320 -12.575 236.845 -11.210 ;
        RECT 311.965 -16.865 312.135 -16.070 ;
        RECT 312.945 -16.865 313.115 -16.070 ;
        RECT 313.925 -16.865 314.095 -16.070 ;
        RECT 316.215 -16.865 316.385 -16.070 ;
        RECT 317.195 -16.865 317.365 -16.070 ;
        RECT 318.175 -16.865 318.345 -16.070 ;
        RECT 311.920 -17.205 318.840 -16.865 ;
        RECT 316.170 -17.890 318.840 -17.205 ;
        RECT 273.215 -18.320 290.625 -18.180 ;
        RECT 272.475 -18.640 290.625 -18.320 ;
        RECT 254.925 -21.105 255.095 -18.640 ;
        RECT 256.105 -21.105 256.275 -18.640 ;
        RECT 257.285 -21.105 257.455 -18.640 ;
        RECT 258.465 -21.105 258.635 -18.640 ;
        RECT 259.645 -21.105 259.815 -18.640 ;
        RECT 260.825 -21.105 260.995 -18.640 ;
        RECT 262.005 -21.105 262.175 -18.640 ;
        RECT 263.185 -21.105 263.355 -18.640 ;
        RECT 264.365 -21.105 264.535 -18.640 ;
        RECT 265.545 -21.105 265.715 -18.640 ;
        RECT 266.725 -21.105 266.895 -18.640 ;
        RECT 267.905 -21.105 268.075 -18.640 ;
        RECT 269.085 -21.105 269.255 -18.640 ;
        RECT 270.265 -21.105 270.435 -18.640 ;
        RECT 271.445 -21.105 271.615 -18.640 ;
        RECT 272.625 -21.105 272.795 -18.640 ;
        RECT 273.215 -20.680 273.385 -18.640 ;
        RECT 273.805 -20.680 273.975 -18.640 ;
        RECT 274.395 -20.680 274.565 -18.640 ;
        RECT 274.985 -20.680 275.155 -18.640 ;
        RECT 275.575 -20.680 275.745 -18.640 ;
        RECT 276.165 -20.680 276.335 -18.640 ;
        RECT 276.755 -20.680 276.925 -18.640 ;
        RECT 277.345 -20.680 277.515 -18.640 ;
        RECT 277.935 -20.680 278.105 -18.640 ;
        RECT 278.525 -20.680 278.695 -18.640 ;
        RECT 279.115 -20.680 279.285 -18.640 ;
        RECT 279.705 -20.680 279.875 -18.640 ;
        RECT 280.295 -20.680 280.465 -18.640 ;
        RECT 280.885 -20.680 281.055 -18.640 ;
        RECT 281.475 -20.680 281.645 -18.640 ;
        RECT 282.065 -20.680 282.235 -18.640 ;
        RECT 282.655 -20.680 282.825 -18.640 ;
        RECT 283.245 -20.680 283.415 -18.640 ;
        RECT 283.835 -20.680 284.005 -18.640 ;
        RECT 284.425 -20.680 284.595 -18.640 ;
        RECT 285.015 -20.680 285.185 -18.640 ;
        RECT 285.605 -20.680 285.775 -18.640 ;
        RECT 286.195 -20.680 286.365 -18.640 ;
        RECT 286.785 -20.680 286.955 -18.640 ;
        RECT 287.375 -20.680 287.545 -18.640 ;
        RECT 287.965 -20.680 288.135 -18.640 ;
        RECT 288.555 -20.680 288.725 -18.640 ;
        RECT 289.145 -20.680 289.315 -18.640 ;
        RECT 289.735 -20.680 289.905 -18.640 ;
        RECT 290.325 -20.680 290.495 -18.640 ;
        RECT 316.215 -18.685 316.385 -17.890 ;
        RECT 317.195 -18.685 317.365 -17.890 ;
        RECT 318.175 -18.685 318.345 -17.890 ;
        RECT 254.715 -21.705 290.650 -21.105 ;
        RECT 233.890 -23.490 236.990 -23.350 ;
        RECT 262.855 -23.490 265.740 -21.705 ;
        RECT 233.890 -26.375 464.795 -23.490 ;
        RECT 233.890 -26.520 237.060 -26.375 ;
        RECT 350.385 -38.335 464.795 -26.375 ;
        RECT 350.385 -39.015 365.230 -38.335 ;
        RECT 407.755 -39.015 422.600 -38.335 ;
        RECT 451.645 -90.205 458.510 -87.520 ;
        RECT 442.140 -92.895 458.510 -90.205 ;
        RECT 451.645 -94.385 458.510 -92.895 ;
        RECT 453.020 -173.160 461.105 -169.440 ;
        RECT 443.815 -175.850 461.105 -173.160 ;
        RECT 453.020 -177.070 461.105 -175.850 ;
        RECT 456.545 -263.715 462.960 -261.010 ;
        RECT 447.000 -266.405 462.960 -263.715 ;
        RECT 456.545 -267.730 462.960 -266.405 ;
      LAYER met1 ;
        RECT -64.360 601.795 -52.250 602.360 ;
        RECT -64.360 584.020 -63.795 601.795 ;
        RECT -52.815 598.820 -52.250 601.795 ;
        RECT -63.255 598.270 -61.755 598.500 ;
        RECT -53.490 597.865 -52.990 598.095 ;
        RECT -63.255 597.060 -61.755 597.290 ;
        RECT -53.490 596.885 -52.990 597.115 ;
        RECT -63.255 596.080 -61.755 596.310 ;
        RECT -51.955 593.840 -50.455 594.070 ;
        RECT -45.545 593.485 -44.045 593.715 ;
        RECT -59.290 592.870 -58.790 593.100 ;
        RECT -59.290 591.890 -58.790 592.120 ;
        RECT -45.545 591.855 -43.045 592.085 ;
        RECT -45.545 591.205 -43.045 591.435 ;
        RECT -52.345 589.955 -51.345 590.185 ;
        RECT -61.825 588.845 -60.325 589.075 ;
        RECT -52.345 588.975 -51.345 589.205 ;
        RECT -45.545 587.250 -44.045 587.480 ;
        RECT -64.360 583.455 -52.095 584.020 ;
        RECT -64.360 580.655 -63.640 583.455 ;
        RECT -64.205 580.635 -63.640 580.655 ;
        RECT -52.660 582.190 -52.095 583.455 ;
        RECT -46.940 583.495 -34.830 584.060 ;
        RECT -46.940 582.190 -46.375 583.495 ;
        RECT -52.660 581.625 -46.370 582.190 ;
        RECT -52.660 580.480 -52.095 581.625 ;
        RECT -46.940 580.675 -46.375 581.625 ;
        RECT -35.395 580.520 -34.830 583.495 ;
        RECT -63.100 579.930 -61.600 580.160 ;
        RECT -45.835 579.970 -44.335 580.200 ;
        RECT -53.335 579.525 -52.835 579.755 ;
        RECT -36.070 579.565 -35.570 579.795 ;
        RECT -63.100 578.720 -61.600 578.950 ;
        RECT -53.335 578.545 -52.835 578.775 ;
        RECT -45.835 578.760 -44.335 578.990 ;
        RECT -36.070 578.585 -35.570 578.815 ;
        RECT -63.100 577.740 -61.600 577.970 ;
        RECT -45.835 577.780 -44.335 578.010 ;
        RECT -51.800 575.500 -50.300 575.730 ;
        RECT -34.535 575.540 -33.035 575.770 ;
        RECT -59.135 574.530 -58.635 574.760 ;
        RECT -41.870 574.570 -41.370 574.800 ;
        RECT -59.135 573.550 -58.635 573.780 ;
        RECT -41.870 573.590 -41.370 573.820 ;
        RECT -52.190 571.615 -51.190 571.845 ;
        RECT -34.925 571.655 -33.925 571.885 ;
        RECT -61.670 570.505 -60.170 570.735 ;
        RECT -52.190 570.635 -51.190 570.865 ;
        RECT -44.405 570.545 -42.905 570.775 ;
        RECT -34.925 570.675 -33.925 570.905 ;
        RECT -64.550 554.975 -52.440 555.540 ;
        RECT -64.550 537.200 -63.985 554.975 ;
        RECT -53.005 552.000 -52.440 554.975 ;
        RECT -63.445 551.450 -61.945 551.680 ;
        RECT -53.680 551.045 -53.180 551.275 ;
        RECT -63.445 550.240 -61.945 550.470 ;
        RECT -53.680 550.065 -53.180 550.295 ;
        RECT -63.445 549.260 -61.945 549.490 ;
        RECT -52.145 547.020 -50.645 547.250 ;
        RECT -45.735 546.665 -44.235 546.895 ;
        RECT -59.480 546.050 -58.980 546.280 ;
        RECT -59.480 545.070 -58.980 545.300 ;
        RECT -45.735 545.035 -43.235 545.265 ;
        RECT -45.735 544.385 -43.235 544.615 ;
        RECT -52.535 543.135 -51.535 543.365 ;
        RECT -62.015 542.025 -60.515 542.255 ;
        RECT -52.535 542.155 -51.535 542.385 ;
        RECT -45.735 540.430 -44.235 540.660 ;
        RECT -64.550 536.635 -52.285 537.200 ;
        RECT -64.550 533.835 -63.830 536.635 ;
        RECT -64.395 533.815 -63.830 533.835 ;
        RECT -52.850 535.370 -52.285 536.635 ;
        RECT -47.130 536.675 -35.020 537.240 ;
        RECT -47.130 535.370 -46.565 536.675 ;
        RECT -52.850 534.805 -46.560 535.370 ;
        RECT -52.850 533.660 -52.285 534.805 ;
        RECT -47.130 533.855 -46.565 534.805 ;
        RECT -35.585 533.700 -35.020 536.675 ;
        RECT -63.290 533.110 -61.790 533.340 ;
        RECT -46.025 533.150 -44.525 533.380 ;
        RECT -53.525 532.705 -53.025 532.935 ;
        RECT -36.260 532.745 -35.760 532.975 ;
        RECT -63.290 531.900 -61.790 532.130 ;
        RECT -53.525 531.725 -53.025 531.955 ;
        RECT -46.025 531.940 -44.525 532.170 ;
        RECT -36.260 531.765 -35.760 531.995 ;
        RECT -63.290 530.920 -61.790 531.150 ;
        RECT -46.025 530.960 -44.525 531.190 ;
        RECT -51.990 528.680 -50.490 528.910 ;
        RECT -34.725 528.720 -33.225 528.950 ;
        RECT -59.325 527.710 -58.825 527.940 ;
        RECT -42.060 527.750 -41.560 527.980 ;
        RECT -59.325 526.730 -58.825 526.960 ;
        RECT -42.060 526.770 -41.560 527.000 ;
        RECT -52.380 524.795 -51.380 525.025 ;
        RECT -35.115 524.835 -34.115 525.065 ;
        RECT -61.860 523.685 -60.360 523.915 ;
        RECT -52.380 523.815 -51.380 524.045 ;
        RECT -44.595 523.725 -43.095 523.955 ;
        RECT -35.115 523.855 -34.115 524.085 ;
        RECT -64.635 509.210 -52.525 509.775 ;
        RECT -64.635 491.435 -64.070 509.210 ;
        RECT -53.090 506.235 -52.525 509.210 ;
        RECT -63.530 505.685 -62.030 505.915 ;
        RECT -53.765 505.280 -53.265 505.510 ;
        RECT -63.530 504.475 -62.030 504.705 ;
        RECT -53.765 504.300 -53.265 504.530 ;
        RECT -63.530 503.495 -62.030 503.725 ;
        RECT -52.230 501.255 -50.730 501.485 ;
        RECT -45.820 500.900 -44.320 501.130 ;
        RECT -59.565 500.285 -59.065 500.515 ;
        RECT -59.565 499.305 -59.065 499.535 ;
        RECT -45.820 499.270 -43.320 499.500 ;
        RECT -45.820 498.620 -43.320 498.850 ;
        RECT -52.620 497.370 -51.620 497.600 ;
        RECT -62.100 496.260 -60.600 496.490 ;
        RECT -52.620 496.390 -51.620 496.620 ;
        RECT -45.820 494.665 -44.320 494.895 ;
        RECT -64.635 490.870 -52.370 491.435 ;
        RECT -64.635 488.070 -63.915 490.870 ;
        RECT -64.480 488.050 -63.915 488.070 ;
        RECT -52.935 489.605 -52.370 490.870 ;
        RECT -47.215 490.910 -35.105 491.475 ;
        RECT -47.215 489.605 -46.650 490.910 ;
        RECT -52.935 489.040 -46.645 489.605 ;
        RECT -52.935 487.895 -52.370 489.040 ;
        RECT -47.215 488.090 -46.650 489.040 ;
        RECT -35.670 487.935 -35.105 490.910 ;
        RECT -63.375 487.345 -61.875 487.575 ;
        RECT -46.110 487.385 -44.610 487.615 ;
        RECT -53.610 486.940 -53.110 487.170 ;
        RECT -36.345 486.980 -35.845 487.210 ;
        RECT -63.375 486.135 -61.875 486.365 ;
        RECT -53.610 485.960 -53.110 486.190 ;
        RECT -46.110 486.175 -44.610 486.405 ;
        RECT -36.345 486.000 -35.845 486.230 ;
        RECT -63.375 485.155 -61.875 485.385 ;
        RECT -46.110 485.195 -44.610 485.425 ;
        RECT -52.075 482.915 -50.575 483.145 ;
        RECT -34.810 482.955 -33.310 483.185 ;
        RECT -59.410 481.945 -58.910 482.175 ;
        RECT -42.145 481.985 -41.645 482.215 ;
        RECT -59.410 480.965 -58.910 481.195 ;
        RECT -42.145 481.005 -41.645 481.235 ;
        RECT -52.465 479.030 -51.465 479.260 ;
        RECT -35.200 479.070 -34.200 479.300 ;
        RECT -61.945 477.920 -60.445 478.150 ;
        RECT -52.465 478.050 -51.465 478.280 ;
        RECT -44.680 477.960 -43.180 478.190 ;
        RECT -35.200 478.090 -34.200 478.320 ;
        RECT -64.965 465.440 -52.855 466.005 ;
        RECT -64.965 447.665 -64.400 465.440 ;
        RECT -53.420 462.465 -52.855 465.440 ;
        RECT -63.860 461.915 -62.360 462.145 ;
        RECT -54.095 461.510 -53.595 461.740 ;
        RECT -63.860 460.705 -62.360 460.935 ;
        RECT -54.095 460.530 -53.595 460.760 ;
        RECT -63.860 459.725 -62.360 459.955 ;
        RECT -52.560 457.485 -51.060 457.715 ;
        RECT -46.150 457.130 -44.650 457.360 ;
        RECT -59.895 456.515 -59.395 456.745 ;
        RECT -59.895 455.535 -59.395 455.765 ;
        RECT -46.150 455.500 -43.650 455.730 ;
        RECT -46.150 454.850 -43.650 455.080 ;
        RECT -52.950 453.600 -51.950 453.830 ;
        RECT -62.430 452.490 -60.930 452.720 ;
        RECT -52.950 452.620 -51.950 452.850 ;
        RECT -46.150 450.895 -44.650 451.125 ;
        RECT -64.965 447.100 -52.700 447.665 ;
        RECT -64.965 444.300 -64.245 447.100 ;
        RECT -64.810 444.280 -64.245 444.300 ;
        RECT -53.265 445.835 -52.700 447.100 ;
        RECT -47.545 447.140 -35.435 447.705 ;
        RECT -47.545 445.835 -46.980 447.140 ;
        RECT -53.265 445.270 -46.975 445.835 ;
        RECT -53.265 444.125 -52.700 445.270 ;
        RECT -47.545 444.320 -46.980 445.270 ;
        RECT -36.000 444.165 -35.435 447.140 ;
        RECT -63.705 443.575 -62.205 443.805 ;
        RECT -46.440 443.615 -44.940 443.845 ;
        RECT -53.940 443.170 -53.440 443.400 ;
        RECT -36.675 443.210 -36.175 443.440 ;
        RECT -63.705 442.365 -62.205 442.595 ;
        RECT -53.940 442.190 -53.440 442.420 ;
        RECT -46.440 442.405 -44.940 442.635 ;
        RECT -36.675 442.230 -36.175 442.460 ;
        RECT -63.705 441.385 -62.205 441.615 ;
        RECT -46.440 441.425 -44.940 441.655 ;
        RECT -52.405 439.145 -50.905 439.375 ;
        RECT -35.140 439.185 -33.640 439.415 ;
        RECT -59.740 438.175 -59.240 438.405 ;
        RECT -42.475 438.215 -41.975 438.445 ;
        RECT -59.740 437.195 -59.240 437.425 ;
        RECT -42.475 437.235 -41.975 437.465 ;
        RECT -52.795 435.260 -51.795 435.490 ;
        RECT -35.530 435.300 -34.530 435.530 ;
        RECT -62.275 434.150 -60.775 434.380 ;
        RECT -52.795 434.280 -51.795 434.510 ;
        RECT -45.010 434.190 -43.510 434.420 ;
        RECT -35.530 434.320 -34.530 434.550 ;
        RECT -65.135 419.450 -53.025 420.015 ;
        RECT -65.135 401.675 -64.570 419.450 ;
        RECT -53.590 416.475 -53.025 419.450 ;
        RECT -64.030 415.925 -62.530 416.155 ;
        RECT -54.265 415.520 -53.765 415.750 ;
        RECT -64.030 414.715 -62.530 414.945 ;
        RECT -54.265 414.540 -53.765 414.770 ;
        RECT -64.030 413.735 -62.530 413.965 ;
        RECT -52.730 411.495 -51.230 411.725 ;
        RECT -46.320 411.140 -44.820 411.370 ;
        RECT -60.065 410.525 -59.565 410.755 ;
        RECT -60.065 409.545 -59.565 409.775 ;
        RECT -46.320 409.510 -43.820 409.740 ;
        RECT -46.320 408.860 -43.820 409.090 ;
        RECT -53.120 407.610 -52.120 407.840 ;
        RECT -62.600 406.500 -61.100 406.730 ;
        RECT -53.120 406.630 -52.120 406.860 ;
        RECT -46.320 404.905 -44.820 405.135 ;
        RECT -65.135 401.110 -52.870 401.675 ;
        RECT -65.135 398.310 -64.415 401.110 ;
        RECT -64.980 398.290 -64.415 398.310 ;
        RECT -53.435 399.845 -52.870 401.110 ;
        RECT -47.715 401.150 -35.605 401.715 ;
        RECT -47.715 399.845 -47.150 401.150 ;
        RECT -53.435 399.280 -47.145 399.845 ;
        RECT -53.435 398.135 -52.870 399.280 ;
        RECT -47.715 398.330 -47.150 399.280 ;
        RECT -36.170 398.175 -35.605 401.150 ;
        RECT -63.875 397.585 -62.375 397.815 ;
        RECT -46.610 397.625 -45.110 397.855 ;
        RECT -54.110 397.180 -53.610 397.410 ;
        RECT -36.845 397.220 -36.345 397.450 ;
        RECT -63.875 396.375 -62.375 396.605 ;
        RECT -54.110 396.200 -53.610 396.430 ;
        RECT -46.610 396.415 -45.110 396.645 ;
        RECT -36.845 396.240 -36.345 396.470 ;
        RECT -63.875 395.395 -62.375 395.625 ;
        RECT -46.610 395.435 -45.110 395.665 ;
        RECT -52.575 393.155 -51.075 393.385 ;
        RECT -35.310 393.195 -33.810 393.425 ;
        RECT -59.910 392.185 -59.410 392.415 ;
        RECT -42.645 392.225 -42.145 392.455 ;
        RECT -59.910 391.205 -59.410 391.435 ;
        RECT -42.645 391.245 -42.145 391.475 ;
        RECT -52.965 389.270 -51.965 389.500 ;
        RECT -35.700 389.310 -34.700 389.540 ;
        RECT -62.445 388.160 -60.945 388.390 ;
        RECT -52.965 388.290 -51.965 388.520 ;
        RECT -45.180 388.200 -43.680 388.430 ;
        RECT -35.700 388.330 -34.700 388.560 ;
        RECT -64.940 375.135 -52.830 375.700 ;
        RECT -64.940 357.360 -64.375 375.135 ;
        RECT -53.395 372.160 -52.830 375.135 ;
        RECT -63.835 371.610 -62.335 371.840 ;
        RECT -54.070 371.205 -53.570 371.435 ;
        RECT -63.835 370.400 -62.335 370.630 ;
        RECT -54.070 370.225 -53.570 370.455 ;
        RECT -63.835 369.420 -62.335 369.650 ;
        RECT -52.535 367.180 -51.035 367.410 ;
        RECT -46.125 366.825 -44.625 367.055 ;
        RECT -59.870 366.210 -59.370 366.440 ;
        RECT -59.870 365.230 -59.370 365.460 ;
        RECT -46.125 365.195 -43.625 365.425 ;
        RECT -46.125 364.545 -43.625 364.775 ;
        RECT -52.925 363.295 -51.925 363.525 ;
        RECT -62.405 362.185 -60.905 362.415 ;
        RECT -52.925 362.315 -51.925 362.545 ;
        RECT -46.125 360.590 -44.625 360.820 ;
        RECT -64.940 356.795 -52.675 357.360 ;
        RECT -64.940 353.995 -64.220 356.795 ;
        RECT -64.785 353.975 -64.220 353.995 ;
        RECT -53.240 355.530 -52.675 356.795 ;
        RECT -47.520 356.835 -35.410 357.400 ;
        RECT -47.520 355.530 -46.955 356.835 ;
        RECT -53.240 354.965 -46.950 355.530 ;
        RECT -53.240 353.820 -52.675 354.965 ;
        RECT -47.520 354.015 -46.955 354.965 ;
        RECT -35.975 353.860 -35.410 356.835 ;
        RECT -63.680 353.270 -62.180 353.500 ;
        RECT -46.415 353.310 -44.915 353.540 ;
        RECT -53.915 352.865 -53.415 353.095 ;
        RECT -36.650 352.905 -36.150 353.135 ;
        RECT -63.680 352.060 -62.180 352.290 ;
        RECT -53.915 351.885 -53.415 352.115 ;
        RECT -46.415 352.100 -44.915 352.330 ;
        RECT -36.650 351.925 -36.150 352.155 ;
        RECT -63.680 351.080 -62.180 351.310 ;
        RECT -46.415 351.120 -44.915 351.350 ;
        RECT -52.380 348.840 -50.880 349.070 ;
        RECT -35.115 348.880 -33.615 349.110 ;
        RECT -59.715 347.870 -59.215 348.100 ;
        RECT -42.450 347.910 -41.950 348.140 ;
        RECT -59.715 346.890 -59.215 347.120 ;
        RECT -42.450 346.930 -41.950 347.160 ;
        RECT -52.770 344.955 -51.770 345.185 ;
        RECT -35.505 344.995 -34.505 345.225 ;
        RECT -62.250 343.845 -60.750 344.075 ;
        RECT -52.770 343.975 -51.770 344.205 ;
        RECT -44.985 343.885 -43.485 344.115 ;
        RECT -35.505 344.015 -34.505 344.245 ;
        RECT -64.885 332.935 -52.775 333.500 ;
        RECT -64.885 315.160 -64.320 332.935 ;
        RECT -53.340 329.960 -52.775 332.935 ;
        RECT -63.780 329.410 -62.280 329.640 ;
        RECT -54.015 329.005 -53.515 329.235 ;
        RECT -63.780 328.200 -62.280 328.430 ;
        RECT -54.015 328.025 -53.515 328.255 ;
        RECT -63.780 327.220 -62.280 327.450 ;
        RECT -52.480 324.980 -50.980 325.210 ;
        RECT -46.070 324.625 -44.570 324.855 ;
        RECT -59.815 324.010 -59.315 324.240 ;
        RECT -59.815 323.030 -59.315 323.260 ;
        RECT -46.070 322.995 -43.570 323.225 ;
        RECT -46.070 322.345 -43.570 322.575 ;
        RECT -52.870 321.095 -51.870 321.325 ;
        RECT -62.350 319.985 -60.850 320.215 ;
        RECT -52.870 320.115 -51.870 320.345 ;
        RECT -46.070 318.390 -44.570 318.620 ;
        RECT -64.885 314.595 -52.620 315.160 ;
        RECT -64.885 311.795 -64.165 314.595 ;
        RECT -64.730 311.775 -64.165 311.795 ;
        RECT -53.185 313.330 -52.620 314.595 ;
        RECT -47.465 314.635 -35.355 315.200 ;
        RECT -47.465 313.330 -46.900 314.635 ;
        RECT -53.185 312.765 -46.895 313.330 ;
        RECT -53.185 311.620 -52.620 312.765 ;
        RECT -47.465 311.815 -46.900 312.765 ;
        RECT -35.920 311.660 -35.355 314.635 ;
        RECT -63.625 311.070 -62.125 311.300 ;
        RECT -46.360 311.110 -44.860 311.340 ;
        RECT -53.860 310.665 -53.360 310.895 ;
        RECT -36.595 310.705 -36.095 310.935 ;
        RECT -63.625 309.860 -62.125 310.090 ;
        RECT -53.860 309.685 -53.360 309.915 ;
        RECT -46.360 309.900 -44.860 310.130 ;
        RECT -36.595 309.725 -36.095 309.955 ;
        RECT -63.625 308.880 -62.125 309.110 ;
        RECT -46.360 308.920 -44.860 309.150 ;
        RECT -52.325 306.640 -50.825 306.870 ;
        RECT -35.060 306.680 -33.560 306.910 ;
        RECT -59.660 305.670 -59.160 305.900 ;
        RECT -42.395 305.710 -41.895 305.940 ;
        RECT -59.660 304.690 -59.160 304.920 ;
        RECT -42.395 304.730 -41.895 304.960 ;
        RECT -52.715 302.755 -51.715 302.985 ;
        RECT -35.450 302.795 -34.450 303.025 ;
        RECT -62.195 301.645 -60.695 301.875 ;
        RECT -52.715 301.775 -51.715 302.005 ;
        RECT -44.930 301.685 -43.430 301.915 ;
        RECT -35.450 301.815 -34.450 302.045 ;
        RECT -40.265 289.110 -39.765 289.340 ;
        RECT -51.940 288.410 -48.440 288.640 ;
        RECT -43.555 288.620 -43.055 288.850 ;
        RECT -42.770 288.095 -42.470 288.215 ;
        RECT -41.380 288.095 -41.080 288.170 ;
        RECT -40.265 288.130 -39.765 288.360 ;
        RECT -43.555 287.640 -43.055 287.870 ;
        RECT -42.770 287.620 -41.080 288.095 ;
        RECT -42.770 287.555 -42.470 287.620 ;
        RECT -41.380 287.485 -41.080 287.620 ;
        RECT -40.265 287.150 -39.765 287.380 ;
        RECT -43.555 286.660 -43.055 286.890 ;
        RECT -51.940 286.410 -48.440 286.640 ;
        RECT -40.265 284.925 -39.765 285.155 ;
        RECT -40.265 283.945 -39.765 284.175 ;
        RECT -51.940 283.410 -48.440 283.640 ;
        RECT -40.265 282.965 -39.765 283.195 ;
        RECT -51.940 281.410 -48.440 281.640 ;
        RECT -43.555 279.905 -43.055 280.135 ;
        RECT -43.555 278.925 -43.055 279.155 ;
        RECT -51.940 278.410 -48.440 278.640 ;
        RECT -43.555 277.945 -43.055 278.175 ;
        RECT -51.940 276.410 -48.440 276.640 ;
        RECT -40.265 275.610 -39.765 275.840 ;
        RECT -43.555 275.120 -43.055 275.350 ;
        RECT -42.750 275.130 -42.450 275.220 ;
        RECT -41.410 275.130 -41.110 275.185 ;
        RECT -42.750 274.655 -41.110 275.130 ;
        RECT -42.750 274.535 -42.450 274.655 ;
        RECT -41.410 274.500 -41.110 274.655 ;
        RECT -40.265 274.630 -39.765 274.860 ;
        RECT -54.820 273.970 -54.320 274.200 ;
        RECT -43.555 274.140 -43.055 274.370 ;
        RECT -40.265 273.650 -39.765 273.880 ;
        RECT -54.820 272.990 -54.320 273.220 ;
        RECT -43.555 273.160 -43.055 273.390 ;
        RECT -52.485 272.260 -51.485 272.490 ;
        RECT -54.820 272.010 -54.320 272.240 ;
        RECT -40.265 271.425 -39.765 271.655 ;
        RECT -40.265 270.445 -39.765 270.675 ;
        RECT -40.265 269.465 -39.765 269.695 ;
        RECT -53.215 268.365 -52.215 268.595 ;
        RECT -43.555 266.405 -43.055 266.635 ;
        RECT -43.555 265.425 -43.055 265.655 ;
        RECT -43.555 264.445 -43.055 264.675 ;
        RECT -53.720 263.205 -52.220 263.435 ;
        RECT -43.555 261.995 -43.055 262.225 ;
        RECT -42.755 261.910 -42.455 262.085 ;
        RECT -41.410 261.910 -41.110 261.995 ;
        RECT -42.755 261.435 -41.110 261.910 ;
        RECT -42.755 261.400 -42.455 261.435 ;
        RECT -41.410 261.335 -41.110 261.435 ;
        RECT -43.555 261.015 -43.055 261.245 ;
        RECT -43.555 260.035 -43.055 260.265 ;
        RECT -53.125 259.605 -52.125 259.835 ;
        RECT -53.125 258.625 -52.125 258.855 ;
        RECT -53.125 254.875 -52.125 255.105 ;
        RECT -40.035 254.900 -39.035 255.130 ;
        RECT -53.125 253.895 -52.125 254.125 ;
        RECT -40.035 253.920 -39.035 254.150 ;
        RECT -66.335 248.470 -65.835 248.700 ;
        RECT -63.045 247.980 -62.545 248.210 ;
        RECT -66.335 247.490 -65.835 247.720 ;
        RECT -65.020 247.455 -64.720 247.530 ;
        RECT -63.630 247.455 -63.330 247.575 ;
        RECT -65.020 246.980 -63.330 247.455 ;
        RECT -63.045 247.000 -62.545 247.230 ;
        RECT -65.020 246.845 -64.720 246.980 ;
        RECT -63.630 246.915 -63.330 246.980 ;
        RECT -66.335 246.510 -65.835 246.740 ;
        RECT -63.045 246.020 -62.545 246.250 ;
        RECT -66.335 244.285 -65.835 244.515 ;
        RECT -66.335 243.305 -65.835 243.535 ;
        RECT -66.335 242.325 -65.835 242.555 ;
        RECT -63.045 239.265 -62.545 239.495 ;
        RECT -63.045 238.285 -62.545 238.515 ;
        RECT -63.045 237.305 -62.545 237.535 ;
        RECT -66.335 234.970 -65.835 235.200 ;
        RECT -64.990 234.490 -64.690 234.545 ;
        RECT -63.650 234.490 -63.350 234.580 ;
        RECT -66.335 233.990 -65.835 234.220 ;
        RECT -64.990 234.015 -63.350 234.490 ;
        RECT -63.045 234.480 -62.545 234.710 ;
        RECT -64.990 233.860 -64.690 234.015 ;
        RECT -63.650 233.895 -63.350 234.015 ;
        RECT -63.045 233.500 -62.545 233.730 ;
        RECT -66.335 233.010 -65.835 233.240 ;
        RECT -63.045 232.520 -62.545 232.750 ;
        RECT -66.335 230.785 -65.835 231.015 ;
        RECT -66.335 229.805 -65.835 230.035 ;
        RECT -66.335 228.825 -65.835 229.055 ;
        RECT -63.045 225.765 -62.545 225.995 ;
        RECT -63.045 224.785 -62.545 225.015 ;
        RECT -63.045 223.805 -62.545 224.035 ;
        RECT -64.990 221.270 -64.690 221.355 ;
        RECT -63.645 221.270 -63.345 221.445 ;
        RECT -63.045 221.355 -62.545 221.585 ;
        RECT -64.990 220.795 -63.345 221.270 ;
        RECT -64.990 220.695 -64.690 220.795 ;
        RECT -63.645 220.760 -63.345 220.795 ;
        RECT -63.045 220.375 -62.545 220.605 ;
        RECT -24.100 220.270 -18.930 220.510 ;
        RECT -9.965 220.270 -4.310 220.350 ;
        RECT -63.045 219.395 -62.545 219.625 ;
        RECT -62.860 212.490 -31.550 212.630 ;
        RECT -80.760 209.495 -80.145 209.725 ;
        RECT -80.760 209.195 -69.720 209.495 ;
        RECT -80.760 209.110 -80.145 209.195 ;
        RECT -78.925 208.790 -78.310 208.970 ;
        RECT -78.925 208.470 -69.900 208.790 ;
        RECT -62.860 208.780 -62.720 212.490 ;
        RECT -62.260 211.680 -32.150 211.820 ;
        RECT -62.260 209.405 -62.120 211.680 ;
        RECT -61.565 210.845 -32.845 211.025 ;
        RECT -61.565 210.230 -61.385 210.845 ;
        RECT -61.585 209.490 -61.345 210.230 ;
        RECT -78.925 208.460 -77.445 208.470 ;
        RECT -78.925 208.355 -78.305 208.460 ;
        RECT -77.400 208.205 -76.810 208.210 ;
        RECT -77.400 207.900 -69.920 208.205 ;
        RECT -62.920 208.060 -62.685 208.780 ;
        RECT -62.265 208.690 -62.030 209.405 ;
        RECT -77.400 207.560 -76.805 207.900 ;
        RECT -76.975 207.555 -76.805 207.560 ;
        RECT -66.020 203.245 -65.020 203.475 ;
        RECT -66.020 201.700 -65.020 201.930 ;
        RECT -66.020 196.380 -65.020 196.610 ;
        RECT -66.020 194.310 -65.020 194.540 ;
        RECT -66.020 188.245 -65.020 188.475 ;
        RECT -66.020 186.700 -65.020 186.930 ;
        RECT -66.020 181.380 -65.020 181.610 ;
        RECT -66.020 179.310 -65.020 179.540 ;
        RECT -62.860 176.825 -62.720 208.060 ;
        RECT -66.725 176.685 -62.720 176.825 ;
        RECT -66.725 174.830 -66.585 176.685 ;
        RECT -66.020 175.745 -65.020 175.975 ;
        RECT -66.730 174.135 -66.460 174.830 ;
        RECT -66.020 174.200 -65.020 174.430 ;
        RECT -66.715 169.440 -66.575 174.135 ;
        RECT -66.760 168.745 -66.490 169.440 ;
        RECT -66.020 168.880 -65.020 169.110 ;
        RECT -66.020 166.810 -65.020 167.040 ;
        RECT -62.260 164.495 -62.120 208.690 ;
        RECT -66.725 164.355 -62.120 164.495 ;
        RECT -66.725 162.330 -66.585 164.355 ;
        RECT -66.020 163.245 -65.020 163.475 ;
        RECT -66.730 161.635 -66.460 162.330 ;
        RECT -66.020 161.700 -65.020 161.930 ;
        RECT -66.715 156.940 -66.575 161.635 ;
        RECT -66.760 156.245 -66.490 156.940 ;
        RECT -66.020 156.380 -65.020 156.610 ;
        RECT -66.020 154.310 -65.020 154.540 ;
        RECT -61.565 152.075 -61.385 209.490 ;
        RECT -54.765 203.295 -53.765 203.525 ;
        RECT -40.645 203.295 -39.645 203.525 ;
        RECT -54.765 201.750 -53.765 201.980 ;
        RECT -40.645 201.750 -39.645 201.980 ;
        RECT -54.765 196.430 -53.765 196.660 ;
        RECT -40.645 196.430 -39.645 196.660 ;
        RECT -54.765 194.360 -53.765 194.590 ;
        RECT -40.645 194.360 -39.645 194.590 ;
        RECT -54.815 191.945 -53.315 192.175 ;
        RECT -41.095 191.945 -39.595 192.175 ;
        RECT -54.310 186.785 -53.310 187.015 ;
        RECT -41.100 186.785 -40.100 187.015 ;
        RECT -55.040 183.180 -53.540 183.410 ;
        RECT -40.870 183.180 -39.370 183.410 ;
        RECT -56.575 180.135 -56.075 180.365 ;
        RECT -38.335 180.135 -37.835 180.365 ;
        RECT -56.575 179.155 -56.075 179.385 ;
        RECT -38.335 179.155 -37.835 179.385 ;
        RECT -55.050 175.155 -53.550 175.385 ;
        RECT -40.860 175.155 -39.360 175.385 ;
        RECT -56.585 172.110 -56.085 172.340 ;
        RECT -38.325 172.110 -37.825 172.340 ;
        RECT -56.585 171.130 -56.085 171.360 ;
        RECT -38.325 171.130 -37.825 171.360 ;
        RECT -54.770 167.135 -53.270 167.365 ;
        RECT -41.140 167.135 -39.640 167.365 ;
        RECT -54.265 161.975 -53.265 162.205 ;
        RECT -41.145 161.975 -40.145 162.205 ;
        RECT -55.990 159.285 -55.490 159.515 ;
        RECT -38.920 159.285 -38.420 159.515 ;
        RECT -40.865 158.765 -40.565 158.865 ;
        RECT -39.520 158.765 -39.220 158.800 ;
        RECT -55.990 158.305 -55.490 158.535 ;
        RECT -40.865 158.290 -39.220 158.765 ;
        RECT -38.920 158.305 -38.420 158.535 ;
        RECT -55.190 158.115 -54.890 158.150 ;
        RECT -53.845 158.115 -53.545 158.215 ;
        RECT -40.865 158.205 -40.565 158.290 ;
        RECT -39.520 158.115 -39.220 158.290 ;
        RECT -55.190 157.640 -53.545 158.115 ;
        RECT -55.990 157.325 -55.490 157.555 ;
        RECT -55.190 157.465 -54.890 157.640 ;
        RECT -53.845 157.555 -53.545 157.640 ;
        RECT -38.920 157.325 -38.420 157.555 ;
        RECT -55.990 154.875 -55.490 155.105 ;
        RECT -38.920 154.875 -38.420 155.105 ;
        RECT -55.990 153.895 -55.490 154.125 ;
        RECT -38.920 153.895 -38.420 154.125 ;
        RECT -55.990 152.915 -55.490 153.145 ;
        RECT -38.920 152.915 -38.420 153.145 ;
        RECT -66.725 151.935 -61.385 152.075 ;
        RECT -33.025 152.075 -32.845 210.845 ;
        RECT -32.290 164.495 -32.150 211.680 ;
        RECT -31.690 176.825 -31.550 212.490 ;
        RECT -24.100 212.515 -3.985 220.270 ;
        RECT -24.100 212.350 -18.930 212.515 ;
        RECT -9.965 212.350 -4.310 212.515 ;
        RECT -29.390 203.245 -28.390 203.475 ;
        RECT -29.390 201.700 -28.390 201.930 ;
        RECT -29.390 196.380 -28.390 196.610 ;
        RECT -29.390 194.310 -28.390 194.540 ;
        RECT -29.390 188.245 -28.390 188.475 ;
        RECT -29.390 186.700 -28.390 186.930 ;
        RECT -29.390 181.380 -28.390 181.610 ;
        RECT -29.390 179.310 -28.390 179.540 ;
        RECT -31.690 176.685 -27.685 176.825 ;
        RECT -29.390 175.745 -28.390 175.975 ;
        RECT -27.825 174.830 -27.685 176.685 ;
        RECT -29.390 174.200 -28.390 174.430 ;
        RECT -27.950 174.135 -27.680 174.830 ;
        RECT -27.835 169.440 -27.695 174.135 ;
        RECT -29.390 168.880 -28.390 169.110 ;
        RECT -27.920 168.745 -27.650 169.440 ;
        RECT -29.390 166.810 -28.390 167.040 ;
        RECT -32.290 164.355 -27.685 164.495 ;
        RECT -29.390 163.245 -28.390 163.475 ;
        RECT -27.825 162.330 -27.685 164.355 ;
        RECT -29.390 161.700 -28.390 161.930 ;
        RECT -27.950 161.635 -27.680 162.330 ;
        RECT -27.835 156.940 -27.695 161.635 ;
        RECT -29.390 156.380 -28.390 156.610 ;
        RECT -27.920 156.245 -27.650 156.940 ;
        RECT -29.390 154.310 -28.390 154.540 ;
        RECT -33.025 151.935 -27.685 152.075 ;
        RECT -66.725 149.830 -66.585 151.935 ;
        RECT -66.020 150.745 -65.020 150.975 ;
        RECT -29.390 150.745 -28.390 150.975 ;
        RECT -52.700 149.855 -52.200 150.085 ;
        RECT -42.210 149.855 -41.710 150.085 ;
        RECT -27.825 149.830 -27.685 151.935 ;
        RECT -66.730 149.135 -66.460 149.830 ;
        RECT -66.020 149.200 -65.020 149.430 ;
        RECT -29.390 149.200 -28.390 149.430 ;
        RECT -27.950 149.135 -27.680 149.830 ;
        RECT -66.715 144.440 -66.575 149.135 ;
        RECT -52.700 148.875 -52.200 149.105 ;
        RECT -42.210 148.875 -41.710 149.105 ;
        RECT -52.700 147.895 -52.200 148.125 ;
        RECT -42.210 147.895 -41.710 148.125 ;
        RECT -55.990 146.160 -55.490 146.390 ;
        RECT -38.920 146.160 -38.420 146.390 ;
        RECT -52.700 145.670 -52.200 145.900 ;
        RECT -42.210 145.670 -41.710 145.900 ;
        RECT -55.990 145.180 -55.490 145.410 ;
        RECT -38.920 145.180 -38.420 145.410 ;
        RECT -55.185 144.895 -54.885 145.015 ;
        RECT -53.845 144.895 -53.545 145.050 ;
        RECT -66.760 143.745 -66.490 144.440 ;
        RECT -55.990 144.200 -55.490 144.430 ;
        RECT -55.185 144.420 -53.545 144.895 ;
        RECT -52.700 144.690 -52.200 144.920 ;
        RECT -42.210 144.690 -41.710 144.920 ;
        RECT -40.865 144.895 -40.565 145.050 ;
        RECT -39.525 144.895 -39.225 145.015 ;
        RECT -55.185 144.330 -54.885 144.420 ;
        RECT -53.845 144.365 -53.545 144.420 ;
        RECT -40.865 144.420 -39.225 144.895 ;
        RECT -27.835 144.440 -27.695 149.135 ;
        RECT -40.865 144.365 -40.565 144.420 ;
        RECT -39.525 144.330 -39.225 144.420 ;
        RECT -38.920 144.200 -38.420 144.430 ;
        RECT -66.020 143.880 -65.020 144.110 ;
        RECT -52.700 143.710 -52.200 143.940 ;
        RECT -42.210 143.710 -41.710 143.940 ;
        RECT -29.390 143.880 -28.390 144.110 ;
        RECT -27.920 143.745 -27.650 144.440 ;
        RECT -66.020 141.810 -65.020 142.040 ;
        RECT -29.390 141.810 -28.390 142.040 ;
        RECT -55.990 141.375 -55.490 141.605 ;
        RECT -38.920 141.375 -38.420 141.605 ;
        RECT -55.990 140.395 -55.490 140.625 ;
        RECT -38.920 140.395 -38.420 140.625 ;
        RECT -55.990 139.415 -55.490 139.645 ;
        RECT -38.920 139.415 -38.420 139.645 ;
        RECT -66.020 138.245 -65.020 138.475 ;
        RECT -29.390 138.245 -28.390 138.475 ;
        RECT -66.020 136.700 -65.020 136.930 ;
        RECT -29.390 136.700 -28.390 136.930 ;
        RECT -52.700 136.355 -52.200 136.585 ;
        RECT -42.210 136.355 -41.710 136.585 ;
        RECT -52.700 135.375 -52.200 135.605 ;
        RECT -42.210 135.375 -41.710 135.605 ;
        RECT -52.700 134.395 -52.200 134.625 ;
        RECT -42.210 134.395 -41.710 134.625 ;
        RECT -31.105 133.455 -30.605 133.685 ;
        RECT -55.990 132.660 -55.490 132.890 ;
        RECT -38.920 132.660 -38.420 132.890 ;
        RECT -31.105 132.475 -30.605 132.705 ;
        RECT -52.700 132.170 -52.200 132.400 ;
        RECT -42.210 132.170 -41.710 132.400 ;
        RECT -55.205 131.930 -54.905 131.995 ;
        RECT -53.815 131.930 -53.515 132.065 ;
        RECT -55.990 131.680 -55.490 131.910 ;
        RECT -66.020 131.380 -65.020 131.610 ;
        RECT -55.230 131.455 -53.515 131.930 ;
        RECT -55.990 130.700 -55.490 130.930 ;
        RECT -66.020 129.310 -65.020 129.540 ;
        RECT -55.230 129.495 -54.755 131.455 ;
        RECT -53.815 131.380 -53.515 131.455 ;
        RECT -40.895 131.930 -40.595 132.065 ;
        RECT -39.505 131.930 -39.205 131.995 ;
        RECT -40.895 131.455 -39.205 131.930 ;
        RECT -38.920 131.680 -38.420 131.910 ;
        RECT -31.105 131.495 -30.605 131.725 ;
        RECT -52.700 131.190 -52.200 131.420 ;
        RECT -42.210 131.190 -41.710 131.420 ;
        RECT -40.895 131.380 -40.595 131.455 ;
        RECT -39.505 131.335 -39.205 131.455 ;
        RECT -29.390 131.380 -28.390 131.610 ;
        RECT -38.920 130.700 -38.420 130.930 ;
        RECT -52.700 130.210 -52.200 130.440 ;
        RECT -42.210 130.210 -41.710 130.440 ;
        RECT -56.100 129.020 -54.755 129.495 ;
        RECT -29.390 129.310 -28.390 129.540 ;
        RECT -56.100 127.945 -55.625 129.020 ;
        RECT -55.110 125.390 -53.610 125.620 ;
        RECT -30.440 125.255 -28.940 125.485 ;
        RECT -55.110 124.410 -53.610 124.640 ;
        RECT -30.440 124.275 -28.940 124.505 ;
        RECT -55.110 123.200 -53.610 123.430 ;
        RECT -30.440 123.065 -28.940 123.295 ;
        RECT -33.910 121.420 -33.345 121.425 ;
        RECT -23.020 121.420 -22.070 205.585 ;
        RECT -33.910 120.945 -22.070 121.420 ;
        RECT -54.655 119.915 -54.155 120.145 ;
        RECT -54.655 118.935 -54.155 119.165 ;
        RECT -53.855 118.745 -53.555 118.780 ;
        RECT -52.510 118.745 -52.210 118.845 ;
        RECT -33.910 118.745 -33.345 120.945 ;
        RECT -30.020 119.915 -29.520 120.145 ;
        RECT -30.020 118.935 -29.520 119.165 ;
        RECT -53.855 118.270 -33.345 118.745 ;
        RECT -54.655 117.955 -54.155 118.185 ;
        RECT -53.855 118.095 -53.555 118.270 ;
        RECT -52.510 118.185 -52.210 118.270 ;
        RECT -54.655 115.505 -54.155 115.735 ;
        RECT -54.655 114.525 -54.155 114.755 ;
        RECT -54.655 113.545 -54.155 113.775 ;
        RECT -51.365 110.485 -50.865 110.715 ;
        RECT -33.910 109.970 -33.345 118.270 ;
        RECT -29.220 118.745 -28.920 118.780 ;
        RECT -28.675 118.745 -28.200 120.945 ;
        RECT -27.875 118.745 -27.575 118.845 ;
        RECT -29.220 118.270 -27.575 118.745 ;
        RECT -30.020 117.955 -29.520 118.185 ;
        RECT -29.220 118.095 -28.920 118.270 ;
        RECT -27.875 118.185 -27.575 118.270 ;
        RECT -30.020 115.505 -29.520 115.735 ;
        RECT -30.020 114.525 -29.520 114.755 ;
        RECT -30.020 113.545 -29.520 113.775 ;
        RECT -26.730 110.485 -26.230 110.715 ;
        RECT -51.365 109.505 -50.865 109.735 ;
        RECT -45.455 109.405 -33.345 109.970 ;
        RECT -26.730 109.505 -26.230 109.735 ;
        RECT -51.365 108.525 -50.865 108.755 ;
        RECT -54.655 106.790 -54.155 107.020 ;
        RECT -51.365 106.300 -50.865 106.530 ;
        RECT -45.455 106.430 -44.890 109.405 ;
        RECT -33.910 106.585 -33.345 109.405 ;
        RECT -26.730 108.525 -26.230 108.755 ;
        RECT -30.020 106.790 -29.520 107.020 ;
        RECT -26.730 106.300 -26.230 106.530 ;
        RECT -54.655 105.810 -54.155 106.040 ;
        RECT -35.950 105.880 -34.450 106.110 ;
        RECT -30.020 105.810 -29.520 106.040 ;
        RECT -53.850 105.525 -53.550 105.645 ;
        RECT -52.510 105.525 -52.210 105.680 ;
        RECT -54.655 104.830 -54.155 105.060 ;
        RECT -53.850 105.050 -52.210 105.525 ;
        RECT -51.365 105.320 -50.865 105.550 ;
        RECT -44.715 105.475 -44.215 105.705 ;
        RECT -29.215 105.525 -28.915 105.645 ;
        RECT -27.875 105.525 -27.575 105.680 ;
        RECT -53.850 104.960 -53.550 105.050 ;
        RECT -52.510 104.995 -52.210 105.050 ;
        RECT -51.365 104.340 -50.865 104.570 ;
        RECT -44.715 104.495 -44.215 104.725 ;
        RECT -35.950 104.670 -34.450 104.900 ;
        RECT -30.020 104.830 -29.520 105.060 ;
        RECT -29.215 105.050 -27.575 105.525 ;
        RECT -26.730 105.320 -26.230 105.550 ;
        RECT -29.215 104.960 -28.915 105.050 ;
        RECT -27.875 104.995 -27.575 105.050 ;
        RECT -26.730 104.340 -26.230 104.570 ;
        RECT -35.950 103.690 -34.450 103.920 ;
        RECT -54.655 102.005 -54.155 102.235 ;
        RECT -30.020 102.005 -29.520 102.235 ;
        RECT -47.250 101.450 -45.750 101.680 ;
        RECT -54.655 101.025 -54.155 101.255 ;
        RECT -30.020 101.025 -29.520 101.255 ;
        RECT -38.915 100.480 -38.415 100.710 ;
        RECT -54.655 100.045 -54.155 100.275 ;
        RECT -30.020 100.045 -29.520 100.275 ;
        RECT -38.915 99.500 -38.415 99.730 ;
        RECT -46.360 97.565 -45.360 97.795 ;
        RECT -51.365 96.985 -50.865 97.215 ;
        RECT -26.730 96.985 -26.230 97.215 ;
        RECT -46.360 96.585 -45.360 96.815 ;
        RECT -37.380 96.455 -35.880 96.685 ;
        RECT -51.365 96.005 -50.865 96.235 ;
        RECT -26.730 96.005 -26.230 96.235 ;
        RECT -51.365 95.025 -50.865 95.255 ;
        RECT -26.730 95.025 -26.230 95.255 ;
        RECT -54.655 93.290 -54.155 93.520 ;
        RECT -30.020 93.290 -29.520 93.520 ;
        RECT -51.365 92.800 -50.865 93.030 ;
        RECT -26.730 92.800 -26.230 93.030 ;
        RECT -53.870 92.560 -53.570 92.625 ;
        RECT -52.480 92.560 -52.180 92.695 ;
        RECT -54.655 92.310 -54.155 92.540 ;
        RECT -53.870 92.085 -52.180 92.560 ;
        RECT -29.235 92.560 -28.935 92.625 ;
        RECT -27.845 92.560 -27.545 92.695 ;
        RECT -30.020 92.310 -29.520 92.540 ;
        RECT -53.870 91.965 -53.570 92.085 ;
        RECT -52.480 92.010 -52.180 92.085 ;
        RECT -29.235 92.085 -27.545 92.560 ;
        RECT -51.365 91.820 -50.865 92.050 ;
        RECT -29.235 91.965 -28.935 92.085 ;
        RECT -27.845 92.010 -27.545 92.085 ;
        RECT -26.730 91.820 -26.230 92.050 ;
        RECT -54.655 91.330 -54.155 91.560 ;
        RECT -30.020 91.330 -29.520 91.560 ;
        RECT -51.365 90.840 -50.865 91.070 ;
        RECT -26.730 90.840 -26.230 91.070 ;
        RECT -65.575 84.495 -28.465 85.025 ;
        RECT -23.020 84.495 -22.070 120.945 ;
        RECT -65.575 84.460 -22.070 84.495 ;
        RECT -65.575 81.485 -65.010 84.460 ;
        RECT -54.030 81.640 -53.465 84.460 ;
        RECT -40.575 81.485 -40.010 84.460 ;
        RECT -29.030 83.545 -22.070 84.460 ;
        RECT -29.030 81.640 -28.465 83.545 ;
        RECT -56.070 80.935 -54.570 81.165 ;
        RECT -31.070 80.935 -29.570 81.165 ;
        RECT -64.835 80.530 -64.335 80.760 ;
        RECT -39.835 80.530 -39.335 80.760 ;
        RECT -64.835 79.550 -64.335 79.780 ;
        RECT -56.070 79.725 -54.570 79.955 ;
        RECT -39.835 79.550 -39.335 79.780 ;
        RECT -31.070 79.725 -29.570 79.955 ;
        RECT -56.070 78.745 -54.570 78.975 ;
        RECT -31.070 78.745 -29.570 78.975 ;
        RECT -67.370 76.505 -65.870 76.735 ;
        RECT -42.370 76.505 -40.870 76.735 ;
        RECT -59.035 75.535 -58.535 75.765 ;
        RECT -34.035 75.535 -33.535 75.765 ;
        RECT -59.035 74.555 -58.535 74.785 ;
        RECT -34.035 74.555 -33.535 74.785 ;
        RECT -66.480 72.620 -65.480 72.850 ;
        RECT -41.480 72.620 -40.480 72.850 ;
        RECT -66.480 71.640 -65.480 71.870 ;
        RECT -57.500 71.510 -56.000 71.740 ;
        RECT -41.480 71.640 -40.480 71.870 ;
        RECT -32.500 71.510 -31.000 71.740 ;
        RECT -42.485 67.645 -41.485 67.875 ;
        RECT -30.525 67.355 -30.025 67.585 ;
        RECT -30.525 66.375 -30.025 66.605 ;
        RECT -58.500 65.480 -57.500 65.710 ;
        RECT -58.500 64.500 -57.500 64.730 ;
        RECT -63.250 63.755 -62.565 63.840 ;
        RECT -57.710 63.755 -57.025 63.870 ;
        RECT -63.250 63.580 -57.025 63.755 ;
        RECT -63.250 63.550 -62.565 63.580 ;
        RECT -62.865 63.370 -62.180 63.375 ;
        RECT -56.850 63.370 -56.165 63.485 ;
        RECT -62.865 63.195 -56.165 63.370 ;
        RECT -33.060 63.330 -31.560 63.560 ;
        RECT -62.865 63.085 -62.180 63.195 ;
        RECT -42.480 62.485 -40.980 62.715 ;
        RECT -35.065 61.335 -34.405 61.410 ;
        RECT -30.855 61.335 -30.565 61.980 ;
        RECT -35.065 61.295 -30.565 61.335 ;
        RECT -58.495 60.955 -57.495 61.185 ;
        RECT -35.065 61.155 -30.650 61.295 ;
        RECT -35.065 61.145 -34.405 61.155 ;
        RECT -58.495 59.975 -57.495 60.205 ;
        RECT -62.470 59.200 -61.785 59.270 ;
        RECT -57.700 59.200 -57.015 59.280 ;
        RECT -62.470 58.990 -57.015 59.200 ;
        RECT -62.470 58.985 -57.035 58.990 ;
        RECT -62.470 58.980 -61.785 58.985 ;
        RECT -32.805 58.495 -31.805 58.725 ;
        RECT -66.445 57.910 -64.945 58.140 ;
        RECT -40.070 57.645 -39.570 57.875 ;
        RECT -64.075 57.080 -63.500 57.125 ;
        RECT -61.440 57.080 -60.690 57.295 ;
        RECT -64.075 56.645 -60.690 57.080 ;
        RECT -40.070 56.665 -39.570 56.895 ;
        RECT 84.745 56.750 86.410 84.195 ;
        RECT -64.075 56.455 -63.500 56.645 ;
        RECT -61.440 56.455 -60.690 56.645 ;
        RECT -64.075 56.020 -60.690 56.455 ;
        RECT -64.075 55.535 -63.500 56.020 ;
        RECT -61.440 55.535 -60.690 56.020 ;
        RECT -64.075 55.100 -60.690 55.535 ;
        RECT -64.075 54.670 -63.500 55.100 ;
        RECT -61.440 54.670 -60.690 55.100 ;
        RECT -60.210 54.925 -59.210 55.155 ;
        RECT -64.075 54.235 -60.690 54.670 ;
        RECT -64.075 53.770 -63.500 54.235 ;
        RECT -61.440 53.770 -60.690 54.235 ;
        RECT -60.210 53.945 -59.210 54.175 ;
        RECT -64.075 53.335 -60.690 53.770 ;
        RECT -42.605 53.620 -41.105 53.850 ;
        RECT -32.800 53.335 -31.300 53.565 ;
        RECT -65.940 52.750 -64.940 52.980 ;
        RECT -64.075 52.210 -63.500 53.335 ;
        RECT -61.440 53.275 -60.690 53.335 ;
        RECT -80.785 51.300 -80.170 51.530 ;
        RECT -80.785 51.000 -39.200 51.300 ;
        RECT -80.785 50.915 -80.170 51.000 ;
        RECT 79.665 50.890 80.090 50.895 ;
        RECT -78.950 50.595 -78.335 50.775 ;
        RECT 79.665 50.660 81.090 50.890 ;
        RECT 84.090 50.660 85.090 50.890 ;
        RECT -78.950 50.275 -41.355 50.595 ;
        RECT -78.950 50.265 -77.470 50.275 ;
        RECT -78.950 50.160 -78.330 50.265 ;
        RECT -77.425 50.010 -76.835 50.015 ;
        RECT -77.425 49.705 -33.995 50.010 ;
        RECT -77.425 49.365 -76.830 49.705 ;
        RECT -77.000 49.360 -76.830 49.365 ;
        RECT 79.665 48.315 79.895 50.660 ;
        RECT 79.665 48.310 80.090 48.315 ;
        RECT 79.665 48.080 81.090 48.310 ;
        RECT 84.090 48.080 85.090 48.310 ;
        RECT 79.665 45.730 79.895 48.080 ;
        RECT 79.665 45.500 81.090 45.730 ;
        RECT 84.090 45.500 85.090 45.730 ;
        RECT 80.215 45.060 80.505 45.500 ;
        RECT 85.655 45.060 86.590 45.905 ;
        RECT 80.165 44.830 86.590 45.060 ;
        RECT 86.010 44.780 86.590 44.830 ;
        RECT -81.385 42.470 -27.190 42.775 ;
        RECT -81.385 40.160 -27.165 42.470 ;
        RECT -32.700 36.365 -27.165 40.160 ;
        RECT 133.765 38.115 190.365 44.220 ;
        RECT 40.870 28.215 41.100 32.215 ;
        RECT 49.450 28.215 49.680 32.215 ;
        RECT 58.030 28.215 58.260 32.215 ;
        RECT 40.870 23.215 41.100 27.215 ;
        RECT 49.450 23.215 49.680 27.215 ;
        RECT 58.030 23.215 58.260 27.215 ;
        RECT 14.330 20.580 16.250 22.800 ;
        RECT 15.305 12.540 16.175 20.580 ;
        RECT 134.180 19.430 140.145 38.115 ;
        RECT 145.555 19.430 151.520 38.115 ;
        RECT 156.375 19.430 162.340 38.115 ;
        RECT 169.420 19.430 175.385 38.115 ;
        RECT 181.905 19.430 187.870 38.115 ;
        RECT 132.915 17.415 194.330 19.430 ;
        RECT 98.940 14.490 99.170 14.990 ;
        RECT 99.920 14.490 100.150 14.990 ;
        RECT 100.900 14.490 101.130 14.990 ;
        RECT 103.190 14.490 103.420 14.990 ;
        RECT 104.170 14.490 104.400 14.990 ;
        RECT 105.150 14.490 105.380 14.990 ;
        RECT 97.760 14.310 98.250 14.460 ;
        RECT 97.760 14.290 98.295 14.310 ;
        RECT 97.760 13.935 101.570 14.290 ;
        RECT 14.045 11.960 16.175 12.540 ;
        RECT 103.190 12.415 103.420 12.915 ;
        RECT 104.170 12.415 104.400 12.915 ;
        RECT 105.150 12.415 105.380 12.915 ;
        RECT 11.955 11.780 16.175 11.960 ;
        RECT 3.535 10.005 3.765 10.425 ;
        RECT 6.095 9.950 6.325 10.550 ;
        RECT 7.545 9.975 7.775 10.575 ;
        RECT 9.705 9.850 9.935 10.610 ;
        RECT 10.885 9.850 11.115 10.610 ;
        RECT 11.955 9.850 12.135 11.780 ;
        RECT 14.045 11.360 16.175 11.780 ;
        RECT 12.470 10.005 12.700 10.425 ;
        RECT 14.015 9.850 14.245 10.425 ;
        RECT 9.705 9.670 14.245 9.850 ;
        RECT 15.305 5.795 16.175 11.360 ;
        RECT 151.620 10.480 151.850 12.480 ;
        RECT 153.200 10.480 153.430 12.480 ;
        RECT 154.780 10.480 155.010 12.480 ;
        RECT 155.570 10.480 155.800 12.480 ;
        RECT 156.360 10.480 156.590 12.480 ;
        RECT 157.150 10.480 157.380 12.480 ;
        RECT 157.940 10.480 158.170 12.480 ;
        RECT 175.295 10.590 175.525 12.590 ;
        RECT 176.875 10.590 177.105 12.590 ;
        RECT 178.455 10.590 178.685 12.590 ;
        RECT 179.245 10.590 179.475 12.590 ;
        RECT 180.035 10.590 180.265 12.590 ;
        RECT 180.825 10.590 181.055 12.590 ;
        RECT 181.615 10.590 181.845 12.590 ;
        RECT 183.900 10.375 184.130 12.375 ;
        RECT 185.480 10.375 185.710 12.375 ;
        RECT 187.060 10.375 187.290 12.375 ;
        RECT 187.850 10.375 188.080 12.375 ;
        RECT 188.640 10.375 188.870 12.375 ;
        RECT 189.430 10.375 189.660 12.375 ;
        RECT 190.220 10.375 190.450 12.375 ;
        RECT 195.900 12.275 196.130 12.775 ;
        RECT 196.880 12.275 197.110 12.775 ;
        RECT 197.860 12.275 198.090 12.775 ;
        RECT 200.310 12.275 200.540 12.775 ;
        RECT 201.290 12.275 201.520 12.775 ;
        RECT 202.270 12.275 202.500 12.775 ;
        RECT 209.025 12.275 209.255 12.775 ;
        RECT 210.005 12.275 210.235 12.775 ;
        RECT 210.985 12.275 211.215 12.775 ;
        RECT 213.810 12.275 214.040 12.775 ;
        RECT 214.790 12.275 215.020 12.775 ;
        RECT 215.770 12.275 216.000 12.775 ;
        RECT 222.525 12.275 222.755 12.775 ;
        RECT 223.505 12.275 223.735 12.775 ;
        RECT 224.485 12.275 224.715 12.775 ;
        RECT 194.025 12.035 194.705 12.040 ;
        RECT 193.900 11.440 194.860 12.035 ;
        RECT 197.265 11.675 197.950 11.975 ;
        RECT 197.300 11.440 197.775 11.675 ;
        RECT 210.400 11.670 211.085 11.970 ;
        RECT 223.420 11.895 224.080 11.990 ;
        RECT 229.020 11.895 229.750 12.205 ;
        RECT 223.420 11.690 229.750 11.895 ;
        RECT 223.485 11.675 229.750 11.690 ;
        RECT 193.900 10.965 197.775 11.440 ;
        RECT 193.900 10.745 194.860 10.965 ;
        RECT 197.300 10.630 197.775 10.965 ;
        RECT 210.520 10.630 210.995 11.670 ;
        RECT 197.200 10.330 197.860 10.630 ;
        RECT 210.365 10.330 211.050 10.630 ;
        RECT 223.485 10.600 223.960 11.675 ;
        RECT 229.020 11.275 229.750 11.675 ;
        RECT 223.350 10.300 224.035 10.600 ;
        RECT 22.545 8.665 22.775 9.165 ;
        RECT 23.525 8.665 23.755 9.165 ;
        RECT 24.505 8.665 24.735 9.165 ;
        RECT 26.795 8.665 27.025 9.165 ;
        RECT 27.775 8.665 28.005 9.165 ;
        RECT 28.755 8.665 28.985 9.165 ;
        RECT 205.330 8.985 205.560 9.485 ;
        RECT 206.310 8.985 206.540 9.485 ;
        RECT 207.290 8.985 207.520 9.485 ;
        RECT 209.515 8.985 209.745 9.485 ;
        RECT 210.495 8.985 210.725 9.485 ;
        RECT 211.475 8.985 211.705 9.485 ;
        RECT 218.830 8.985 219.060 9.485 ;
        RECT 219.810 8.985 220.040 9.485 ;
        RECT 220.790 8.985 221.020 9.485 ;
        RECT 223.015 8.985 223.245 9.485 ;
        RECT 223.995 8.985 224.225 9.485 ;
        RECT 224.975 8.985 225.205 9.485 ;
        RECT 227.865 9.435 228.095 9.935 ;
        RECT 228.845 9.435 229.075 9.935 ;
        RECT 229.825 9.435 230.055 9.935 ;
        RECT 255.910 9.130 256.140 11.130 ;
        RECT 257.090 9.130 257.320 11.130 ;
        RECT 258.270 9.130 258.500 11.130 ;
        RECT 259.450 9.130 259.680 11.130 ;
        RECT 260.630 9.130 260.860 11.130 ;
        RECT 261.810 9.130 262.040 11.130 ;
        RECT 262.990 9.130 263.220 11.130 ;
        RECT 264.170 9.130 264.400 11.130 ;
        RECT 265.350 9.130 265.580 11.130 ;
        RECT 266.530 9.130 266.760 11.130 ;
        RECT 267.710 9.130 267.940 11.130 ;
        RECT 268.890 9.130 269.120 11.130 ;
        RECT 270.070 9.130 270.300 11.130 ;
        RECT 271.250 9.130 271.480 11.130 ;
        RECT 272.430 9.130 272.660 11.130 ;
        RECT 273.610 9.130 273.840 11.130 ;
        RECT 274.200 9.130 274.430 11.130 ;
        RECT 274.790 9.130 275.020 11.130 ;
        RECT 275.380 9.130 275.610 11.130 ;
        RECT 275.970 9.130 276.200 11.130 ;
        RECT 276.560 9.130 276.790 11.130 ;
        RECT 277.150 9.130 277.380 11.130 ;
        RECT 277.740 9.130 277.970 11.130 ;
        RECT 278.330 9.130 278.560 11.130 ;
        RECT 278.920 9.130 279.150 11.130 ;
        RECT 279.510 9.130 279.740 11.130 ;
        RECT 280.100 9.130 280.330 11.130 ;
        RECT 280.690 9.130 280.920 11.130 ;
        RECT 281.280 9.130 281.510 11.130 ;
        RECT 281.870 9.130 282.100 11.130 ;
        RECT 282.460 9.130 282.690 11.130 ;
        RECT 283.050 9.130 283.280 11.130 ;
        RECT 283.640 9.130 283.870 11.130 ;
        RECT 284.230 9.130 284.460 11.130 ;
        RECT 284.820 9.130 285.050 11.130 ;
        RECT 285.410 9.130 285.640 11.130 ;
        RECT 286.000 9.130 286.230 11.130 ;
        RECT 286.590 9.130 286.820 11.130 ;
        RECT 287.180 9.130 287.410 11.130 ;
        RECT 287.770 9.130 288.000 11.130 ;
        RECT 288.360 9.130 288.590 11.130 ;
        RECT 288.950 9.130 289.180 11.130 ;
        RECT 289.540 9.130 289.770 11.130 ;
        RECT 290.130 9.130 290.360 11.130 ;
        RECT 290.720 9.130 290.950 11.130 ;
        RECT 291.310 9.130 291.540 11.130 ;
        RECT 20.930 6.925 24.815 7.595 ;
        RECT 22.900 6.920 24.135 6.925 ;
        RECT 26.795 6.590 27.025 7.090 ;
        RECT 27.775 6.590 28.005 7.090 ;
        RECT 28.755 6.590 28.985 7.090 ;
        RECT 15.305 5.505 19.495 5.795 ;
        RECT 9.705 4.460 14.245 4.640 ;
        RECT 3.535 3.885 3.765 4.305 ;
        RECT 6.095 3.760 6.325 4.360 ;
        RECT 7.545 3.735 7.775 4.335 ;
        RECT 9.705 3.700 9.935 4.460 ;
        RECT 10.885 3.700 11.115 4.460 ;
        RECT 11.955 2.530 12.135 4.460 ;
        RECT 12.470 3.885 12.700 4.305 ;
        RECT 14.015 3.885 14.245 4.460 ;
        RECT 15.305 2.945 16.175 5.505 ;
        RECT 13.970 2.530 16.175 2.945 ;
        RECT 11.955 2.350 16.175 2.530 ;
        RECT 13.970 2.195 16.175 2.350 ;
        RECT 13.970 1.775 15.495 2.195 ;
        RECT 19.205 -5.055 19.495 5.505 ;
        RECT 39.520 5.245 39.750 7.245 ;
        RECT 40.700 5.245 40.930 7.245 ;
        RECT 41.880 5.245 42.110 7.245 ;
        RECT 43.060 5.245 43.290 7.245 ;
        RECT 44.240 5.245 44.470 7.245 ;
        RECT 45.420 5.245 45.650 7.245 ;
        RECT 46.600 5.245 46.830 7.245 ;
        RECT 47.780 5.245 48.010 7.245 ;
        RECT 48.960 5.245 49.190 7.245 ;
        RECT 50.140 5.245 50.370 7.245 ;
        RECT 51.320 5.245 51.550 7.245 ;
        RECT 52.500 5.245 52.730 7.245 ;
        RECT 53.680 5.245 53.910 7.245 ;
        RECT 54.860 5.245 55.090 7.245 ;
        RECT 56.040 5.245 56.270 7.245 ;
        RECT 57.220 5.245 57.450 7.245 ;
        RECT 57.810 5.245 58.040 7.245 ;
        RECT 58.400 5.245 58.630 7.245 ;
        RECT 58.990 5.245 59.220 7.245 ;
        RECT 59.580 5.245 59.810 7.245 ;
        RECT 60.170 5.245 60.400 7.245 ;
        RECT 60.760 5.245 60.990 7.245 ;
        RECT 61.350 5.245 61.580 7.245 ;
        RECT 61.940 5.245 62.170 7.245 ;
        RECT 62.530 5.245 62.760 7.245 ;
        RECT 63.120 5.245 63.350 7.245 ;
        RECT 63.710 5.245 63.940 7.245 ;
        RECT 64.300 5.245 64.530 7.245 ;
        RECT 64.890 5.245 65.120 7.245 ;
        RECT 65.480 5.245 65.710 7.245 ;
        RECT 66.070 5.245 66.300 7.245 ;
        RECT 66.660 5.245 66.890 7.245 ;
        RECT 67.250 5.245 67.480 7.245 ;
        RECT 67.840 5.245 68.070 7.245 ;
        RECT 68.430 5.245 68.660 7.245 ;
        RECT 69.020 5.245 69.250 7.245 ;
        RECT 69.610 5.245 69.840 7.245 ;
        RECT 70.200 5.245 70.430 7.245 ;
        RECT 70.790 5.245 71.020 7.245 ;
        RECT 71.380 5.245 71.610 7.245 ;
        RECT 71.970 5.245 72.200 7.245 ;
        RECT 72.560 5.245 72.790 7.245 ;
        RECT 73.150 5.245 73.380 7.245 ;
        RECT 73.740 5.245 73.970 7.245 ;
        RECT 74.330 5.245 74.560 7.245 ;
        RECT 74.920 5.245 75.150 7.245 ;
        RECT 112.180 6.205 114.625 6.585 ;
        RECT 97.360 4.715 114.625 6.205 ;
        RECT 97.360 -2.480 97.710 4.715 ;
        RECT 112.180 4.475 114.625 4.715 ;
        RECT 139.050 1.990 139.280 5.705 ;
        RECT 139.840 2.445 140.070 5.705 ;
        RECT 145.580 4.685 145.810 5.685 ;
        RECT 146.370 4.685 146.600 5.685 ;
        RECT 145.575 2.445 145.805 3.445 ;
        RECT 138.445 1.760 139.280 1.990 ;
        RECT 146.365 1.845 146.595 3.445 ;
        RECT 163.325 1.955 163.555 5.670 ;
        RECT 164.115 2.410 164.345 5.670 ;
        RECT 169.855 4.650 170.085 5.650 ;
        RECT 170.645 4.650 170.875 5.650 ;
        RECT 169.850 2.410 170.080 3.410 ;
        RECT 137.655 -0.115 137.885 0.885 ;
        RECT 138.445 -0.115 138.675 1.760 ;
        RECT 146.365 1.615 147.730 1.845 ;
        RECT 139.805 -0.105 140.035 0.895 ;
        RECT 141.385 -0.105 141.615 0.895 ;
        RECT 142.965 -0.105 143.195 0.895 ;
        RECT 144.545 -0.105 144.775 0.895 ;
        RECT 146.125 -0.105 146.355 0.895 ;
        RECT 147.500 -0.105 147.730 1.615 ;
        RECT 162.720 1.725 163.555 1.955 ;
        RECT 170.640 1.810 170.870 3.410 ;
        RECT 148.290 -0.105 148.520 0.895 ;
        RECT 151.620 -1.080 151.850 0.920 ;
        RECT 153.200 -1.080 153.430 0.920 ;
        RECT 154.780 -1.080 155.010 0.920 ;
        RECT 155.570 -1.080 155.800 0.920 ;
        RECT 156.360 -1.080 156.590 0.920 ;
        RECT 157.150 -1.080 157.380 0.920 ;
        RECT 157.940 -1.080 158.170 0.920 ;
        RECT 161.930 -0.150 162.160 0.850 ;
        RECT 162.720 -0.150 162.950 1.725 ;
        RECT 170.640 1.580 172.005 1.810 ;
        RECT 164.080 -0.140 164.310 0.860 ;
        RECT 165.660 -0.140 165.890 0.860 ;
        RECT 167.240 -0.140 167.470 0.860 ;
        RECT 168.820 -0.140 169.050 0.860 ;
        RECT 170.400 -0.140 170.630 0.860 ;
        RECT 171.775 -0.140 172.005 1.580 ;
        RECT 172.565 -0.140 172.795 0.860 ;
        RECT 175.295 -0.965 175.525 1.035 ;
        RECT 176.875 -0.965 177.105 1.035 ;
        RECT 178.455 -0.965 178.685 1.035 ;
        RECT 179.245 -0.965 179.475 1.035 ;
        RECT 180.035 -0.965 180.265 1.035 ;
        RECT 180.825 -0.965 181.055 1.035 ;
        RECT 181.615 -0.965 181.845 1.035 ;
        RECT 183.900 -0.750 184.130 1.250 ;
        RECT 185.480 -0.750 185.710 1.250 ;
        RECT 187.060 -0.750 187.290 1.250 ;
        RECT 187.850 -0.750 188.080 1.250 ;
        RECT 188.640 -0.750 188.870 1.250 ;
        RECT 189.430 -0.750 189.660 1.250 ;
        RECT 190.220 -0.750 190.450 1.250 ;
        RECT 99.800 -2.260 100.030 -1.760 ;
        RECT 100.780 -2.260 101.010 -1.760 ;
        RECT 101.760 -2.260 101.990 -1.760 ;
        RECT 104.050 -2.260 104.280 -1.760 ;
        RECT 105.030 -2.260 105.260 -1.760 ;
        RECT 106.010 -2.260 106.240 -1.760 ;
        RECT 97.360 -2.830 102.585 -2.480 ;
        RECT 22.620 -4.785 22.850 -4.285 ;
        RECT 23.600 -4.785 23.830 -4.285 ;
        RECT 24.580 -4.785 24.810 -4.285 ;
        RECT 26.870 -4.785 27.100 -4.285 ;
        RECT 27.850 -4.785 28.080 -4.285 ;
        RECT 28.830 -4.785 29.060 -4.285 ;
        RECT 104.050 -4.335 104.280 -3.835 ;
        RECT 105.030 -4.335 105.260 -3.835 ;
        RECT 106.010 -4.335 106.240 -3.835 ;
        RECT 19.205 -5.330 24.995 -5.055 ;
        RECT 19.205 -5.345 23.005 -5.330 ;
        RECT 254.895 -5.425 255.125 -3.425 ;
        RECT 256.075 -5.425 256.305 -3.425 ;
        RECT 257.255 -5.425 257.485 -3.425 ;
        RECT 258.435 -5.425 258.665 -3.425 ;
        RECT 259.615 -5.425 259.845 -3.425 ;
        RECT 260.795 -5.425 261.025 -3.425 ;
        RECT 261.975 -5.425 262.205 -3.425 ;
        RECT 263.155 -5.425 263.385 -3.425 ;
        RECT 264.335 -5.425 264.565 -3.425 ;
        RECT 265.515 -5.425 265.745 -3.425 ;
        RECT 266.695 -5.425 266.925 -3.425 ;
        RECT 267.875 -5.425 268.105 -3.425 ;
        RECT 269.055 -5.425 269.285 -3.425 ;
        RECT 270.235 -5.425 270.465 -3.425 ;
        RECT 271.415 -5.425 271.645 -3.425 ;
        RECT 272.595 -5.425 272.825 -3.425 ;
        RECT 273.185 -5.425 273.415 -3.425 ;
        RECT 273.775 -5.425 274.005 -3.425 ;
        RECT 274.365 -5.425 274.595 -3.425 ;
        RECT 274.955 -5.425 275.185 -3.425 ;
        RECT 275.545 -5.425 275.775 -3.425 ;
        RECT 276.135 -5.425 276.365 -3.425 ;
        RECT 276.725 -5.425 276.955 -3.425 ;
        RECT 277.315 -5.425 277.545 -3.425 ;
        RECT 277.905 -5.425 278.135 -3.425 ;
        RECT 278.495 -5.425 278.725 -3.425 ;
        RECT 279.085 -5.425 279.315 -3.425 ;
        RECT 279.675 -5.425 279.905 -3.425 ;
        RECT 280.265 -5.425 280.495 -3.425 ;
        RECT 280.855 -5.425 281.085 -3.425 ;
        RECT 281.445 -5.425 281.675 -3.425 ;
        RECT 282.035 -5.425 282.265 -3.425 ;
        RECT 282.625 -5.425 282.855 -3.425 ;
        RECT 283.215 -5.425 283.445 -3.425 ;
        RECT 283.805 -5.425 284.035 -3.425 ;
        RECT 284.395 -5.425 284.625 -3.425 ;
        RECT 284.985 -5.425 285.215 -3.425 ;
        RECT 285.575 -5.425 285.805 -3.425 ;
        RECT 286.165 -5.425 286.395 -3.425 ;
        RECT 286.755 -5.425 286.985 -3.425 ;
        RECT 287.345 -5.425 287.575 -3.425 ;
        RECT 287.935 -5.425 288.165 -3.425 ;
        RECT 288.525 -5.425 288.755 -3.425 ;
        RECT 289.115 -5.425 289.345 -3.425 ;
        RECT 289.705 -5.425 289.935 -3.425 ;
        RECT 290.295 -5.425 290.525 -3.425 ;
        RECT 26.870 -6.860 27.100 -6.360 ;
        RECT 27.850 -6.860 28.080 -6.360 ;
        RECT 28.830 -6.860 29.060 -6.360 ;
        RECT 39.315 -8.535 39.545 -6.535 ;
        RECT 40.495 -8.535 40.725 -6.535 ;
        RECT 41.675 -8.535 41.905 -6.535 ;
        RECT 42.855 -8.535 43.085 -6.535 ;
        RECT 44.035 -8.535 44.265 -6.535 ;
        RECT 45.215 -8.535 45.445 -6.535 ;
        RECT 46.395 -8.535 46.625 -6.535 ;
        RECT 47.575 -8.535 47.805 -6.535 ;
        RECT 48.755 -8.535 48.985 -6.535 ;
        RECT 49.935 -8.535 50.165 -6.535 ;
        RECT 51.115 -8.535 51.345 -6.535 ;
        RECT 52.295 -8.535 52.525 -6.535 ;
        RECT 53.475 -8.535 53.705 -6.535 ;
        RECT 54.655 -8.535 54.885 -6.535 ;
        RECT 55.835 -8.535 56.065 -6.535 ;
        RECT 57.015 -8.535 57.245 -6.535 ;
        RECT 57.605 -8.535 57.835 -6.535 ;
        RECT 58.195 -8.535 58.425 -6.535 ;
        RECT 58.785 -8.535 59.015 -6.535 ;
        RECT 59.375 -8.535 59.605 -6.535 ;
        RECT 59.965 -8.535 60.195 -6.535 ;
        RECT 60.555 -8.535 60.785 -6.535 ;
        RECT 61.145 -8.535 61.375 -6.535 ;
        RECT 61.735 -8.535 61.965 -6.535 ;
        RECT 62.325 -8.535 62.555 -6.535 ;
        RECT 62.915 -8.535 63.145 -6.535 ;
        RECT 63.505 -8.535 63.735 -6.535 ;
        RECT 64.095 -8.535 64.325 -6.535 ;
        RECT 64.685 -8.535 64.915 -6.535 ;
        RECT 65.275 -8.535 65.505 -6.535 ;
        RECT 65.865 -8.535 66.095 -6.535 ;
        RECT 66.455 -8.535 66.685 -6.535 ;
        RECT 67.045 -8.535 67.275 -6.535 ;
        RECT 67.635 -8.535 67.865 -6.535 ;
        RECT 68.225 -8.535 68.455 -6.535 ;
        RECT 68.815 -8.535 69.045 -6.535 ;
        RECT 69.405 -8.535 69.635 -6.535 ;
        RECT 69.995 -8.535 70.225 -6.535 ;
        RECT 70.585 -8.535 70.815 -6.535 ;
        RECT 71.175 -8.535 71.405 -6.535 ;
        RECT 71.765 -8.535 71.995 -6.535 ;
        RECT 72.355 -8.535 72.585 -6.535 ;
        RECT 72.945 -8.535 73.175 -6.535 ;
        RECT 73.535 -8.535 73.765 -6.535 ;
        RECT 74.125 -8.535 74.355 -6.535 ;
        RECT 74.715 -8.535 74.945 -6.535 ;
        RECT 234.250 -23.350 237.060 -9.800 ;
        RECT 306.765 -16.465 310.880 -16.140 ;
        RECT 254.895 -20.660 255.125 -18.660 ;
        RECT 256.075 -20.660 256.305 -18.660 ;
        RECT 257.255 -20.660 257.485 -18.660 ;
        RECT 258.435 -20.660 258.665 -18.660 ;
        RECT 259.615 -20.660 259.845 -18.660 ;
        RECT 260.795 -20.660 261.025 -18.660 ;
        RECT 261.975 -20.660 262.205 -18.660 ;
        RECT 263.155 -20.660 263.385 -18.660 ;
        RECT 264.335 -20.660 264.565 -18.660 ;
        RECT 265.515 -20.660 265.745 -18.660 ;
        RECT 266.695 -20.660 266.925 -18.660 ;
        RECT 267.875 -20.660 268.105 -18.660 ;
        RECT 269.055 -20.660 269.285 -18.660 ;
        RECT 270.235 -20.660 270.465 -18.660 ;
        RECT 271.415 -20.660 271.645 -18.660 ;
        RECT 272.595 -20.660 272.825 -18.660 ;
        RECT 273.185 -20.660 273.415 -18.660 ;
        RECT 273.775 -20.660 274.005 -18.660 ;
        RECT 274.365 -20.660 274.595 -18.660 ;
        RECT 274.955 -20.660 275.185 -18.660 ;
        RECT 275.545 -20.660 275.775 -18.660 ;
        RECT 276.135 -20.660 276.365 -18.660 ;
        RECT 276.725 -20.660 276.955 -18.660 ;
        RECT 277.315 -20.660 277.545 -18.660 ;
        RECT 277.905 -20.660 278.135 -18.660 ;
        RECT 278.495 -20.660 278.725 -18.660 ;
        RECT 279.085 -20.660 279.315 -18.660 ;
        RECT 279.675 -20.660 279.905 -18.660 ;
        RECT 280.265 -20.660 280.495 -18.660 ;
        RECT 280.855 -20.660 281.085 -18.660 ;
        RECT 281.445 -20.660 281.675 -18.660 ;
        RECT 282.035 -20.660 282.265 -18.660 ;
        RECT 282.625 -20.660 282.855 -18.660 ;
        RECT 283.215 -20.660 283.445 -18.660 ;
        RECT 283.805 -20.660 284.035 -18.660 ;
        RECT 284.395 -20.660 284.625 -18.660 ;
        RECT 284.985 -20.660 285.215 -18.660 ;
        RECT 285.575 -20.660 285.805 -18.660 ;
        RECT 286.165 -20.660 286.395 -18.660 ;
        RECT 286.755 -20.660 286.985 -18.660 ;
        RECT 287.345 -20.660 287.575 -18.660 ;
        RECT 287.935 -20.660 288.165 -18.660 ;
        RECT 288.525 -20.660 288.755 -18.660 ;
        RECT 289.115 -20.660 289.345 -18.660 ;
        RECT 289.705 -20.660 289.935 -18.660 ;
        RECT 290.295 -20.660 290.525 -18.660 ;
        RECT 233.890 -26.520 237.060 -23.350 ;
        RECT 306.765 -23.895 307.090 -16.465 ;
        RECT 310.555 -16.800 310.880 -16.465 ;
        RECT 311.935 -16.590 312.165 -16.090 ;
        RECT 312.915 -16.590 313.145 -16.090 ;
        RECT 313.895 -16.590 314.125 -16.090 ;
        RECT 316.185 -16.590 316.415 -16.090 ;
        RECT 317.165 -16.590 317.395 -16.090 ;
        RECT 318.145 -16.590 318.375 -16.090 ;
        RECT 310.555 -17.125 314.550 -16.800 ;
        RECT 311.935 -17.155 314.550 -17.125 ;
        RECT 316.185 -18.665 316.415 -18.165 ;
        RECT 317.165 -18.665 317.395 -18.165 ;
        RECT 318.145 -18.665 318.375 -18.165 ;
        RECT 306.305 -25.205 307.410 -23.895 ;
        RECT 449.950 -38.335 464.795 -23.490 ;
        RECT 450.595 -271.390 463.655 -38.335 ;
      LAYER met2 ;
        RECT 84.745 56.750 86.410 84.195 ;
      LAYER met3 ;
        RECT 91.300 419.320 116.700 446.180 ;
        RECT 117.900 419.320 143.300 446.180 ;
        RECT 144.500 419.320 169.900 446.180 ;
        RECT 171.100 419.320 196.500 446.180 ;
        RECT 197.700 419.320 223.100 446.180 ;
        RECT 224.300 419.320 249.700 446.180 ;
        RECT 250.900 419.320 276.300 446.180 ;
        RECT 277.500 419.320 302.900 446.180 ;
        RECT 304.100 419.320 329.500 446.180 ;
        RECT 330.700 419.320 356.100 446.180 ;
        RECT 357.300 419.320 382.700 446.180 ;
        RECT 383.900 419.320 409.300 446.180 ;
        RECT 410.500 419.320 435.900 446.180 ;
        RECT 437.100 419.320 462.500 446.180 ;
        RECT 91.300 391.260 116.700 418.120 ;
        RECT 117.900 391.260 143.300 418.120 ;
        RECT 144.500 391.260 169.900 418.120 ;
        RECT 171.100 391.260 196.500 418.120 ;
        RECT 197.700 391.260 223.100 418.120 ;
        RECT 224.300 391.260 249.700 418.120 ;
        RECT 250.900 391.260 276.300 418.120 ;
        RECT 277.500 391.260 302.900 418.120 ;
        RECT 304.100 391.260 329.500 418.120 ;
        RECT 330.700 391.260 356.100 418.120 ;
        RECT 357.300 391.260 382.700 418.120 ;
        RECT 383.900 391.260 409.300 418.120 ;
        RECT 410.500 391.260 435.900 418.120 ;
        RECT 437.100 391.260 462.500 418.120 ;
        RECT 91.300 363.200 116.700 390.060 ;
        RECT 117.900 363.200 143.300 390.060 ;
        RECT 144.500 363.200 169.900 390.060 ;
        RECT 171.100 363.200 196.500 390.060 ;
        RECT 197.700 363.200 223.100 390.060 ;
        RECT 224.300 363.200 249.700 390.060 ;
        RECT 250.900 363.200 276.300 390.060 ;
        RECT 277.500 363.200 302.900 390.060 ;
        RECT 304.100 363.200 329.500 390.060 ;
        RECT 330.700 363.200 356.100 390.060 ;
        RECT 357.300 363.200 382.700 390.060 ;
        RECT 383.900 363.200 409.300 390.060 ;
        RECT 410.500 363.200 435.900 390.060 ;
        RECT 437.100 363.200 462.500 390.060 ;
        RECT 91.300 335.140 116.700 362.000 ;
        RECT 117.900 335.140 143.300 362.000 ;
        RECT 144.500 335.140 169.900 362.000 ;
        RECT 171.100 335.140 196.500 362.000 ;
        RECT 197.700 335.140 223.100 362.000 ;
        RECT 224.300 335.140 249.700 362.000 ;
        RECT 250.900 335.140 276.300 362.000 ;
        RECT 277.500 335.140 302.900 362.000 ;
        RECT 304.100 335.140 329.500 362.000 ;
        RECT 330.700 335.140 356.100 362.000 ;
        RECT 357.300 335.140 382.700 362.000 ;
        RECT 383.900 335.140 409.300 362.000 ;
        RECT 410.500 335.140 435.900 362.000 ;
        RECT 437.100 335.140 462.500 362.000 ;
        RECT 91.300 307.080 116.700 333.940 ;
        RECT 117.900 307.080 143.300 333.940 ;
        RECT 144.500 307.080 169.900 333.940 ;
        RECT 171.100 307.080 196.500 333.940 ;
        RECT 197.700 307.080 223.100 333.940 ;
        RECT 224.300 307.080 249.700 333.940 ;
        RECT 250.900 307.080 276.300 333.940 ;
        RECT 277.500 307.080 302.900 333.940 ;
        RECT 304.100 307.080 329.500 333.940 ;
        RECT 330.700 307.080 356.100 333.940 ;
        RECT 357.300 307.080 382.700 333.940 ;
        RECT 383.900 307.080 409.300 333.940 ;
        RECT 410.500 307.080 435.900 333.940 ;
        RECT 437.100 307.080 462.500 333.940 ;
        RECT 91.300 279.020 116.700 305.880 ;
        RECT 117.900 279.020 143.300 305.880 ;
        RECT 144.500 279.020 169.900 305.880 ;
        RECT 171.100 279.020 196.500 305.880 ;
        RECT 197.700 279.020 223.100 305.880 ;
        RECT 224.300 279.020 249.700 305.880 ;
        RECT 250.900 279.020 276.300 305.880 ;
        RECT 277.500 279.020 302.900 305.880 ;
        RECT 304.100 279.020 329.500 305.880 ;
        RECT 330.700 279.020 356.100 305.880 ;
        RECT 357.300 279.020 382.700 305.880 ;
        RECT 383.900 279.020 409.300 305.880 ;
        RECT 410.500 279.020 435.900 305.880 ;
        RECT 437.100 279.020 462.500 305.880 ;
        RECT 91.300 250.960 116.700 277.820 ;
        RECT 117.900 250.960 143.300 277.820 ;
        RECT 144.500 250.960 169.900 277.820 ;
        RECT 171.100 250.960 196.500 277.820 ;
        RECT 197.700 250.960 223.100 277.820 ;
        RECT 224.300 250.960 249.700 277.820 ;
        RECT 250.900 250.960 276.300 277.820 ;
        RECT 277.500 250.960 302.900 277.820 ;
        RECT 304.100 250.960 329.500 277.820 ;
        RECT 330.700 250.960 356.100 277.820 ;
        RECT 357.300 250.960 382.700 277.820 ;
        RECT 383.900 250.960 409.300 277.820 ;
        RECT 410.500 250.960 435.900 277.820 ;
        RECT 437.100 250.960 462.500 277.820 ;
        RECT 91.300 222.900 116.700 249.760 ;
        RECT 117.900 222.900 143.300 249.760 ;
        RECT 144.500 222.900 169.900 249.760 ;
        RECT 171.100 222.900 196.500 249.760 ;
        RECT 197.700 222.900 223.100 249.760 ;
        RECT 224.300 222.900 249.700 249.760 ;
        RECT 250.900 222.900 276.300 249.760 ;
        RECT 277.500 222.900 302.900 249.760 ;
        RECT 304.100 222.900 329.500 249.760 ;
        RECT 330.700 222.900 356.100 249.760 ;
        RECT 357.300 222.900 382.700 249.760 ;
        RECT 383.900 222.900 409.300 249.760 ;
        RECT 410.500 222.900 435.900 249.760 ;
        RECT 437.100 222.900 462.500 249.760 ;
        RECT 91.300 194.840 116.700 221.700 ;
        RECT 117.900 194.840 143.300 221.700 ;
        RECT 144.500 194.840 169.900 221.700 ;
        RECT 171.100 194.840 196.500 221.700 ;
        RECT 197.700 194.840 223.100 221.700 ;
        RECT 224.300 194.840 249.700 221.700 ;
        RECT 250.900 194.840 276.300 221.700 ;
        RECT 277.500 194.840 302.900 221.700 ;
        RECT 304.100 194.840 329.500 221.700 ;
        RECT 330.700 194.840 356.100 221.700 ;
        RECT 357.300 194.840 382.700 221.700 ;
        RECT 383.900 194.840 409.300 221.700 ;
        RECT 410.500 194.840 435.900 221.700 ;
        RECT 437.100 194.840 462.500 221.700 ;
        RECT 91.300 166.780 116.700 193.640 ;
        RECT 117.900 166.780 143.300 193.640 ;
        RECT 144.500 166.780 169.900 193.640 ;
        RECT 171.100 166.780 196.500 193.640 ;
        RECT 197.700 166.780 223.100 193.640 ;
        RECT 224.300 166.780 249.700 193.640 ;
        RECT 250.900 166.780 276.300 193.640 ;
        RECT 277.500 166.780 302.900 193.640 ;
        RECT 304.100 166.780 329.500 193.640 ;
        RECT 330.700 166.780 356.100 193.640 ;
        RECT 357.300 166.780 382.700 193.640 ;
        RECT 383.900 166.780 409.300 193.640 ;
        RECT 410.500 166.780 435.900 193.640 ;
        RECT 437.100 166.780 462.500 193.640 ;
        RECT 1.585 132.435 11.985 144.295 ;
        RECT 13.185 132.435 23.585 144.295 ;
        RECT 24.785 132.435 35.185 144.295 ;
        RECT 36.385 132.435 46.785 144.295 ;
        RECT 47.985 132.435 58.385 144.295 ;
        RECT 59.585 132.435 69.985 144.295 ;
        RECT 71.185 132.435 81.585 144.295 ;
        RECT 91.300 138.720 116.700 165.580 ;
        RECT 117.900 138.720 143.300 165.580 ;
        RECT 144.500 138.720 169.900 165.580 ;
        RECT 171.100 138.720 196.500 165.580 ;
        RECT 197.700 138.720 223.100 165.580 ;
        RECT 224.300 138.720 249.700 165.580 ;
        RECT 250.900 138.720 276.300 165.580 ;
        RECT 277.500 138.720 302.900 165.580 ;
        RECT 304.100 138.720 329.500 165.580 ;
        RECT 330.700 138.720 356.100 165.580 ;
        RECT 357.300 138.720 382.700 165.580 ;
        RECT 383.900 138.720 409.300 165.580 ;
        RECT 410.500 138.720 435.900 165.580 ;
        RECT 437.100 138.720 462.500 165.580 ;
        RECT 1.585 119.375 11.985 131.235 ;
        RECT 13.185 119.375 23.585 131.235 ;
        RECT 24.785 119.375 35.185 131.235 ;
        RECT 36.385 119.375 46.785 131.235 ;
        RECT 47.985 119.375 58.385 131.235 ;
        RECT 59.585 119.375 69.985 131.235 ;
        RECT 71.185 119.375 81.585 131.235 ;
        RECT 1.585 106.315 11.985 118.175 ;
        RECT 13.185 106.315 23.585 118.175 ;
        RECT 24.785 106.315 35.185 118.175 ;
        RECT 36.385 106.315 46.785 118.175 ;
        RECT 47.985 106.315 58.385 118.175 ;
        RECT 59.585 106.315 69.985 118.175 ;
        RECT 71.185 106.315 81.585 118.175 ;
        RECT 91.300 110.660 116.700 137.520 ;
        RECT 117.900 110.660 143.300 137.520 ;
        RECT 144.500 110.660 169.900 137.520 ;
        RECT 171.100 110.660 196.500 137.520 ;
        RECT 197.700 110.660 223.100 137.520 ;
        RECT 224.300 110.660 249.700 137.520 ;
        RECT 250.900 110.660 276.300 137.520 ;
        RECT 277.500 110.660 302.900 137.520 ;
        RECT 304.100 110.660 329.500 137.520 ;
        RECT 330.700 110.660 356.100 137.520 ;
        RECT 357.300 110.660 382.700 137.520 ;
        RECT 383.900 110.660 409.300 137.520 ;
        RECT 410.500 110.660 435.900 137.520 ;
        RECT 437.100 110.660 462.500 137.520 ;
        RECT 1.585 93.255 11.985 105.115 ;
        RECT 13.185 93.255 23.585 105.115 ;
        RECT 24.785 93.255 35.185 105.115 ;
        RECT 36.385 93.255 46.785 105.115 ;
        RECT 47.985 93.255 58.385 105.115 ;
        RECT 59.585 93.255 69.985 105.115 ;
        RECT 71.185 93.255 81.585 105.115 ;
        RECT 1.585 80.195 11.985 92.055 ;
        RECT 13.185 80.195 23.585 92.055 ;
        RECT 24.785 80.195 35.185 92.055 ;
        RECT 36.385 80.195 46.785 92.055 ;
        RECT 47.985 80.195 58.385 92.055 ;
        RECT 59.585 80.195 69.985 92.055 ;
        RECT 71.185 80.195 81.585 92.055 ;
        RECT 1.585 67.135 11.985 78.995 ;
        RECT 13.185 67.135 23.585 78.995 ;
        RECT 24.785 67.135 35.185 78.995 ;
        RECT 36.385 67.135 46.785 78.995 ;
        RECT 47.985 67.135 58.385 78.995 ;
        RECT 59.585 67.135 69.985 78.995 ;
        RECT 71.185 67.135 81.585 78.995 ;
        RECT 1.585 54.075 11.985 65.935 ;
        RECT 13.185 54.075 23.585 65.935 ;
        RECT 24.785 54.075 35.185 65.935 ;
        RECT 36.385 54.075 46.785 65.935 ;
        RECT 47.985 54.075 58.385 65.935 ;
        RECT 59.585 54.075 69.985 65.935 ;
        RECT 71.185 54.075 81.585 65.935 ;
        RECT 84.745 56.750 86.410 84.195 ;
        RECT 91.300 82.600 116.700 109.460 ;
        RECT 117.900 82.600 143.300 109.460 ;
        RECT 144.500 82.600 169.900 109.460 ;
        RECT 171.100 82.600 196.500 109.460 ;
        RECT 197.700 82.600 223.100 109.460 ;
        RECT 224.300 82.600 249.700 109.460 ;
        RECT 250.900 82.600 276.300 109.460 ;
        RECT 277.500 82.600 302.900 109.460 ;
        RECT 304.100 82.600 329.500 109.460 ;
        RECT 330.700 82.600 356.100 109.460 ;
        RECT 357.300 82.600 382.700 109.460 ;
        RECT 383.900 82.600 409.300 109.460 ;
        RECT 410.500 82.600 435.900 109.460 ;
        RECT 437.100 82.600 462.500 109.460 ;
        RECT 91.300 54.540 116.700 81.400 ;
        RECT 117.900 54.540 143.300 81.400 ;
        RECT 144.500 54.540 169.900 81.400 ;
        RECT 171.100 54.540 196.500 81.400 ;
        RECT 197.700 54.540 223.100 81.400 ;
        RECT 224.300 54.540 249.700 81.400 ;
        RECT 250.900 54.540 276.300 81.400 ;
        RECT 277.500 54.540 302.900 81.400 ;
        RECT 304.100 54.540 329.500 81.400 ;
        RECT 330.700 54.540 356.100 81.400 ;
        RECT 357.300 54.540 382.700 81.400 ;
        RECT 383.900 54.540 409.300 81.400 ;
        RECT 410.500 54.540 435.900 81.400 ;
        RECT 437.100 54.540 462.500 81.400 ;
      LAYER met4 ;
        RECT 85.870 446.180 90.150 446.540 ;
        RECT 85.870 445.660 463.100 446.180 ;
        RECT 85.870 418.120 90.150 445.660 ;
        RECT 85.870 417.600 463.100 418.120 ;
        RECT 85.870 390.060 90.150 417.600 ;
        RECT 85.870 389.540 463.100 390.060 ;
        RECT 85.870 362.000 90.150 389.540 ;
        RECT 85.870 361.480 463.100 362.000 ;
        RECT 85.870 333.940 90.150 361.480 ;
        RECT 85.870 333.420 463.100 333.940 ;
        RECT 85.870 305.880 90.150 333.420 ;
        RECT 85.870 305.360 463.100 305.880 ;
        RECT 85.870 277.820 90.150 305.360 ;
        RECT 85.870 277.300 463.100 277.820 ;
        RECT 85.870 249.760 90.150 277.300 ;
        RECT 85.870 249.240 463.100 249.760 ;
        RECT 85.870 221.700 90.150 249.240 ;
        RECT 85.870 221.180 463.100 221.700 ;
        RECT 85.870 193.640 90.150 221.180 ;
        RECT 85.870 193.120 463.100 193.640 ;
        RECT 85.870 165.580 90.150 193.120 ;
        RECT 85.870 165.060 463.100 165.580 ;
        RECT 85.870 144.295 90.150 165.060 ;
        RECT 0.985 143.775 90.150 144.295 ;
        RECT 84.060 137.520 90.150 143.775 ;
        RECT 84.060 137.000 463.100 137.520 ;
        RECT 84.060 131.235 90.150 137.000 ;
        RECT 0.985 130.715 90.150 131.235 ;
        RECT 84.060 118.175 90.150 130.715 ;
        RECT 0.985 117.655 90.150 118.175 ;
        RECT 84.060 109.460 90.150 117.655 ;
        RECT 84.060 108.940 463.100 109.460 ;
        RECT 84.060 105.115 90.150 108.940 ;
        RECT 0.985 104.595 90.150 105.115 ;
        RECT 84.060 92.055 90.150 104.595 ;
        RECT 0.985 91.535 90.150 92.055 ;
        RECT 84.060 81.400 90.150 91.535 ;
        RECT 84.060 80.880 463.100 81.400 ;
        RECT 84.060 78.995 90.150 80.880 ;
        RECT 0.985 78.475 90.150 78.995 ;
        RECT 84.060 65.935 90.150 78.475 ;
        RECT 0.985 65.415 90.150 65.935 ;
        RECT 84.060 57.545 90.150 65.415 ;
        RECT 84.060 56.225 86.960 57.545 ;
    END
  END VSS
  OBS
      LAYER pwell ;
        RECT -63.385 598.110 -61.625 599.150 ;
        RECT -63.385 595.920 -61.625 597.450 ;
        RECT -53.620 596.725 -52.860 598.745 ;
        RECT -59.420 591.730 -58.660 593.750 ;
        RECT -52.085 593.190 -50.325 595.700 ;
        RECT -45.675 593.325 -43.915 594.365 ;
        RECT -45.675 591.695 -42.915 593.225 ;
        RECT -61.955 588.195 -60.195 590.705 ;
        RECT -52.475 588.815 -51.215 590.835 ;
        RECT -45.675 590.555 -42.915 591.595 ;
        RECT -45.675 589.440 -42.915 590.480 ;
        RECT -45.675 587.090 -43.915 588.130 ;
        RECT -63.230 579.770 -61.470 580.810 ;
        RECT -63.230 577.580 -61.470 579.110 ;
        RECT -53.465 578.385 -52.705 580.405 ;
        RECT -45.965 579.810 -44.205 580.850 ;
        RECT -45.965 577.620 -44.205 579.150 ;
        RECT -36.200 578.425 -35.440 580.445 ;
        RECT -59.265 573.390 -58.505 575.410 ;
        RECT -51.930 574.850 -50.170 577.360 ;
        RECT -42.000 573.430 -41.240 575.450 ;
        RECT -34.665 574.890 -32.905 577.400 ;
        RECT -61.800 569.855 -60.040 572.365 ;
        RECT -52.320 570.475 -51.060 572.495 ;
        RECT -44.535 569.895 -42.775 572.405 ;
        RECT -35.055 570.515 -33.795 572.535 ;
        RECT -63.575 551.290 -61.815 552.330 ;
        RECT -63.575 549.100 -61.815 550.630 ;
        RECT -53.810 549.905 -53.050 551.925 ;
        RECT -59.610 544.910 -58.850 546.930 ;
        RECT -52.275 546.370 -50.515 548.880 ;
        RECT -45.865 546.505 -44.105 547.545 ;
        RECT -45.865 544.875 -43.105 546.405 ;
        RECT -62.145 541.375 -60.385 543.885 ;
        RECT -52.665 541.995 -51.405 544.015 ;
        RECT -45.865 543.735 -43.105 544.775 ;
        RECT -45.865 542.620 -43.105 543.660 ;
        RECT -45.865 540.270 -44.105 541.310 ;
        RECT -63.420 532.950 -61.660 533.990 ;
        RECT -63.420 530.760 -61.660 532.290 ;
        RECT -53.655 531.565 -52.895 533.585 ;
        RECT -46.155 532.990 -44.395 534.030 ;
        RECT -46.155 530.800 -44.395 532.330 ;
        RECT -36.390 531.605 -35.630 533.625 ;
        RECT -59.455 526.570 -58.695 528.590 ;
        RECT -52.120 528.030 -50.360 530.540 ;
        RECT -42.190 526.610 -41.430 528.630 ;
        RECT -34.855 528.070 -33.095 530.580 ;
        RECT -61.990 523.035 -60.230 525.545 ;
        RECT -52.510 523.655 -51.250 525.675 ;
        RECT -44.725 523.075 -42.965 525.585 ;
        RECT -35.245 523.695 -33.985 525.715 ;
        RECT -63.660 505.525 -61.900 506.565 ;
        RECT -63.660 503.335 -61.900 504.865 ;
        RECT -53.895 504.140 -53.135 506.160 ;
        RECT -59.695 499.145 -58.935 501.165 ;
        RECT -52.360 500.605 -50.600 503.115 ;
        RECT -45.950 500.740 -44.190 501.780 ;
        RECT -45.950 499.110 -43.190 500.640 ;
        RECT -62.230 495.610 -60.470 498.120 ;
        RECT -52.750 496.230 -51.490 498.250 ;
        RECT -45.950 497.970 -43.190 499.010 ;
        RECT -45.950 496.855 -43.190 497.895 ;
        RECT -45.950 494.505 -44.190 495.545 ;
        RECT -63.505 487.185 -61.745 488.225 ;
        RECT -63.505 484.995 -61.745 486.525 ;
        RECT -53.740 485.800 -52.980 487.820 ;
        RECT -46.240 487.225 -44.480 488.265 ;
        RECT -46.240 485.035 -44.480 486.565 ;
        RECT -36.475 485.840 -35.715 487.860 ;
        RECT -59.540 480.805 -58.780 482.825 ;
        RECT -52.205 482.265 -50.445 484.775 ;
        RECT -42.275 480.845 -41.515 482.865 ;
        RECT -34.940 482.305 -33.180 484.815 ;
        RECT -62.075 477.270 -60.315 479.780 ;
        RECT -52.595 477.890 -51.335 479.910 ;
        RECT -44.810 477.310 -43.050 479.820 ;
        RECT -35.330 477.930 -34.070 479.950 ;
        RECT -63.990 461.755 -62.230 462.795 ;
        RECT -63.990 459.565 -62.230 461.095 ;
        RECT -54.225 460.370 -53.465 462.390 ;
        RECT -60.025 455.375 -59.265 457.395 ;
        RECT -52.690 456.835 -50.930 459.345 ;
        RECT -46.280 456.970 -44.520 458.010 ;
        RECT -46.280 455.340 -43.520 456.870 ;
        RECT -62.560 451.840 -60.800 454.350 ;
        RECT -53.080 452.460 -51.820 454.480 ;
        RECT -46.280 454.200 -43.520 455.240 ;
        RECT -46.280 453.085 -43.520 454.125 ;
        RECT -46.280 450.735 -44.520 451.775 ;
        RECT -63.835 443.415 -62.075 444.455 ;
        RECT -63.835 441.225 -62.075 442.755 ;
        RECT -54.070 442.030 -53.310 444.050 ;
        RECT -46.570 443.455 -44.810 444.495 ;
        RECT -46.570 441.265 -44.810 442.795 ;
        RECT -36.805 442.070 -36.045 444.090 ;
        RECT -59.870 437.035 -59.110 439.055 ;
        RECT -52.535 438.495 -50.775 441.005 ;
        RECT -42.605 437.075 -41.845 439.095 ;
        RECT -35.270 438.535 -33.510 441.045 ;
        RECT -62.405 433.500 -60.645 436.010 ;
        RECT -52.925 434.120 -51.665 436.140 ;
        RECT -45.140 433.540 -43.380 436.050 ;
        RECT -35.660 434.160 -34.400 436.180 ;
        RECT -64.160 415.765 -62.400 416.805 ;
        RECT -64.160 413.575 -62.400 415.105 ;
        RECT -54.395 414.380 -53.635 416.400 ;
        RECT -60.195 409.385 -59.435 411.405 ;
        RECT -52.860 410.845 -51.100 413.355 ;
        RECT -46.450 410.980 -44.690 412.020 ;
        RECT -46.450 409.350 -43.690 410.880 ;
        RECT -62.730 405.850 -60.970 408.360 ;
        RECT -53.250 406.470 -51.990 408.490 ;
        RECT -46.450 408.210 -43.690 409.250 ;
        RECT -46.450 407.095 -43.690 408.135 ;
        RECT -46.450 404.745 -44.690 405.785 ;
        RECT -64.005 397.425 -62.245 398.465 ;
        RECT -64.005 395.235 -62.245 396.765 ;
        RECT -54.240 396.040 -53.480 398.060 ;
        RECT -46.740 397.465 -44.980 398.505 ;
        RECT -46.740 395.275 -44.980 396.805 ;
        RECT -36.975 396.080 -36.215 398.100 ;
        RECT -60.040 391.045 -59.280 393.065 ;
        RECT -52.705 392.505 -50.945 395.015 ;
        RECT -42.775 391.085 -42.015 393.105 ;
        RECT -35.440 392.545 -33.680 395.055 ;
        RECT -62.575 387.510 -60.815 390.020 ;
        RECT -53.095 388.130 -51.835 390.150 ;
        RECT -45.310 387.550 -43.550 390.060 ;
        RECT -35.830 388.170 -34.570 390.190 ;
        RECT -63.965 371.450 -62.205 372.490 ;
        RECT -63.965 369.260 -62.205 370.790 ;
        RECT -54.200 370.065 -53.440 372.085 ;
        RECT -60.000 365.070 -59.240 367.090 ;
        RECT -52.665 366.530 -50.905 369.040 ;
        RECT -46.255 366.665 -44.495 367.705 ;
        RECT -46.255 365.035 -43.495 366.565 ;
        RECT -62.535 361.535 -60.775 364.045 ;
        RECT -53.055 362.155 -51.795 364.175 ;
        RECT -46.255 363.895 -43.495 364.935 ;
        RECT -46.255 362.780 -43.495 363.820 ;
        RECT -46.255 360.430 -44.495 361.470 ;
        RECT -63.810 353.110 -62.050 354.150 ;
        RECT -63.810 350.920 -62.050 352.450 ;
        RECT -54.045 351.725 -53.285 353.745 ;
        RECT -46.545 353.150 -44.785 354.190 ;
        RECT -46.545 350.960 -44.785 352.490 ;
        RECT -36.780 351.765 -36.020 353.785 ;
        RECT -59.845 346.730 -59.085 348.750 ;
        RECT -52.510 348.190 -50.750 350.700 ;
        RECT -42.580 346.770 -41.820 348.790 ;
        RECT -35.245 348.230 -33.485 350.740 ;
        RECT -62.380 343.195 -60.620 345.705 ;
        RECT -52.900 343.815 -51.640 345.835 ;
        RECT -45.115 343.235 -43.355 345.745 ;
        RECT -35.635 343.855 -34.375 345.875 ;
        RECT -63.910 329.250 -62.150 330.290 ;
        RECT -63.910 327.060 -62.150 328.590 ;
        RECT -54.145 327.865 -53.385 329.885 ;
        RECT -59.945 322.870 -59.185 324.890 ;
        RECT -52.610 324.330 -50.850 326.840 ;
        RECT -46.200 324.465 -44.440 325.505 ;
        RECT -46.200 322.835 -43.440 324.365 ;
        RECT -62.480 319.335 -60.720 321.845 ;
        RECT -53.000 319.955 -51.740 321.975 ;
        RECT -46.200 321.695 -43.440 322.735 ;
        RECT -46.200 320.580 -43.440 321.620 ;
        RECT -46.200 318.230 -44.440 319.270 ;
        RECT -63.755 310.910 -61.995 311.950 ;
        RECT -63.755 308.720 -61.995 310.250 ;
        RECT -53.990 309.525 -53.230 311.545 ;
        RECT -46.490 310.950 -44.730 311.990 ;
        RECT -46.490 308.760 -44.730 310.290 ;
        RECT -36.725 309.565 -35.965 311.585 ;
        RECT -59.790 304.530 -59.030 306.550 ;
        RECT -52.455 305.990 -50.695 308.500 ;
        RECT -42.525 304.570 -41.765 306.590 ;
        RECT -35.190 306.030 -33.430 308.540 ;
        RECT -62.325 300.995 -60.565 303.505 ;
        RECT -52.845 301.615 -51.585 303.635 ;
        RECT -45.060 301.035 -43.300 303.545 ;
        RECT -35.580 301.655 -34.320 303.675 ;
        RECT -52.070 288.250 -48.310 289.290 ;
        RECT -52.070 286.250 -48.310 287.290 ;
        RECT -43.685 286.500 -42.925 289.500 ;
        RECT -40.395 286.500 -39.635 289.500 ;
        RECT -52.070 283.250 -48.310 284.290 ;
        RECT -52.070 281.250 -48.310 282.290 ;
        RECT -43.435 281.330 -42.675 285.310 ;
        RECT -40.395 282.315 -39.635 285.315 ;
        RECT -52.070 278.250 -48.310 279.290 ;
        RECT -43.685 277.785 -42.925 280.785 ;
        RECT -40.645 277.790 -39.885 281.770 ;
        RECT -52.070 276.250 -48.310 277.290 ;
        RECT -54.950 271.850 -54.190 274.850 ;
        RECT -52.615 273.150 -51.355 274.190 ;
        RECT -52.615 272.100 -51.355 273.140 ;
        RECT -43.685 273.000 -42.925 276.000 ;
        RECT -40.395 273.000 -39.635 276.000 ;
        RECT -53.345 268.205 -52.085 269.245 ;
        RECT -43.435 267.830 -42.675 271.810 ;
        RECT -40.395 268.815 -39.635 271.815 ;
        RECT -53.845 265.650 -52.085 267.180 ;
        RECT -53.845 264.105 -52.085 265.635 ;
        RECT -43.685 264.285 -42.925 267.285 ;
        RECT -40.645 264.290 -39.885 268.270 ;
        RECT -53.850 262.555 -52.090 264.085 ;
        RECT -53.255 258.465 -51.995 259.995 ;
        RECT -43.685 259.875 -42.925 262.875 ;
        RECT -53.255 253.735 -51.995 255.265 ;
        RECT -40.165 253.760 -38.905 255.780 ;
        RECT -66.465 245.860 -65.705 248.860 ;
        RECT -63.175 245.860 -62.415 248.860 ;
        RECT -66.465 241.675 -65.705 244.675 ;
        RECT -66.215 237.150 -65.455 241.130 ;
        RECT -63.425 240.690 -62.665 244.670 ;
        RECT -63.175 237.145 -62.415 240.145 ;
        RECT -66.465 232.360 -65.705 235.360 ;
        RECT -63.175 232.360 -62.415 235.360 ;
        RECT -66.465 228.175 -65.705 231.175 ;
        RECT -66.215 223.650 -65.455 227.630 ;
        RECT -63.425 227.190 -62.665 231.170 ;
        RECT -63.175 223.645 -62.415 226.645 ;
        RECT -63.175 219.235 -62.415 222.235 ;
        RECT -66.150 202.595 -64.890 203.635 ;
        RECT -54.895 202.645 -53.635 203.685 ;
        RECT -40.775 202.645 -39.515 203.685 ;
        RECT -29.520 202.595 -28.260 203.635 ;
        RECT -66.150 201.050 -64.890 202.090 ;
        RECT -54.895 201.100 -53.635 202.140 ;
        RECT -40.775 201.100 -39.515 202.140 ;
        RECT -29.520 201.050 -28.260 202.090 ;
        RECT -66.150 199.500 -64.890 200.540 ;
        RECT -54.895 199.550 -53.635 200.590 ;
        RECT -40.775 199.550 -39.515 200.590 ;
        RECT -29.520 199.500 -28.260 200.540 ;
        RECT -66.150 198.030 -64.890 199.070 ;
        RECT -54.895 198.080 -53.635 199.120 ;
        RECT -40.775 198.080 -39.515 199.120 ;
        RECT -29.520 198.030 -28.260 199.070 ;
        RECT -66.150 196.220 -64.890 197.260 ;
        RECT -54.895 196.270 -53.635 197.310 ;
        RECT -40.775 196.270 -39.515 197.310 ;
        RECT -29.520 196.220 -28.260 197.260 ;
        RECT -66.150 194.150 -64.890 195.190 ;
        RECT -54.895 194.200 -53.635 195.240 ;
        RECT -40.775 194.200 -39.515 195.240 ;
        RECT -29.520 194.150 -28.260 195.190 ;
        RECT -54.945 191.295 -53.185 192.825 ;
        RECT -41.225 191.295 -39.465 192.825 ;
        RECT -54.940 189.745 -53.180 191.275 ;
        RECT -41.230 189.745 -39.470 191.275 ;
        RECT -66.150 187.595 -64.890 188.635 ;
        RECT -54.940 188.200 -53.180 189.730 ;
        RECT -41.230 188.200 -39.470 189.730 ;
        RECT -29.520 187.595 -28.260 188.635 ;
        RECT -66.150 186.050 -64.890 187.090 ;
        RECT -54.440 186.135 -53.180 187.175 ;
        RECT -41.230 186.135 -39.970 187.175 ;
        RECT -29.520 186.050 -28.260 187.090 ;
        RECT -66.150 184.500 -64.890 185.540 ;
        RECT -29.520 184.500 -28.260 185.540 ;
        RECT -66.150 183.030 -64.890 184.070 ;
        RECT -66.150 181.220 -64.890 182.260 ;
        RECT -55.170 181.550 -53.410 184.060 ;
        RECT -41.000 181.550 -39.240 184.060 ;
        RECT -29.520 183.030 -28.260 184.070 ;
        RECT -29.520 181.220 -28.260 182.260 ;
        RECT -66.150 179.150 -64.890 180.190 ;
        RECT -56.705 178.505 -55.945 180.525 ;
        RECT -38.465 178.505 -37.705 180.525 ;
        RECT -29.520 179.150 -28.260 180.190 ;
        RECT -66.150 175.095 -64.890 176.135 ;
        RECT -66.150 173.550 -64.890 174.590 ;
        RECT -55.180 173.525 -53.420 176.035 ;
        RECT -40.990 173.525 -39.230 176.035 ;
        RECT -29.520 175.095 -28.260 176.135 ;
        RECT -29.520 173.550 -28.260 174.590 ;
        RECT -66.150 172.000 -64.890 173.040 ;
        RECT -66.150 170.530 -64.890 171.570 ;
        RECT -56.715 170.480 -55.955 172.500 ;
        RECT -38.455 170.480 -37.695 172.500 ;
        RECT -29.520 172.000 -28.260 173.040 ;
        RECT -29.520 170.530 -28.260 171.570 ;
        RECT -66.150 168.720 -64.890 169.760 ;
        RECT -29.520 168.720 -28.260 169.760 ;
        RECT -66.150 166.650 -64.890 167.690 ;
        RECT -54.900 166.485 -53.140 168.015 ;
        RECT -41.270 166.485 -39.510 168.015 ;
        RECT -29.520 166.650 -28.260 167.690 ;
        RECT -54.895 164.935 -53.135 166.465 ;
        RECT -41.275 164.935 -39.515 166.465 ;
        RECT -66.150 162.595 -64.890 163.635 ;
        RECT -54.895 163.390 -53.135 164.920 ;
        RECT -41.275 163.390 -39.515 164.920 ;
        RECT -29.520 162.595 -28.260 163.635 ;
        RECT -66.150 161.050 -64.890 162.090 ;
        RECT -54.395 161.325 -53.135 162.365 ;
        RECT -41.275 161.325 -40.015 162.365 ;
        RECT -29.520 161.050 -28.260 162.090 ;
        RECT -66.150 159.500 -64.890 160.540 ;
        RECT -66.150 158.030 -64.890 159.070 ;
        RECT -66.150 156.220 -64.890 157.260 ;
        RECT -56.120 156.675 -55.360 159.675 ;
        RECT -39.050 156.675 -38.290 159.675 ;
        RECT -29.520 159.500 -28.260 160.540 ;
        RECT -29.520 158.030 -28.260 159.070 ;
        RECT -29.520 156.220 -28.260 157.260 ;
        RECT -66.150 154.150 -64.890 155.190 ;
        RECT -56.120 152.265 -55.360 155.265 ;
        RECT -66.150 150.095 -64.890 151.135 ;
        RECT -66.150 148.550 -64.890 149.590 ;
        RECT -66.150 147.000 -64.890 148.040 ;
        RECT -55.870 147.740 -55.110 151.720 ;
        RECT -53.080 151.280 -52.320 155.260 ;
        RECT -42.090 151.280 -41.330 155.260 ;
        RECT -39.050 152.265 -38.290 155.265 ;
        RECT -29.520 154.150 -28.260 155.190 ;
        RECT -52.830 147.735 -52.070 150.735 ;
        RECT -42.340 147.735 -41.580 150.735 ;
        RECT -39.300 147.740 -38.540 151.720 ;
        RECT -29.520 150.095 -28.260 151.135 ;
        RECT -29.520 148.550 -28.260 149.590 ;
        RECT -29.520 147.000 -28.260 148.040 ;
        RECT -66.150 145.530 -64.890 146.570 ;
        RECT -66.150 143.720 -64.890 144.760 ;
        RECT -56.120 143.550 -55.360 146.550 ;
        RECT -52.830 143.550 -52.070 146.550 ;
        RECT -42.340 143.550 -41.580 146.550 ;
        RECT -39.050 143.550 -38.290 146.550 ;
        RECT -29.520 145.530 -28.260 146.570 ;
        RECT -29.520 143.720 -28.260 144.760 ;
        RECT -66.150 141.650 -64.890 142.690 ;
        RECT -56.120 138.765 -55.360 141.765 ;
        RECT -66.150 137.595 -64.890 138.635 ;
        RECT -66.150 136.050 -64.890 137.090 ;
        RECT -66.150 134.500 -64.890 135.540 ;
        RECT -55.870 134.240 -55.110 138.220 ;
        RECT -53.080 137.780 -52.320 141.760 ;
        RECT -42.090 137.780 -41.330 141.760 ;
        RECT -39.050 138.765 -38.290 141.765 ;
        RECT -29.520 141.650 -28.260 142.690 ;
        RECT -52.830 134.235 -52.070 137.235 ;
        RECT -42.340 134.235 -41.580 137.235 ;
        RECT -39.300 134.240 -38.540 138.220 ;
        RECT -29.520 137.595 -28.260 138.635 ;
        RECT -29.520 136.050 -28.260 137.090 ;
        RECT -29.520 134.500 -28.260 135.540 ;
        RECT -66.150 133.030 -64.890 134.070 ;
        RECT -66.150 131.220 -64.890 132.260 ;
        RECT -66.150 129.150 -64.890 130.190 ;
        RECT -56.120 130.050 -55.360 133.050 ;
        RECT -52.830 130.050 -52.070 133.050 ;
        RECT -42.340 130.050 -41.580 133.050 ;
        RECT -39.050 130.050 -38.290 133.050 ;
        RECT -31.235 131.335 -30.475 134.335 ;
        RECT -29.520 133.030 -28.260 134.070 ;
        RECT -29.520 131.220 -28.260 132.260 ;
        RECT -29.520 129.150 -28.260 130.190 ;
        RECT -55.240 124.250 -53.480 125.780 ;
        RECT -30.570 124.115 -28.810 125.645 ;
        RECT -55.240 122.550 -53.480 123.590 ;
        RECT -30.570 122.415 -28.810 123.455 ;
        RECT -54.785 117.305 -54.025 120.305 ;
        RECT -30.150 117.305 -29.390 120.305 ;
        RECT -54.785 112.895 -54.025 115.895 ;
        RECT -54.535 108.370 -53.775 112.350 ;
        RECT -51.745 111.910 -50.985 115.890 ;
        RECT -30.150 112.895 -29.390 115.895 ;
        RECT -51.495 108.365 -50.735 111.365 ;
        RECT -29.900 108.370 -29.140 112.350 ;
        RECT -27.110 111.910 -26.350 115.890 ;
        RECT -26.860 108.365 -26.100 111.365 ;
        RECT -54.785 104.180 -54.025 107.180 ;
        RECT -51.495 104.180 -50.735 107.180 ;
        RECT -44.845 104.335 -44.085 106.355 ;
        RECT -36.080 105.720 -34.320 106.760 ;
        RECT -36.080 103.530 -34.320 105.060 ;
        RECT -30.150 104.180 -29.390 107.180 ;
        RECT -26.860 104.180 -26.100 107.180 ;
        RECT -54.785 99.395 -54.025 102.395 ;
        RECT -54.535 94.870 -53.775 98.850 ;
        RECT -51.745 98.410 -50.985 102.390 ;
        RECT -47.380 100.800 -45.620 103.310 ;
        RECT -39.045 99.340 -38.285 101.360 ;
        RECT -30.150 99.395 -29.390 102.395 ;
        RECT -51.495 94.865 -50.735 97.865 ;
        RECT -46.490 96.425 -45.230 98.445 ;
        RECT -37.510 95.805 -35.750 98.315 ;
        RECT -29.900 94.870 -29.140 98.850 ;
        RECT -27.110 98.410 -26.350 102.390 ;
        RECT -26.860 94.865 -26.100 97.865 ;
        RECT -54.785 90.680 -54.025 93.680 ;
        RECT -51.495 90.680 -50.735 93.680 ;
        RECT -30.150 90.680 -29.390 93.680 ;
        RECT -26.860 90.680 -26.100 93.680 ;
        RECT -64.965 79.390 -64.205 81.410 ;
        RECT -56.200 80.775 -54.440 81.815 ;
        RECT -56.200 78.585 -54.440 80.115 ;
        RECT -39.965 79.390 -39.205 81.410 ;
        RECT -31.200 80.775 -29.440 81.815 ;
        RECT -31.200 78.585 -29.440 80.115 ;
        RECT -67.500 75.855 -65.740 78.365 ;
        RECT -59.165 74.395 -58.405 76.415 ;
        RECT -42.500 75.855 -40.740 78.365 ;
        RECT -34.165 74.395 -33.405 76.415 ;
        RECT -66.610 71.480 -65.350 73.500 ;
        RECT -57.630 70.860 -55.870 73.370 ;
        RECT -41.610 71.480 -40.350 73.500 ;
        RECT -32.630 70.860 -30.870 73.370 ;
        RECT -42.615 67.485 -41.355 68.525 ;
        RECT -58.630 64.340 -57.370 65.870 ;
        RECT -42.615 64.930 -40.855 66.460 ;
        RECT -30.655 66.215 -29.895 68.235 ;
        RECT -42.615 63.385 -40.855 64.915 ;
        RECT -42.610 61.835 -40.850 63.365 ;
        RECT -33.190 62.680 -31.430 65.190 ;
        RECT -58.625 59.815 -57.365 61.345 ;
        RECT -66.575 57.260 -64.815 58.790 ;
        RECT -66.570 55.710 -64.810 57.240 ;
        RECT -40.200 56.505 -39.440 58.525 ;
        RECT -32.935 58.335 -31.675 59.375 ;
        RECT -66.570 54.165 -64.810 55.695 ;
        RECT -60.340 53.785 -59.080 55.805 ;
        RECT -32.935 55.780 -31.175 57.310 ;
        RECT -66.070 52.100 -64.810 53.140 ;
        RECT -42.735 52.970 -40.975 55.480 ;
        RECT -32.935 54.235 -31.175 55.765 ;
        RECT -32.930 52.685 -31.170 54.215 ;
        RECT 79.960 45.340 81.220 51.050 ;
        RECT 81.960 45.340 83.220 51.050 ;
        RECT 83.960 45.340 85.220 51.050 ;
        RECT 80.035 44.080 80.715 45.220 ;
        RECT 40.710 28.085 58.420 32.345 ;
        RECT 40.710 23.085 62.710 27.345 ;
        RECT 98.780 14.360 101.780 15.120 ;
        RECT 103.030 14.360 106.030 15.120 ;
        RECT 106.260 14.030 110.730 15.290 ;
        RECT 103.030 12.285 106.030 13.045 ;
        RECT 106.260 12.115 110.730 13.375 ;
        RECT 2.935 9.875 3.925 10.555 ;
        RECT 4.165 9.820 7.365 10.680 ;
        RECT 7.385 9.845 8.815 10.705 ;
        RECT 8.955 9.880 11.865 10.740 ;
        RECT 12.310 9.875 13.300 10.555 ;
        RECT 13.855 9.875 14.845 10.555 ;
        RECT 151.460 10.350 158.330 12.610 ;
        RECT 175.135 10.460 182.005 12.720 ;
        RECT 183.740 10.245 190.610 12.505 ;
        RECT 195.740 12.145 198.740 12.905 ;
        RECT 200.150 12.145 203.150 12.905 ;
        RECT 203.695 11.895 207.675 12.655 ;
        RECT 208.865 12.145 211.865 12.905 ;
        RECT 213.650 12.145 216.650 12.905 ;
        RECT 217.195 11.895 221.175 12.655 ;
        RECT 222.365 12.145 225.365 12.905 ;
        RECT -21.110 7.265 -20.410 7.740 ;
        RECT -18.110 7.655 -15.110 8.415 ;
        RECT -13.860 7.655 -10.860 8.415 ;
        RECT -18.095 7.040 -15.165 7.640 ;
        RECT -13.845 7.040 -10.915 7.640 ;
        RECT -10.630 7.325 -6.160 8.585 ;
        RECT 22.385 8.535 25.385 9.295 ;
        RECT 26.635 8.535 29.635 9.295 ;
        RECT 29.865 8.205 34.335 9.465 ;
        RECT 200.155 9.105 204.135 9.865 ;
        RECT 204.680 8.855 207.680 9.615 ;
        RECT 208.865 8.855 211.865 9.615 ;
        RECT 213.655 9.105 217.635 9.865 ;
        RECT 218.180 8.855 221.180 9.615 ;
        RECT 222.365 8.855 225.365 9.615 ;
        RECT 227.705 9.305 230.705 10.065 ;
        RECT 255.750 9.000 291.700 11.260 ;
        RECT -13.845 6.355 -10.915 6.955 ;
        RECT -66.745 3.705 -30.795 5.965 ;
        RECT -13.860 5.580 -10.860 6.340 ;
        RECT -10.630 5.410 -6.160 6.670 ;
        RECT 26.635 6.460 29.635 7.220 ;
        RECT 29.865 6.290 34.335 7.550 ;
        RECT 39.360 5.115 75.310 7.375 ;
        RECT 138.890 4.575 140.230 5.835 ;
        RECT 140.290 4.565 144.000 5.825 ;
        RECT 144.040 4.565 145.380 5.825 ;
        RECT 145.420 4.555 146.760 5.815 ;
        RECT 163.165 4.540 164.505 5.800 ;
        RECT 164.565 4.530 168.275 5.790 ;
        RECT 168.315 4.530 169.655 5.790 ;
        RECT 169.695 4.520 171.035 5.780 ;
        RECT 2.935 3.755 3.925 4.435 ;
        RECT 4.165 3.630 7.365 4.490 ;
        RECT 7.385 3.605 8.815 4.465 ;
        RECT 8.955 3.570 11.865 4.430 ;
        RECT 12.310 3.755 13.300 4.435 ;
        RECT 13.855 3.755 14.845 4.435 ;
        RECT -66.880 2.655 -30.615 3.545 ;
        RECT 138.890 2.315 140.230 3.575 ;
        RECT 140.290 2.315 144.000 3.575 ;
        RECT 144.040 2.315 145.380 3.575 ;
        RECT 145.415 2.315 146.755 3.575 ;
        RECT 163.165 2.280 164.505 3.540 ;
        RECT 164.565 2.280 168.275 3.540 ;
        RECT 168.315 2.280 169.655 3.540 ;
        RECT 169.690 2.280 171.030 3.540 ;
        RECT 137.495 -0.245 138.835 1.015 ;
        RECT 138.855 -0.235 147.305 1.025 ;
        RECT 147.340 -0.235 148.680 1.025 ;
        RECT 151.460 -1.210 158.330 1.050 ;
        RECT 161.770 -0.280 163.110 0.980 ;
        RECT 163.130 -0.270 171.580 0.990 ;
        RECT 171.615 -0.270 172.955 0.990 ;
        RECT 175.135 -1.095 182.005 1.165 ;
        RECT 183.740 -0.880 190.610 1.380 ;
        RECT 99.640 -2.390 102.640 -1.630 ;
        RECT 103.890 -2.390 106.890 -1.630 ;
        RECT 107.120 -2.720 111.590 -1.460 ;
        RECT -25.450 -4.205 -22.450 -3.445 ;
        RECT -21.200 -4.205 -18.200 -3.445 ;
        RECT -25.435 -4.820 -22.505 -4.220 ;
        RECT -21.185 -4.820 -18.255 -4.220 ;
        RECT -17.970 -4.535 -13.500 -3.275 ;
        RECT -21.185 -5.505 -18.255 -4.905 ;
        RECT 22.460 -4.915 25.460 -4.155 ;
        RECT 26.710 -4.915 29.710 -4.155 ;
        RECT -21.200 -6.280 -18.200 -5.520 ;
        RECT -17.970 -6.450 -13.500 -5.190 ;
        RECT 29.940 -5.245 34.410 -3.985 ;
        RECT 103.890 -4.465 106.890 -3.705 ;
        RECT 107.120 -4.635 111.590 -3.375 ;
        RECT 254.735 -5.555 290.685 -3.295 ;
        RECT 26.710 -6.990 29.710 -6.230 ;
        RECT 29.940 -7.160 34.410 -5.900 ;
        RECT 39.155 -8.665 75.105 -6.405 ;
        RECT 311.775 -16.720 314.775 -15.960 ;
        RECT 316.025 -16.720 319.025 -15.960 ;
        RECT 319.255 -17.050 323.725 -15.790 ;
        RECT 254.735 -20.790 290.685 -18.530 ;
        RECT 316.025 -18.795 319.025 -18.035 ;
        RECT 319.255 -18.965 323.725 -17.705 ;
        RECT -75.080 -76.350 -38.815 -75.460 ;
        RECT -74.945 -78.770 -38.995 -76.510 ;
        RECT -75.885 -94.515 -72.885 -93.755 ;
        RECT -71.700 -94.515 -68.700 -93.755 ;
        RECT -75.870 -95.130 -72.940 -94.530 ;
        RECT -71.685 -95.130 -68.755 -94.530 ;
        RECT -68.155 -94.765 -64.175 -94.005 ;
        RECT -62.385 -94.515 -59.385 -93.755 ;
        RECT -58.200 -94.515 -55.200 -93.755 ;
        RECT -62.370 -95.130 -59.440 -94.530 ;
        RECT -58.185 -95.130 -55.255 -94.530 ;
        RECT -54.655 -94.765 -50.675 -94.005 ;
        RECT -88.365 -96.810 -84.370 -96.140 ;
        RECT -75.830 -97.030 -72.900 -96.430 ;
        RECT -100.350 -98.310 -98.330 -97.550 ;
        RECT -113.880 -100.585 -112.350 -98.825 ;
        RECT -112.330 -100.590 -110.800 -98.830 ;
        RECT -110.785 -100.590 -109.255 -98.830 ;
        RECT -100.710 -98.975 -97.805 -98.320 ;
        RECT -95.745 -98.505 -93.240 -97.940 ;
        RECT -108.230 -100.590 -107.190 -99.330 ;
        RECT -103.885 -100.845 -101.375 -99.085 ;
        RECT -95.705 -100.285 -93.195 -98.525 ;
        RECT -87.980 -98.855 -86.450 -97.095 ;
        RECT -85.790 -98.855 -84.750 -97.095 ;
        RECT -75.885 -97.805 -72.885 -97.045 ;
        RECT -71.695 -97.555 -67.715 -96.795 ;
        RECT -67.115 -97.030 -64.185 -96.430 ;
        RECT -62.330 -97.030 -59.400 -96.430 ;
        RECT -67.170 -97.805 -64.170 -97.045 ;
        RECT -62.385 -97.805 -59.385 -97.045 ;
        RECT -58.195 -97.555 -54.215 -96.795 ;
        RECT -53.615 -97.030 -50.685 -96.430 ;
        RECT -49.205 -97.030 -46.275 -96.430 ;
        RECT -53.670 -97.805 -50.670 -97.045 ;
        RECT -49.260 -97.805 -46.260 -97.045 ;
        RECT -44.150 -98.225 -43.110 -96.465 ;
        RECT -42.450 -98.225 -40.920 -96.465 ;
        RECT -37.415 -97.175 -36.375 -95.915 ;
        RECT -35.345 -97.175 -34.305 -95.915 ;
        RECT -33.535 -97.175 -32.495 -95.915 ;
        RECT -32.065 -97.175 -31.025 -95.915 ;
        RECT -30.515 -97.175 -29.475 -95.915 ;
        RECT -28.970 -97.175 -27.930 -95.915 ;
        RECT -24.915 -97.175 -23.875 -95.915 ;
        RECT -22.845 -97.175 -21.805 -95.915 ;
        RECT -21.035 -97.175 -19.995 -95.915 ;
        RECT -19.565 -97.175 -18.525 -95.915 ;
        RECT -18.015 -97.175 -16.975 -95.915 ;
        RECT -16.470 -97.175 -15.430 -95.915 ;
        RECT -12.415 -97.175 -11.375 -95.915 ;
        RECT -10.345 -97.175 -9.305 -95.915 ;
        RECT -8.535 -97.175 -7.495 -95.915 ;
        RECT -7.065 -97.175 -6.025 -95.915 ;
        RECT -5.515 -97.175 -4.475 -95.915 ;
        RECT -3.970 -97.175 -2.930 -95.915 ;
        RECT 0.085 -97.175 1.125 -95.915 ;
        RECT 2.155 -97.175 3.195 -95.915 ;
        RECT 3.965 -97.175 5.005 -95.915 ;
        RECT 5.435 -97.175 6.475 -95.915 ;
        RECT 6.985 -97.175 8.025 -95.915 ;
        RECT 8.530 -97.175 9.570 -95.915 ;
        RECT 12.585 -97.175 13.625 -95.915 ;
        RECT 14.655 -97.175 15.695 -95.915 ;
        RECT 16.465 -97.175 17.505 -95.915 ;
        RECT 17.935 -97.175 18.975 -95.915 ;
        RECT 19.485 -97.175 20.525 -95.915 ;
        RECT 21.030 -97.175 22.070 -95.915 ;
        RECT 27.585 -97.175 28.625 -95.915 ;
        RECT 29.655 -97.175 30.695 -95.915 ;
        RECT 31.465 -97.175 32.505 -95.915 ;
        RECT 32.935 -97.175 33.975 -95.915 ;
        RECT 34.485 -97.175 35.525 -95.915 ;
        RECT 36.030 -97.175 37.070 -95.915 ;
        RECT -35.215 -98.115 -32.285 -97.515 ;
        RECT -31.370 -98.060 -27.950 -97.320 ;
        RECT -18.870 -98.060 -15.450 -97.320 ;
        RECT -6.370 -98.060 -2.950 -97.320 ;
        RECT 6.130 -98.060 9.550 -97.320 ;
        RECT 18.630 -98.060 22.050 -97.320 ;
        RECT 33.630 -98.060 37.050 -97.320 ;
        RECT -44.530 -99.180 -40.535 -98.510 ;
        RECT -35.230 -98.890 -32.230 -98.130 ;
        RECT -113.820 -101.875 -107.190 -101.290 ;
        RECT -103.925 -101.430 -101.420 -100.865 ;
        RECT -92.530 -101.050 -89.625 -100.395 ;
        RECT -92.170 -101.820 -90.150 -101.060 ;
        RECT -63.420 -101.690 -59.425 -101.020 ;
        RECT 139.425 -101.065 141.930 -100.500 ;
        RECT 134.730 -101.965 137.635 -101.310 ;
        RECT -70.800 -103.385 -68.295 -102.820 ;
        RECT -70.760 -105.165 -68.250 -103.405 ;
        RECT -63.035 -103.735 -61.505 -101.975 ;
        RECT -60.845 -103.735 -59.805 -101.975 ;
        RECT 135.090 -103.235 137.110 -101.975 ;
        RECT 139.465 -102.845 141.975 -101.085 ;
        RECT 181.625 -101.120 184.130 -100.555 ;
        RECT 176.930 -102.020 179.835 -101.365 ;
        RECT 142.640 -103.610 145.545 -102.955 ;
        RECT 177.290 -103.290 179.310 -102.030 ;
        RECT 181.665 -102.900 184.175 -101.140 ;
        RECT 225.940 -101.315 228.445 -100.750 ;
        RECT 271.930 -101.145 274.435 -100.580 ;
        RECT 315.700 -100.815 318.205 -100.250 ;
        RECT 361.465 -100.730 363.970 -100.165 ;
        RECT 408.285 -100.540 410.790 -99.975 ;
        RECT 221.245 -102.215 224.150 -101.560 ;
        RECT 143.000 -104.380 145.020 -103.620 ;
        RECT 184.840 -103.665 187.745 -103.010 ;
        RECT 221.605 -103.485 223.625 -102.225 ;
        RECT 225.980 -103.095 228.490 -101.335 ;
        RECT 267.235 -102.045 270.140 -101.390 ;
        RECT 185.200 -104.435 187.220 -103.675 ;
        RECT 229.155 -103.860 232.060 -103.205 ;
        RECT 267.595 -103.315 269.615 -102.055 ;
        RECT 271.970 -102.925 274.480 -101.165 ;
        RECT 311.005 -101.715 313.910 -101.060 ;
        RECT 311.365 -102.985 313.385 -101.725 ;
        RECT 315.740 -102.595 318.250 -100.835 ;
        RECT 356.770 -101.630 359.675 -100.975 ;
        RECT 275.145 -103.690 278.050 -103.035 ;
        RECT 318.915 -103.360 321.820 -102.705 ;
        RECT 357.130 -102.900 359.150 -101.640 ;
        RECT 361.505 -102.510 364.015 -100.750 ;
        RECT 403.590 -101.440 406.495 -100.785 ;
        RECT 364.680 -103.275 367.585 -102.620 ;
        RECT 403.950 -102.710 405.970 -101.450 ;
        RECT 408.325 -102.320 410.835 -100.560 ;
        RECT 411.500 -103.085 414.405 -102.430 ;
        RECT 229.515 -104.630 231.535 -103.870 ;
        RECT 275.505 -104.460 277.525 -103.700 ;
        RECT 319.275 -104.130 321.295 -103.370 ;
        RECT 365.040 -104.045 367.060 -103.285 ;
        RECT 411.860 -103.855 413.880 -103.095 ;
        RECT -67.585 -105.930 -64.680 -105.275 ;
        RECT -67.225 -106.700 -65.205 -105.940 ;
        RECT -36.515 -106.705 -33.515 -105.945 ;
        RECT -110.060 -107.855 -108.040 -107.095 ;
        RECT -87.175 -107.620 -85.155 -106.860 ;
        RECT -36.460 -107.320 -33.530 -106.720 ;
        RECT -32.325 -106.955 -28.345 -106.195 ;
        RECT -27.800 -106.705 -24.800 -105.945 ;
        RECT -23.015 -106.705 -20.015 -105.945 ;
        RECT -27.745 -107.320 -24.815 -106.720 ;
        RECT -22.960 -107.320 -20.030 -106.720 ;
        RECT -18.825 -106.955 -14.845 -106.195 ;
        RECT -14.300 -106.705 -11.300 -105.945 ;
        RECT -9.890 -106.705 -6.890 -105.945 ;
        RECT 3.915 -106.110 5.935 -105.350 ;
        RECT 11.940 -106.120 13.960 -105.360 ;
        RECT -14.245 -107.320 -11.315 -106.720 ;
        RECT -9.835 -107.320 -6.905 -106.720 ;
        RECT 3.390 -106.775 6.295 -106.120 ;
        RECT 11.415 -106.785 14.320 -106.130 ;
        RECT 86.710 -106.255 91.255 -105.465 ;
        RECT -110.420 -108.520 -107.515 -107.865 ;
        RECT -113.595 -110.390 -111.085 -108.630 ;
        RECT -104.730 -110.265 -103.200 -108.505 ;
        RECT -103.180 -110.270 -101.650 -108.510 ;
        RECT -101.635 -110.270 -100.105 -108.510 ;
        RECT -99.080 -110.270 -98.040 -109.010 ;
        RECT -95.085 -109.265 -93.065 -108.005 ;
        RECT -87.535 -108.285 -84.630 -107.630 ;
        RECT -95.445 -109.930 -92.540 -109.275 ;
        RECT -90.710 -110.155 -88.200 -108.395 ;
        RECT -36.500 -109.220 -33.570 -108.620 ;
        RECT -32.315 -109.220 -29.385 -108.620 ;
        RECT -36.515 -109.995 -33.515 -109.235 ;
        RECT -32.330 -109.995 -29.330 -109.235 ;
        RECT -28.785 -109.745 -24.805 -108.985 ;
        RECT -23.000 -109.220 -20.070 -108.620 ;
        RECT -18.815 -109.220 -15.885 -108.620 ;
        RECT -5.240 -108.930 -4.200 -107.670 ;
        RECT -3.175 -108.930 -1.645 -107.170 ;
        RECT -1.630 -108.930 -0.100 -107.170 ;
        RECT -0.080 -108.925 1.450 -107.165 ;
        RECT 6.960 -108.645 9.470 -106.885 ;
        RECT 14.985 -108.655 17.495 -106.895 ;
        RECT -23.015 -109.995 -20.015 -109.235 ;
        RECT -18.830 -109.995 -15.830 -109.235 ;
        RECT -15.285 -109.745 -11.305 -108.985 ;
        RECT 7.005 -109.230 9.510 -108.665 ;
        RECT 15.030 -109.240 17.535 -108.675 ;
        RECT 19.570 -108.885 20.610 -107.625 ;
        RECT 21.635 -108.885 23.165 -107.125 ;
        RECT 23.180 -108.885 24.710 -107.125 ;
        RECT 24.730 -108.880 26.260 -107.120 ;
        RECT 27.635 -108.430 28.675 -107.170 ;
        RECT 29.705 -108.430 30.745 -107.170 ;
        RECT 31.515 -108.430 32.555 -107.170 ;
        RECT 32.985 -108.430 34.025 -107.170 ;
        RECT 34.535 -108.430 35.575 -107.170 ;
        RECT 36.080 -108.430 37.120 -107.170 ;
        RECT 87.195 -107.820 89.215 -106.560 ;
        RECT 97.725 -108.300 101.705 -107.540 ;
        RECT 102.250 -108.050 105.250 -107.290 ;
        RECT 106.435 -108.050 109.435 -107.290 ;
        RECT 33.680 -109.315 37.100 -108.575 ;
        RECT 102.305 -108.665 105.235 -108.065 ;
        RECT 106.490 -108.665 109.420 -108.065 ;
        RECT 111.225 -108.300 115.205 -107.540 ;
        RECT 115.750 -108.050 118.750 -107.290 ;
        RECT 119.935 -108.050 122.935 -107.290 ;
        RECT 115.805 -108.665 118.735 -108.065 ;
        RECT 119.990 -108.665 122.920 -108.065 ;
        RECT -113.635 -110.975 -111.130 -110.410 ;
        RECT -90.750 -110.740 -88.245 -110.175 ;
        RECT -5.240 -110.215 1.390 -109.630 ;
        RECT 19.570 -110.170 26.200 -109.585 ;
        RECT 93.325 -110.565 96.255 -109.965 ;
        RECT 97.735 -110.565 100.665 -109.965 ;
        RECT -104.670 -111.555 -98.040 -110.970 ;
        RECT 93.310 -111.340 96.310 -110.580 ;
        RECT 97.720 -111.340 100.720 -110.580 ;
        RECT 101.265 -111.090 105.245 -110.330 ;
        RECT 106.450 -110.565 109.380 -109.965 ;
        RECT 111.235 -110.565 114.165 -109.965 ;
        RECT 106.435 -111.340 109.435 -110.580 ;
        RECT 111.220 -111.340 114.220 -110.580 ;
        RECT 114.765 -111.090 118.745 -110.330 ;
        RECT 119.950 -110.565 122.880 -109.965 ;
        RECT 138.005 -110.180 140.025 -109.420 ;
        RECT 119.935 -111.340 122.935 -110.580 ;
        RECT 137.645 -110.845 140.550 -110.190 ;
        RECT 180.205 -110.235 182.225 -109.475 ;
        RECT 179.845 -110.900 182.750 -110.245 ;
        RECT 224.520 -110.430 226.540 -109.670 ;
        RECT 270.510 -110.260 272.530 -109.500 ;
        RECT 314.280 -109.930 316.300 -109.170 ;
        RECT 360.045 -109.845 362.065 -109.085 ;
        RECT 406.865 -109.655 408.885 -108.895 ;
        RECT -62.230 -112.500 -60.210 -111.740 ;
        RECT -70.140 -114.145 -68.120 -112.885 ;
        RECT -62.590 -113.165 -59.685 -112.510 ;
        RECT 134.470 -112.715 136.980 -110.955 ;
        RECT -70.500 -114.810 -67.595 -114.155 ;
        RECT -65.765 -115.035 -63.255 -113.275 ;
        RECT 134.430 -113.300 136.935 -112.735 ;
        RECT 142.195 -114.145 143.725 -112.385 ;
        RECT 144.385 -114.145 145.425 -112.385 ;
        RECT 151.665 -113.855 152.705 -112.095 ;
        RECT 154.015 -113.855 155.055 -111.095 ;
        RECT 155.130 -113.855 156.170 -111.095 ;
        RECT 156.270 -113.855 157.800 -111.095 ;
        RECT 157.900 -113.855 158.940 -112.095 ;
        RECT 176.670 -112.770 179.180 -111.010 ;
        RECT 224.160 -111.095 227.065 -110.440 ;
        RECT 270.150 -110.925 273.055 -110.270 ;
        RECT 313.920 -110.595 316.825 -109.940 ;
        RECT 359.685 -110.510 362.590 -109.855 ;
        RECT 406.505 -110.320 409.410 -109.665 ;
        RECT 176.630 -113.355 179.135 -112.790 ;
        RECT -65.805 -115.620 -63.300 -115.055 ;
        RECT 109.260 -115.640 123.155 -114.895 ;
        RECT 141.810 -115.100 145.805 -114.430 ;
        RECT 151.335 -115.170 158.960 -114.105 ;
        RECT 184.395 -114.200 185.925 -112.440 ;
        RECT 186.585 -114.200 187.625 -112.440 ;
        RECT 193.865 -113.910 194.905 -112.150 ;
        RECT 196.215 -113.910 197.255 -111.150 ;
        RECT 197.330 -113.910 198.370 -111.150 ;
        RECT 198.470 -113.910 200.000 -111.150 ;
        RECT 200.100 -113.910 201.140 -112.150 ;
        RECT 220.985 -112.965 223.495 -111.205 ;
        RECT 220.945 -113.550 223.450 -112.985 ;
        RECT 184.010 -115.155 188.005 -114.485 ;
        RECT 193.535 -115.225 201.160 -114.160 ;
        RECT 228.710 -114.395 230.240 -112.635 ;
        RECT 230.900 -114.395 231.940 -112.635 ;
        RECT 238.180 -114.105 239.220 -112.345 ;
        RECT 240.530 -114.105 241.570 -111.345 ;
        RECT 241.645 -114.105 242.685 -111.345 ;
        RECT 242.785 -114.105 244.315 -111.345 ;
        RECT 244.415 -114.105 245.455 -112.345 ;
        RECT 266.975 -112.795 269.485 -111.035 ;
        RECT 266.935 -113.380 269.440 -112.815 ;
        RECT 274.700 -114.225 276.230 -112.465 ;
        RECT 276.890 -114.225 277.930 -112.465 ;
        RECT 284.170 -113.935 285.210 -112.175 ;
        RECT 286.520 -113.935 287.560 -111.175 ;
        RECT 287.635 -113.935 288.675 -111.175 ;
        RECT 288.775 -113.935 290.305 -111.175 ;
        RECT 290.405 -113.935 291.445 -112.175 ;
        RECT 310.745 -112.465 313.255 -110.705 ;
        RECT 310.705 -113.050 313.210 -112.485 ;
        RECT 318.470 -113.895 320.000 -112.135 ;
        RECT 320.660 -113.895 321.700 -112.135 ;
        RECT 327.940 -113.605 328.980 -111.845 ;
        RECT 330.290 -113.605 331.330 -110.845 ;
        RECT 331.405 -113.605 332.445 -110.845 ;
        RECT 332.545 -113.605 334.075 -110.845 ;
        RECT 334.175 -113.605 335.215 -111.845 ;
        RECT 356.510 -112.380 359.020 -110.620 ;
        RECT 356.470 -112.965 358.975 -112.400 ;
        RECT 364.235 -113.810 365.765 -112.050 ;
        RECT 366.425 -113.810 367.465 -112.050 ;
        RECT 373.705 -113.520 374.745 -111.760 ;
        RECT 376.055 -113.520 377.095 -110.760 ;
        RECT 377.170 -113.520 378.210 -110.760 ;
        RECT 378.310 -113.520 379.840 -110.760 ;
        RECT 379.940 -113.520 380.980 -111.760 ;
        RECT 403.330 -112.190 405.840 -110.430 ;
        RECT 403.290 -112.775 405.795 -112.210 ;
        RECT 411.055 -113.620 412.585 -111.860 ;
        RECT 413.245 -113.620 414.285 -111.860 ;
        RECT 420.525 -113.330 421.565 -111.570 ;
        RECT 422.875 -113.330 423.915 -110.570 ;
        RECT 423.990 -113.330 425.030 -110.570 ;
        RECT 425.130 -113.330 426.660 -110.570 ;
        RECT 426.760 -113.330 427.800 -111.570 ;
        RECT 228.325 -115.350 232.320 -114.680 ;
        RECT 237.850 -115.420 245.475 -114.355 ;
        RECT 274.315 -115.180 278.310 -114.510 ;
        RECT 283.840 -115.250 291.465 -114.185 ;
        RECT 318.085 -114.850 322.080 -114.180 ;
        RECT 327.610 -114.920 335.235 -113.855 ;
        RECT 363.850 -114.765 367.845 -114.095 ;
        RECT 373.375 -114.835 381.000 -113.770 ;
        RECT 410.670 -114.575 414.665 -113.905 ;
        RECT 420.195 -114.645 427.820 -113.580 ;
        RECT -75.885 -119.150 -72.885 -118.390 ;
        RECT -71.700 -119.150 -68.700 -118.390 ;
        RECT -75.870 -119.765 -72.940 -119.165 ;
        RECT -71.685 -119.765 -68.755 -119.165 ;
        RECT -68.155 -119.400 -64.175 -118.640 ;
        RECT -62.385 -119.150 -59.385 -118.390 ;
        RECT -58.200 -119.150 -55.200 -118.390 ;
        RECT -62.370 -119.765 -59.440 -119.165 ;
        RECT -58.185 -119.765 -55.255 -119.165 ;
        RECT -54.655 -119.400 -50.675 -118.640 ;
        RECT 86.565 -119.375 89.810 -118.670 ;
        RECT 91.295 -119.375 94.540 -118.670 ;
        RECT 96.050 -119.040 102.680 -118.455 ;
        RECT -36.515 -120.485 -33.515 -119.725 ;
        RECT -32.330 -120.485 -29.330 -119.725 ;
        RECT -88.365 -121.810 -84.370 -121.140 ;
        RECT -75.830 -121.665 -72.900 -121.065 ;
        RECT -95.745 -123.505 -93.240 -122.940 ;
        RECT -106.750 -126.280 -105.220 -125.020 ;
        RECT -102.225 -126.285 -100.695 -125.025 ;
        RECT -95.705 -125.285 -93.195 -123.525 ;
        RECT -87.980 -123.855 -86.450 -122.095 ;
        RECT -85.790 -123.855 -84.750 -122.095 ;
        RECT -75.885 -122.440 -72.885 -121.680 ;
        RECT -71.695 -122.190 -67.715 -121.430 ;
        RECT -67.115 -121.665 -64.185 -121.065 ;
        RECT -62.330 -121.665 -59.400 -121.065 ;
        RECT -67.170 -122.440 -64.170 -121.680 ;
        RECT -62.385 -122.440 -59.385 -121.680 ;
        RECT -58.195 -122.190 -54.215 -121.430 ;
        RECT -53.615 -121.665 -50.685 -121.065 ;
        RECT -49.205 -121.665 -46.275 -121.065 ;
        RECT -36.500 -121.100 -33.570 -120.500 ;
        RECT -32.315 -121.100 -29.385 -120.500 ;
        RECT -28.785 -120.735 -24.805 -119.975 ;
        RECT -23.015 -120.485 -20.015 -119.725 ;
        RECT -18.830 -120.485 -15.830 -119.725 ;
        RECT -23.000 -121.100 -20.070 -120.500 ;
        RECT -18.815 -121.100 -15.885 -120.500 ;
        RECT -15.285 -120.735 -11.305 -119.975 ;
        RECT -5.240 -120.090 1.390 -119.505 ;
        RECT 19.570 -120.135 26.200 -119.550 ;
        RECT -53.670 -122.440 -50.670 -121.680 ;
        RECT -49.260 -122.440 -46.260 -121.680 ;
        RECT -44.015 -122.895 -42.975 -121.135 ;
        RECT -42.315 -122.895 -40.785 -121.135 ;
        RECT -5.240 -122.050 -4.200 -120.790 ;
        RECT -36.460 -123.000 -33.530 -122.400 ;
        RECT -44.395 -123.850 -40.400 -123.180 ;
        RECT -36.515 -123.775 -33.515 -123.015 ;
        RECT -32.325 -123.525 -28.345 -122.765 ;
        RECT -27.745 -123.000 -24.815 -122.400 ;
        RECT -22.960 -123.000 -20.030 -122.400 ;
        RECT -27.800 -123.775 -24.800 -123.015 ;
        RECT -23.015 -123.775 -20.015 -123.015 ;
        RECT -18.825 -123.525 -14.845 -122.765 ;
        RECT -14.245 -123.000 -11.315 -122.400 ;
        RECT -9.835 -123.000 -6.905 -122.400 ;
        RECT -3.175 -122.550 -1.645 -120.790 ;
        RECT -1.630 -122.550 -0.100 -120.790 ;
        RECT -0.080 -122.555 1.450 -120.795 ;
        RECT 7.005 -121.055 9.510 -120.490 ;
        RECT 15.030 -121.045 17.535 -120.480 ;
        RECT 6.960 -122.835 9.470 -121.075 ;
        RECT 14.985 -122.825 17.495 -121.065 ;
        RECT 19.570 -122.095 20.610 -120.835 ;
        RECT 21.635 -122.595 23.165 -120.835 ;
        RECT 23.180 -122.595 24.710 -120.835 ;
        RECT 24.730 -122.600 26.260 -120.840 ;
        RECT 33.680 -121.145 37.100 -120.405 ;
        RECT 87.170 -120.910 88.700 -119.650 ;
        RECT 91.900 -120.910 93.430 -119.650 ;
        RECT 27.635 -122.550 28.675 -121.290 ;
        RECT 29.705 -122.550 30.745 -121.290 ;
        RECT 31.515 -122.550 32.555 -121.290 ;
        RECT 32.985 -122.550 34.025 -121.290 ;
        RECT 34.535 -122.550 35.575 -121.290 ;
        RECT 36.080 -122.550 37.120 -121.290 ;
        RECT 95.990 -121.505 97.520 -119.745 ;
        RECT 97.540 -121.500 99.070 -119.740 ;
        RECT 99.085 -121.500 100.615 -119.740 ;
        RECT 101.640 -121.000 102.680 -119.740 ;
        RECT 105.535 -120.270 106.575 -119.010 ;
        RECT 106.585 -120.270 107.625 -119.010 ;
        RECT 109.685 -119.725 110.725 -115.965 ;
        RECT 111.685 -119.725 112.725 -115.965 ;
        RECT 114.685 -119.725 115.725 -115.965 ;
        RECT 116.685 -119.725 117.725 -115.965 ;
        RECT 119.685 -119.725 120.725 -115.965 ;
        RECT 121.685 -119.725 122.725 -115.965 ;
        RECT 139.385 -118.330 141.890 -117.765 ;
        RECT 134.690 -119.230 137.595 -118.575 ;
        RECT 135.050 -120.500 137.070 -119.240 ;
        RECT 139.425 -120.110 141.935 -118.350 ;
        RECT 157.725 -118.485 160.230 -117.920 ;
        RECT 181.585 -118.385 184.090 -117.820 ;
        RECT 153.030 -119.385 155.935 -118.730 ;
        RECT 105.430 -121.215 108.085 -120.550 ;
        RECT 142.600 -120.875 145.505 -120.220 ;
        RECT 153.390 -120.655 155.410 -119.395 ;
        RECT 157.765 -120.265 160.275 -118.505 ;
        RECT 176.890 -119.285 179.795 -118.630 ;
        RECT 105.300 -121.830 108.230 -121.230 ;
        RECT 142.960 -121.645 144.980 -120.885 ;
        RECT 160.940 -121.030 163.845 -120.375 ;
        RECT 177.250 -120.555 179.270 -119.295 ;
        RECT 181.625 -120.165 184.135 -118.405 ;
        RECT 199.925 -118.540 202.430 -117.975 ;
        RECT 195.230 -119.440 198.135 -118.785 ;
        RECT 184.800 -120.930 187.705 -120.275 ;
        RECT 195.590 -120.710 197.610 -119.450 ;
        RECT 199.965 -120.320 202.475 -118.560 ;
        RECT 225.900 -118.580 228.405 -118.015 ;
        RECT 221.205 -119.480 224.110 -118.825 ;
        RECT 161.300 -121.800 163.320 -121.040 ;
        RECT 185.160 -121.700 187.180 -120.940 ;
        RECT 203.140 -121.085 206.045 -120.430 ;
        RECT 221.565 -120.750 223.585 -119.490 ;
        RECT 225.940 -120.360 228.450 -118.600 ;
        RECT 244.240 -118.735 246.745 -118.170 ;
        RECT 271.890 -118.410 274.395 -117.845 ;
        RECT 239.545 -119.635 242.450 -118.980 ;
        RECT 105.285 -122.605 108.285 -121.845 ;
        RECT 203.500 -121.855 205.520 -121.095 ;
        RECT 229.115 -121.125 232.020 -120.470 ;
        RECT 239.905 -120.905 241.925 -119.645 ;
        RECT 244.280 -120.515 246.790 -118.755 ;
        RECT 267.195 -119.310 270.100 -118.655 ;
        RECT 267.555 -120.580 269.575 -119.320 ;
        RECT 271.930 -120.190 274.440 -118.430 ;
        RECT 290.230 -118.565 292.735 -118.000 ;
        RECT 315.660 -118.080 318.165 -117.515 ;
        RECT 285.535 -119.465 288.440 -118.810 ;
        RECT 229.475 -121.895 231.495 -121.135 ;
        RECT 247.455 -121.280 250.360 -120.625 ;
        RECT 275.105 -120.955 278.010 -120.300 ;
        RECT 285.895 -120.735 287.915 -119.475 ;
        RECT 290.270 -120.345 292.780 -118.585 ;
        RECT 310.965 -118.980 313.870 -118.325 ;
        RECT 311.325 -120.250 313.345 -118.990 ;
        RECT 315.700 -119.860 318.210 -118.100 ;
        RECT 334.000 -118.235 336.505 -117.670 ;
        RECT 361.425 -117.995 363.930 -117.430 ;
        RECT 329.305 -119.135 332.210 -118.480 ;
        RECT 247.815 -122.050 249.835 -121.290 ;
        RECT 275.465 -121.725 277.485 -120.965 ;
        RECT 293.445 -121.110 296.350 -120.455 ;
        RECT 318.875 -120.625 321.780 -119.970 ;
        RECT 329.665 -120.405 331.685 -119.145 ;
        RECT 334.040 -120.015 336.550 -118.255 ;
        RECT 356.730 -118.895 359.635 -118.240 ;
        RECT 293.805 -121.880 295.825 -121.120 ;
        RECT 319.235 -121.395 321.255 -120.635 ;
        RECT 337.215 -120.780 340.120 -120.125 ;
        RECT 357.090 -120.165 359.110 -118.905 ;
        RECT 361.465 -119.775 363.975 -118.015 ;
        RECT 379.765 -118.150 382.270 -117.585 ;
        RECT 408.245 -117.805 410.750 -117.240 ;
        RECT 375.070 -119.050 377.975 -118.395 ;
        RECT 364.640 -120.540 367.545 -119.885 ;
        RECT 375.430 -120.320 377.450 -119.060 ;
        RECT 379.805 -119.930 382.315 -118.170 ;
        RECT 403.550 -118.705 406.455 -118.050 ;
        RECT 403.910 -119.975 405.930 -118.715 ;
        RECT 408.285 -119.585 410.795 -117.825 ;
        RECT 426.585 -117.960 429.090 -117.395 ;
        RECT 421.890 -118.860 424.795 -118.205 ;
        RECT 337.575 -121.550 339.595 -120.790 ;
        RECT 365.000 -121.310 367.020 -120.550 ;
        RECT 382.980 -120.695 385.885 -120.040 ;
        RECT 411.460 -120.350 414.365 -119.695 ;
        RECT 422.250 -120.130 424.270 -118.870 ;
        RECT 426.625 -119.740 429.135 -117.980 ;
        RECT 383.340 -121.465 385.360 -120.705 ;
        RECT 411.820 -121.120 413.840 -120.360 ;
        RECT 429.800 -120.505 432.705 -119.850 ;
        RECT 430.160 -121.275 432.180 -120.515 ;
        RECT -14.300 -123.775 -11.300 -123.015 ;
        RECT -9.890 -123.775 -6.890 -123.015 ;
        RECT 3.390 -123.600 6.295 -122.945 ;
        RECT 11.415 -123.590 14.320 -122.935 ;
        RECT 3.915 -124.370 5.935 -123.610 ;
        RECT 11.940 -124.360 13.960 -123.600 ;
        RECT -92.530 -126.050 -89.625 -125.395 ;
        RECT -112.780 -127.995 -110.760 -126.735 ;
        RECT -107.355 -127.260 -104.110 -126.555 ;
        RECT -102.830 -127.265 -99.585 -126.560 ;
        RECT -92.170 -126.820 -90.150 -126.060 ;
        RECT 137.965 -127.445 139.985 -126.685 ;
        RECT 137.605 -128.110 140.510 -127.455 ;
        RECT 156.305 -127.600 158.325 -126.840 ;
        RECT 180.165 -127.500 182.185 -126.740 ;
        RECT -113.265 -129.090 -108.720 -128.300 ;
        RECT 134.430 -129.980 136.940 -128.220 ;
        RECT 155.945 -128.265 158.850 -127.610 ;
        RECT 179.805 -128.165 182.710 -127.510 ;
        RECT 198.505 -127.655 200.525 -126.895 ;
        RECT 52.670 -130.830 55.670 -130.070 ;
        RECT 57.080 -130.830 60.080 -130.070 ;
        RECT -114.465 -131.765 -107.835 -131.180 ;
        RECT 52.685 -131.445 55.615 -130.845 ;
        RECT 57.095 -131.445 60.025 -130.845 ;
        RECT 60.625 -131.080 64.605 -130.320 ;
        RECT 65.795 -130.830 68.795 -130.070 ;
        RECT 70.580 -130.830 73.580 -130.070 ;
        RECT 65.810 -131.445 68.740 -130.845 ;
        RECT 70.595 -131.445 73.525 -130.845 ;
        RECT 74.125 -131.080 78.105 -130.320 ;
        RECT 79.295 -130.830 82.295 -130.070 ;
        RECT 134.390 -130.565 136.895 -130.000 ;
        RECT 79.310 -131.445 82.240 -130.845 ;
        RECT 142.155 -131.410 143.685 -129.650 ;
        RECT 144.345 -131.410 145.385 -129.650 ;
        RECT 152.770 -130.135 155.280 -128.375 ;
        RECT 152.730 -130.720 155.235 -130.155 ;
        RECT 160.495 -131.565 162.025 -129.805 ;
        RECT 162.685 -131.565 163.725 -129.805 ;
        RECT 176.630 -130.035 179.140 -128.275 ;
        RECT 198.145 -128.320 201.050 -127.665 ;
        RECT 224.480 -127.695 226.500 -126.935 ;
        RECT 224.120 -128.360 227.025 -127.705 ;
        RECT 242.820 -127.850 244.840 -127.090 ;
        RECT 270.470 -127.525 272.490 -126.765 ;
        RECT 176.590 -130.620 179.095 -130.055 ;
        RECT 184.355 -131.465 185.885 -129.705 ;
        RECT 186.545 -131.465 187.585 -129.705 ;
        RECT 194.970 -130.190 197.480 -128.430 ;
        RECT 194.930 -130.775 197.435 -130.210 ;
        RECT 202.695 -131.620 204.225 -129.860 ;
        RECT 204.885 -131.620 205.925 -129.860 ;
        RECT 220.945 -130.230 223.455 -128.470 ;
        RECT 242.460 -128.515 245.365 -127.860 ;
        RECT 270.110 -128.190 273.015 -127.535 ;
        RECT 288.810 -127.680 290.830 -126.920 ;
        RECT 314.240 -127.195 316.260 -126.435 ;
        RECT 220.905 -130.815 223.410 -130.250 ;
        RECT 228.670 -131.660 230.200 -129.900 ;
        RECT 230.860 -131.660 231.900 -129.900 ;
        RECT 239.285 -130.385 241.795 -128.625 ;
        RECT 239.245 -130.970 241.750 -130.405 ;
        RECT -114.465 -133.725 -113.425 -132.465 ;
        RECT -112.400 -134.225 -110.870 -132.465 ;
        RECT -110.855 -134.225 -109.325 -132.465 ;
        RECT -109.305 -134.230 -107.775 -132.470 ;
        RECT -87.175 -132.620 -85.155 -131.860 ;
        RECT -31.370 -132.400 -27.950 -131.660 ;
        RECT -18.870 -132.400 -15.450 -131.660 ;
        RECT -6.370 -132.400 -2.950 -131.660 ;
        RECT 6.130 -132.400 9.550 -131.660 ;
        RECT 18.630 -132.400 22.050 -131.660 ;
        RECT 33.630 -132.400 37.050 -131.660 ;
        RECT 141.770 -132.365 145.765 -131.695 ;
        RECT 160.110 -132.520 164.105 -131.850 ;
        RECT 183.970 -132.420 187.965 -131.750 ;
        RECT 247.010 -131.815 248.540 -130.055 ;
        RECT 249.200 -131.815 250.240 -130.055 ;
        RECT 266.935 -130.060 269.445 -128.300 ;
        RECT 288.450 -128.345 291.355 -127.690 ;
        RECT 313.880 -127.860 316.785 -127.205 ;
        RECT 332.580 -127.350 334.600 -126.590 ;
        RECT 360.005 -127.110 362.025 -126.350 ;
        RECT 266.895 -130.645 269.400 -130.080 ;
        RECT 274.660 -131.490 276.190 -129.730 ;
        RECT 276.850 -131.490 277.890 -129.730 ;
        RECT 285.275 -130.215 287.785 -128.455 ;
        RECT 310.705 -129.730 313.215 -127.970 ;
        RECT 332.220 -128.015 335.125 -127.360 ;
        RECT 359.645 -127.775 362.550 -127.120 ;
        RECT 378.345 -127.265 380.365 -126.505 ;
        RECT 406.825 -126.920 408.845 -126.160 ;
        RECT 285.235 -130.800 287.740 -130.235 ;
        RECT 293.000 -131.645 294.530 -129.885 ;
        RECT 295.190 -131.645 296.230 -129.885 ;
        RECT 310.665 -130.315 313.170 -129.750 ;
        RECT 318.430 -131.160 319.960 -129.400 ;
        RECT 320.620 -131.160 321.660 -129.400 ;
        RECT 329.045 -129.885 331.555 -128.125 ;
        RECT 329.005 -130.470 331.510 -129.905 ;
        RECT 336.770 -131.315 338.300 -129.555 ;
        RECT 338.960 -131.315 340.000 -129.555 ;
        RECT 356.470 -129.645 358.980 -127.885 ;
        RECT 377.985 -127.930 380.890 -127.275 ;
        RECT 406.465 -127.585 409.370 -126.930 ;
        RECT 425.165 -127.075 427.185 -126.315 ;
        RECT 356.430 -130.230 358.935 -129.665 ;
        RECT 364.195 -131.075 365.725 -129.315 ;
        RECT 366.385 -131.075 367.425 -129.315 ;
        RECT 374.810 -129.800 377.320 -128.040 ;
        RECT 403.290 -129.455 405.800 -127.695 ;
        RECT 424.805 -127.740 427.710 -127.085 ;
        RECT 374.770 -130.385 377.275 -129.820 ;
        RECT 382.535 -131.230 384.065 -129.470 ;
        RECT 384.725 -131.230 385.765 -129.470 ;
        RECT 403.250 -130.040 405.755 -129.475 ;
        RECT 411.015 -130.885 412.545 -129.125 ;
        RECT 413.205 -130.885 414.245 -129.125 ;
        RECT 421.630 -129.610 424.140 -127.850 ;
        RECT 421.590 -130.195 424.095 -129.630 ;
        RECT 429.355 -131.040 430.885 -129.280 ;
        RECT 431.545 -131.040 432.585 -129.280 ;
        RECT -95.085 -134.265 -93.065 -133.005 ;
        RECT -87.535 -133.285 -84.630 -132.630 ;
        RECT -95.445 -134.930 -92.540 -134.275 ;
        RECT -90.710 -135.155 -88.200 -133.395 ;
        RECT -37.415 -133.805 -36.375 -132.545 ;
        RECT -35.345 -133.805 -34.305 -132.545 ;
        RECT -33.535 -133.805 -32.495 -132.545 ;
        RECT -32.065 -133.805 -31.025 -132.545 ;
        RECT -30.515 -133.805 -29.475 -132.545 ;
        RECT -28.970 -133.805 -27.930 -132.545 ;
        RECT -24.915 -133.805 -23.875 -132.545 ;
        RECT -22.845 -133.805 -21.805 -132.545 ;
        RECT -21.035 -133.805 -19.995 -132.545 ;
        RECT -19.565 -133.805 -18.525 -132.545 ;
        RECT -18.015 -133.805 -16.975 -132.545 ;
        RECT -16.470 -133.805 -15.430 -132.545 ;
        RECT -12.415 -133.805 -11.375 -132.545 ;
        RECT -10.345 -133.805 -9.305 -132.545 ;
        RECT -8.535 -133.805 -7.495 -132.545 ;
        RECT -7.065 -133.805 -6.025 -132.545 ;
        RECT -5.515 -133.805 -4.475 -132.545 ;
        RECT -3.970 -133.805 -2.930 -132.545 ;
        RECT 0.085 -133.805 1.125 -132.545 ;
        RECT 2.155 -133.805 3.195 -132.545 ;
        RECT 3.965 -133.805 5.005 -132.545 ;
        RECT 5.435 -133.805 6.475 -132.545 ;
        RECT 6.985 -133.805 8.025 -132.545 ;
        RECT 8.530 -133.805 9.570 -132.545 ;
        RECT 12.585 -133.805 13.625 -132.545 ;
        RECT 14.655 -133.805 15.695 -132.545 ;
        RECT 16.465 -133.805 17.505 -132.545 ;
        RECT 17.935 -133.805 18.975 -132.545 ;
        RECT 19.485 -133.805 20.525 -132.545 ;
        RECT 21.030 -133.805 22.070 -132.545 ;
        RECT 27.585 -133.805 28.625 -132.545 ;
        RECT 29.655 -133.805 30.695 -132.545 ;
        RECT 31.465 -133.805 32.505 -132.545 ;
        RECT 32.935 -133.805 33.975 -132.545 ;
        RECT 34.485 -133.805 35.525 -132.545 ;
        RECT 36.030 -133.805 37.070 -132.545 ;
        RECT 202.310 -132.575 206.305 -131.905 ;
        RECT 228.285 -132.615 232.280 -131.945 ;
        RECT 57.085 -133.870 61.065 -133.110 ;
        RECT 61.665 -133.345 64.595 -132.745 ;
        RECT 65.850 -133.345 68.780 -132.745 ;
        RECT 61.610 -134.120 64.610 -133.360 ;
        RECT 65.795 -134.120 68.795 -133.360 ;
        RECT 70.585 -133.870 74.565 -133.110 ;
        RECT 75.165 -133.345 78.095 -132.745 ;
        RECT 79.350 -133.345 82.280 -132.745 ;
        RECT 246.625 -132.770 250.620 -132.100 ;
        RECT 274.275 -132.445 278.270 -131.775 ;
        RECT 292.615 -132.600 296.610 -131.930 ;
        RECT 318.045 -132.115 322.040 -131.445 ;
        RECT 336.385 -132.270 340.380 -131.600 ;
        RECT 363.810 -132.030 367.805 -131.360 ;
        RECT 382.150 -132.185 386.145 -131.515 ;
        RECT 410.630 -131.840 414.625 -131.170 ;
        RECT 428.970 -131.995 432.965 -131.325 ;
        RECT 75.110 -134.120 78.110 -133.360 ;
        RECT 79.295 -134.120 82.295 -133.360 ;
        RECT -90.750 -135.740 -88.245 -135.175 ;
        RECT -135.280 -206.525 -134.390 -170.260 ;
        RECT -134.230 -206.345 -131.970 -170.395 ;
        RECT -72.395 -177.470 -69.395 -176.710 ;
        RECT -68.210 -177.470 -65.210 -176.710 ;
        RECT -72.380 -178.085 -69.450 -177.485 ;
        RECT -68.195 -178.085 -65.265 -177.485 ;
        RECT -64.665 -177.720 -60.685 -176.960 ;
        RECT -58.895 -177.470 -55.895 -176.710 ;
        RECT -54.710 -177.470 -51.710 -176.710 ;
        RECT -58.880 -178.085 -55.950 -177.485 ;
        RECT -54.695 -178.085 -51.765 -177.485 ;
        RECT -51.165 -177.720 -47.185 -176.960 ;
        RECT -84.875 -179.765 -80.880 -179.095 ;
        RECT -72.340 -179.985 -69.410 -179.385 ;
        RECT -96.860 -181.265 -94.840 -180.505 ;
        RECT -110.390 -183.540 -108.860 -181.780 ;
        RECT -108.840 -183.545 -107.310 -181.785 ;
        RECT -107.295 -183.545 -105.765 -181.785 ;
        RECT -97.220 -181.930 -94.315 -181.275 ;
        RECT -92.255 -181.460 -89.750 -180.895 ;
        RECT -104.740 -183.545 -103.700 -182.285 ;
        RECT -100.395 -183.800 -97.885 -182.040 ;
        RECT -92.215 -183.240 -89.705 -181.480 ;
        RECT -84.490 -181.810 -82.960 -180.050 ;
        RECT -82.300 -181.810 -81.260 -180.050 ;
        RECT -72.395 -180.760 -69.395 -180.000 ;
        RECT -68.205 -180.510 -64.225 -179.750 ;
        RECT -63.625 -179.985 -60.695 -179.385 ;
        RECT -58.840 -179.985 -55.910 -179.385 ;
        RECT -63.680 -180.760 -60.680 -180.000 ;
        RECT -58.895 -180.760 -55.895 -180.000 ;
        RECT -54.705 -180.510 -50.725 -179.750 ;
        RECT -50.125 -179.985 -47.195 -179.385 ;
        RECT -45.715 -179.985 -42.785 -179.385 ;
        RECT -50.180 -180.760 -47.180 -180.000 ;
        RECT -45.770 -180.760 -42.770 -180.000 ;
        RECT -40.660 -181.180 -39.620 -179.420 ;
        RECT -38.960 -181.180 -37.430 -179.420 ;
        RECT -33.925 -180.130 -32.885 -178.870 ;
        RECT -31.855 -180.130 -30.815 -178.870 ;
        RECT -30.045 -180.130 -29.005 -178.870 ;
        RECT -28.575 -180.130 -27.535 -178.870 ;
        RECT -27.025 -180.130 -25.985 -178.870 ;
        RECT -25.480 -180.130 -24.440 -178.870 ;
        RECT -21.425 -180.130 -20.385 -178.870 ;
        RECT -19.355 -180.130 -18.315 -178.870 ;
        RECT -17.545 -180.130 -16.505 -178.870 ;
        RECT -16.075 -180.130 -15.035 -178.870 ;
        RECT -14.525 -180.130 -13.485 -178.870 ;
        RECT -12.980 -180.130 -11.940 -178.870 ;
        RECT -8.925 -180.130 -7.885 -178.870 ;
        RECT -6.855 -180.130 -5.815 -178.870 ;
        RECT -5.045 -180.130 -4.005 -178.870 ;
        RECT -3.575 -180.130 -2.535 -178.870 ;
        RECT -2.025 -180.130 -0.985 -178.870 ;
        RECT -0.480 -180.130 0.560 -178.870 ;
        RECT 3.575 -180.130 4.615 -178.870 ;
        RECT 5.645 -180.130 6.685 -178.870 ;
        RECT 7.455 -180.130 8.495 -178.870 ;
        RECT 8.925 -180.130 9.965 -178.870 ;
        RECT 10.475 -180.130 11.515 -178.870 ;
        RECT 12.020 -180.130 13.060 -178.870 ;
        RECT 16.075 -180.130 17.115 -178.870 ;
        RECT 18.145 -180.130 19.185 -178.870 ;
        RECT 19.955 -180.130 20.995 -178.870 ;
        RECT 21.425 -180.130 22.465 -178.870 ;
        RECT 22.975 -180.130 24.015 -178.870 ;
        RECT 24.520 -180.130 25.560 -178.870 ;
        RECT 31.075 -180.130 32.115 -178.870 ;
        RECT 33.145 -180.130 34.185 -178.870 ;
        RECT 34.955 -180.130 35.995 -178.870 ;
        RECT 36.425 -180.130 37.465 -178.870 ;
        RECT 37.975 -180.130 39.015 -178.870 ;
        RECT 39.520 -180.130 40.560 -178.870 ;
        RECT -31.725 -181.070 -28.795 -180.470 ;
        RECT -27.880 -181.015 -24.460 -180.275 ;
        RECT -15.380 -181.015 -11.960 -180.275 ;
        RECT -2.880 -181.015 0.540 -180.275 ;
        RECT 9.620 -181.015 13.040 -180.275 ;
        RECT 22.120 -181.015 25.540 -180.275 ;
        RECT 37.120 -181.015 40.540 -180.275 ;
        RECT -41.040 -182.135 -37.045 -181.465 ;
        RECT -31.740 -181.845 -28.740 -181.085 ;
        RECT -110.330 -184.830 -103.700 -184.245 ;
        RECT -100.435 -184.385 -97.930 -183.820 ;
        RECT -89.040 -184.005 -86.135 -183.350 ;
        RECT -88.680 -184.775 -86.660 -184.015 ;
        RECT -59.930 -184.645 -55.935 -183.975 ;
        RECT 142.915 -184.020 145.420 -183.455 ;
        RECT 138.220 -184.920 141.125 -184.265 ;
        RECT -67.310 -186.340 -64.805 -185.775 ;
        RECT -67.270 -188.120 -64.760 -186.360 ;
        RECT -59.545 -186.690 -58.015 -184.930 ;
        RECT -57.355 -186.690 -56.315 -184.930 ;
        RECT 138.580 -186.190 140.600 -184.930 ;
        RECT 142.955 -185.800 145.465 -184.040 ;
        RECT 185.115 -184.075 187.620 -183.510 ;
        RECT 180.420 -184.975 183.325 -184.320 ;
        RECT 146.130 -186.565 149.035 -185.910 ;
        RECT 180.780 -186.245 182.800 -184.985 ;
        RECT 185.155 -185.855 187.665 -184.095 ;
        RECT 229.430 -184.270 231.935 -183.705 ;
        RECT 275.420 -184.100 277.925 -183.535 ;
        RECT 319.190 -183.770 321.695 -183.205 ;
        RECT 364.955 -183.685 367.460 -183.120 ;
        RECT 411.775 -183.495 414.280 -182.930 ;
        RECT 224.735 -185.170 227.640 -184.515 ;
        RECT 146.490 -187.335 148.510 -186.575 ;
        RECT 188.330 -186.620 191.235 -185.965 ;
        RECT 225.095 -186.440 227.115 -185.180 ;
        RECT 229.470 -186.050 231.980 -184.290 ;
        RECT 270.725 -185.000 273.630 -184.345 ;
        RECT 188.690 -187.390 190.710 -186.630 ;
        RECT 232.645 -186.815 235.550 -186.160 ;
        RECT 271.085 -186.270 273.105 -185.010 ;
        RECT 275.460 -185.880 277.970 -184.120 ;
        RECT 314.495 -184.670 317.400 -184.015 ;
        RECT 314.855 -185.940 316.875 -184.680 ;
        RECT 319.230 -185.550 321.740 -183.790 ;
        RECT 360.260 -184.585 363.165 -183.930 ;
        RECT 278.635 -186.645 281.540 -185.990 ;
        RECT 322.405 -186.315 325.310 -185.660 ;
        RECT 360.620 -185.855 362.640 -184.595 ;
        RECT 364.995 -185.465 367.505 -183.705 ;
        RECT 407.080 -184.395 409.985 -183.740 ;
        RECT 368.170 -186.230 371.075 -185.575 ;
        RECT 407.440 -185.665 409.460 -184.405 ;
        RECT 411.815 -185.275 414.325 -183.515 ;
        RECT 414.990 -186.040 417.895 -185.385 ;
        RECT 233.005 -187.585 235.025 -186.825 ;
        RECT 278.995 -187.415 281.015 -186.655 ;
        RECT 322.765 -187.085 324.785 -186.325 ;
        RECT 368.530 -187.000 370.550 -186.240 ;
        RECT 415.350 -186.810 417.370 -186.050 ;
        RECT -64.095 -188.885 -61.190 -188.230 ;
        RECT -63.735 -189.655 -61.715 -188.895 ;
        RECT -33.025 -189.660 -30.025 -188.900 ;
        RECT -106.570 -190.810 -104.550 -190.050 ;
        RECT -83.685 -190.575 -81.665 -189.815 ;
        RECT -32.970 -190.275 -30.040 -189.675 ;
        RECT -28.835 -189.910 -24.855 -189.150 ;
        RECT -24.310 -189.660 -21.310 -188.900 ;
        RECT -19.525 -189.660 -16.525 -188.900 ;
        RECT -24.255 -190.275 -21.325 -189.675 ;
        RECT -19.470 -190.275 -16.540 -189.675 ;
        RECT -15.335 -189.910 -11.355 -189.150 ;
        RECT -10.810 -189.660 -7.810 -188.900 ;
        RECT -6.400 -189.660 -3.400 -188.900 ;
        RECT 7.405 -189.065 9.425 -188.305 ;
        RECT 15.430 -189.075 17.450 -188.315 ;
        RECT -10.755 -190.275 -7.825 -189.675 ;
        RECT -6.345 -190.275 -3.415 -189.675 ;
        RECT 6.880 -189.730 9.785 -189.075 ;
        RECT 14.905 -189.740 17.810 -189.085 ;
        RECT 90.200 -189.210 94.745 -188.420 ;
        RECT -106.930 -191.475 -104.025 -190.820 ;
        RECT -110.105 -193.345 -107.595 -191.585 ;
        RECT -101.240 -193.220 -99.710 -191.460 ;
        RECT -99.690 -193.225 -98.160 -191.465 ;
        RECT -98.145 -193.225 -96.615 -191.465 ;
        RECT -95.590 -193.225 -94.550 -191.965 ;
        RECT -91.595 -192.220 -89.575 -190.960 ;
        RECT -84.045 -191.240 -81.140 -190.585 ;
        RECT -91.955 -192.885 -89.050 -192.230 ;
        RECT -87.220 -193.110 -84.710 -191.350 ;
        RECT -33.010 -192.175 -30.080 -191.575 ;
        RECT -28.825 -192.175 -25.895 -191.575 ;
        RECT -33.025 -192.950 -30.025 -192.190 ;
        RECT -28.840 -192.950 -25.840 -192.190 ;
        RECT -25.295 -192.700 -21.315 -191.940 ;
        RECT -19.510 -192.175 -16.580 -191.575 ;
        RECT -15.325 -192.175 -12.395 -191.575 ;
        RECT -1.750 -191.885 -0.710 -190.625 ;
        RECT 0.315 -191.885 1.845 -190.125 ;
        RECT 1.860 -191.885 3.390 -190.125 ;
        RECT 3.410 -191.880 4.940 -190.120 ;
        RECT 10.450 -191.600 12.960 -189.840 ;
        RECT 18.475 -191.610 20.985 -189.850 ;
        RECT -19.525 -192.950 -16.525 -192.190 ;
        RECT -15.340 -192.950 -12.340 -192.190 ;
        RECT -11.795 -192.700 -7.815 -191.940 ;
        RECT 10.495 -192.185 13.000 -191.620 ;
        RECT 18.520 -192.195 21.025 -191.630 ;
        RECT 23.060 -191.840 24.100 -190.580 ;
        RECT 25.125 -191.840 26.655 -190.080 ;
        RECT 26.670 -191.840 28.200 -190.080 ;
        RECT 28.220 -191.835 29.750 -190.075 ;
        RECT 31.125 -191.385 32.165 -190.125 ;
        RECT 33.195 -191.385 34.235 -190.125 ;
        RECT 35.005 -191.385 36.045 -190.125 ;
        RECT 36.475 -191.385 37.515 -190.125 ;
        RECT 38.025 -191.385 39.065 -190.125 ;
        RECT 39.570 -191.385 40.610 -190.125 ;
        RECT 90.685 -190.775 92.705 -189.515 ;
        RECT 101.215 -191.255 105.195 -190.495 ;
        RECT 105.740 -191.005 108.740 -190.245 ;
        RECT 109.925 -191.005 112.925 -190.245 ;
        RECT 37.170 -192.270 40.590 -191.530 ;
        RECT 105.795 -191.620 108.725 -191.020 ;
        RECT 109.980 -191.620 112.910 -191.020 ;
        RECT 114.715 -191.255 118.695 -190.495 ;
        RECT 119.240 -191.005 122.240 -190.245 ;
        RECT 123.425 -191.005 126.425 -190.245 ;
        RECT 119.295 -191.620 122.225 -191.020 ;
        RECT 123.480 -191.620 126.410 -191.020 ;
        RECT -110.145 -193.930 -107.640 -193.365 ;
        RECT -87.260 -193.695 -84.755 -193.130 ;
        RECT -1.750 -193.170 4.880 -192.585 ;
        RECT 23.060 -193.125 29.690 -192.540 ;
        RECT 96.815 -193.520 99.745 -192.920 ;
        RECT 101.225 -193.520 104.155 -192.920 ;
        RECT -101.180 -194.510 -94.550 -193.925 ;
        RECT 96.800 -194.295 99.800 -193.535 ;
        RECT 101.210 -194.295 104.210 -193.535 ;
        RECT 104.755 -194.045 108.735 -193.285 ;
        RECT 109.940 -193.520 112.870 -192.920 ;
        RECT 114.725 -193.520 117.655 -192.920 ;
        RECT 109.925 -194.295 112.925 -193.535 ;
        RECT 114.710 -194.295 117.710 -193.535 ;
        RECT 118.255 -194.045 122.235 -193.285 ;
        RECT 123.440 -193.520 126.370 -192.920 ;
        RECT 141.495 -193.135 143.515 -192.375 ;
        RECT 123.425 -194.295 126.425 -193.535 ;
        RECT 141.135 -193.800 144.040 -193.145 ;
        RECT 183.695 -193.190 185.715 -192.430 ;
        RECT 183.335 -193.855 186.240 -193.200 ;
        RECT 228.010 -193.385 230.030 -192.625 ;
        RECT 274.000 -193.215 276.020 -192.455 ;
        RECT 317.770 -192.885 319.790 -192.125 ;
        RECT 363.535 -192.800 365.555 -192.040 ;
        RECT 410.355 -192.610 412.375 -191.850 ;
        RECT -58.740 -195.455 -56.720 -194.695 ;
        RECT -66.650 -197.100 -64.630 -195.840 ;
        RECT -59.100 -196.120 -56.195 -195.465 ;
        RECT 137.960 -195.670 140.470 -193.910 ;
        RECT -67.010 -197.765 -64.105 -197.110 ;
        RECT -62.275 -197.990 -59.765 -196.230 ;
        RECT 137.920 -196.255 140.425 -195.690 ;
        RECT 145.685 -197.100 147.215 -195.340 ;
        RECT 147.875 -197.100 148.915 -195.340 ;
        RECT 155.155 -196.810 156.195 -195.050 ;
        RECT 157.505 -196.810 158.545 -194.050 ;
        RECT 158.620 -196.810 159.660 -194.050 ;
        RECT 159.760 -196.810 161.290 -194.050 ;
        RECT 161.390 -196.810 162.430 -195.050 ;
        RECT 180.160 -195.725 182.670 -193.965 ;
        RECT 227.650 -194.050 230.555 -193.395 ;
        RECT 273.640 -193.880 276.545 -193.225 ;
        RECT 317.410 -193.550 320.315 -192.895 ;
        RECT 363.175 -193.465 366.080 -192.810 ;
        RECT 409.995 -193.275 412.900 -192.620 ;
        RECT 180.120 -196.310 182.625 -195.745 ;
        RECT -62.315 -198.575 -59.810 -198.010 ;
        RECT 112.750 -198.595 126.645 -197.850 ;
        RECT 145.300 -198.055 149.295 -197.385 ;
        RECT 154.825 -198.125 162.450 -197.060 ;
        RECT 187.885 -197.155 189.415 -195.395 ;
        RECT 190.075 -197.155 191.115 -195.395 ;
        RECT 197.355 -196.865 198.395 -195.105 ;
        RECT 199.705 -196.865 200.745 -194.105 ;
        RECT 200.820 -196.865 201.860 -194.105 ;
        RECT 201.960 -196.865 203.490 -194.105 ;
        RECT 203.590 -196.865 204.630 -195.105 ;
        RECT 224.475 -195.920 226.985 -194.160 ;
        RECT 224.435 -196.505 226.940 -195.940 ;
        RECT 187.500 -198.110 191.495 -197.440 ;
        RECT 197.025 -198.180 204.650 -197.115 ;
        RECT 232.200 -197.350 233.730 -195.590 ;
        RECT 234.390 -197.350 235.430 -195.590 ;
        RECT 241.670 -197.060 242.710 -195.300 ;
        RECT 244.020 -197.060 245.060 -194.300 ;
        RECT 245.135 -197.060 246.175 -194.300 ;
        RECT 246.275 -197.060 247.805 -194.300 ;
        RECT 247.905 -197.060 248.945 -195.300 ;
        RECT 270.465 -195.750 272.975 -193.990 ;
        RECT 270.425 -196.335 272.930 -195.770 ;
        RECT 278.190 -197.180 279.720 -195.420 ;
        RECT 280.380 -197.180 281.420 -195.420 ;
        RECT 287.660 -196.890 288.700 -195.130 ;
        RECT 290.010 -196.890 291.050 -194.130 ;
        RECT 291.125 -196.890 292.165 -194.130 ;
        RECT 292.265 -196.890 293.795 -194.130 ;
        RECT 293.895 -196.890 294.935 -195.130 ;
        RECT 314.235 -195.420 316.745 -193.660 ;
        RECT 314.195 -196.005 316.700 -195.440 ;
        RECT 321.960 -196.850 323.490 -195.090 ;
        RECT 324.150 -196.850 325.190 -195.090 ;
        RECT 331.430 -196.560 332.470 -194.800 ;
        RECT 333.780 -196.560 334.820 -193.800 ;
        RECT 334.895 -196.560 335.935 -193.800 ;
        RECT 336.035 -196.560 337.565 -193.800 ;
        RECT 337.665 -196.560 338.705 -194.800 ;
        RECT 360.000 -195.335 362.510 -193.575 ;
        RECT 359.960 -195.920 362.465 -195.355 ;
        RECT 367.725 -196.765 369.255 -195.005 ;
        RECT 369.915 -196.765 370.955 -195.005 ;
        RECT 377.195 -196.475 378.235 -194.715 ;
        RECT 379.545 -196.475 380.585 -193.715 ;
        RECT 380.660 -196.475 381.700 -193.715 ;
        RECT 381.800 -196.475 383.330 -193.715 ;
        RECT 383.430 -196.475 384.470 -194.715 ;
        RECT 406.820 -195.145 409.330 -193.385 ;
        RECT 406.780 -195.730 409.285 -195.165 ;
        RECT 414.545 -196.575 416.075 -194.815 ;
        RECT 416.735 -196.575 417.775 -194.815 ;
        RECT 424.015 -196.285 425.055 -194.525 ;
        RECT 426.365 -196.285 427.405 -193.525 ;
        RECT 427.480 -196.285 428.520 -193.525 ;
        RECT 428.620 -196.285 430.150 -193.525 ;
        RECT 430.250 -196.285 431.290 -194.525 ;
        RECT 231.815 -198.305 235.810 -197.635 ;
        RECT 241.340 -198.375 248.965 -197.310 ;
        RECT 277.805 -198.135 281.800 -197.465 ;
        RECT 287.330 -198.205 294.955 -197.140 ;
        RECT 321.575 -197.805 325.570 -197.135 ;
        RECT 331.100 -197.875 338.725 -196.810 ;
        RECT 367.340 -197.720 371.335 -197.050 ;
        RECT 376.865 -197.790 384.490 -196.725 ;
        RECT 414.160 -197.530 418.155 -196.860 ;
        RECT 423.685 -197.600 431.310 -196.535 ;
        RECT -72.395 -202.105 -69.395 -201.345 ;
        RECT -68.210 -202.105 -65.210 -201.345 ;
        RECT -72.380 -202.720 -69.450 -202.120 ;
        RECT -68.195 -202.720 -65.265 -202.120 ;
        RECT -64.665 -202.355 -60.685 -201.595 ;
        RECT -58.895 -202.105 -55.895 -201.345 ;
        RECT -54.710 -202.105 -51.710 -201.345 ;
        RECT -58.880 -202.720 -55.950 -202.120 ;
        RECT -54.695 -202.720 -51.765 -202.120 ;
        RECT -51.165 -202.355 -47.185 -201.595 ;
        RECT 90.055 -202.330 93.300 -201.625 ;
        RECT 94.785 -202.330 98.030 -201.625 ;
        RECT 99.540 -201.995 106.170 -201.410 ;
        RECT -33.025 -203.440 -30.025 -202.680 ;
        RECT -28.840 -203.440 -25.840 -202.680 ;
        RECT -84.875 -204.765 -80.880 -204.095 ;
        RECT -72.340 -204.620 -69.410 -204.020 ;
        RECT -92.255 -206.460 -89.750 -205.895 ;
        RECT -103.260 -209.235 -101.730 -207.975 ;
        RECT -98.735 -209.240 -97.205 -207.980 ;
        RECT -92.215 -208.240 -89.705 -206.480 ;
        RECT -84.490 -206.810 -82.960 -205.050 ;
        RECT -82.300 -206.810 -81.260 -205.050 ;
        RECT -72.395 -205.395 -69.395 -204.635 ;
        RECT -68.205 -205.145 -64.225 -204.385 ;
        RECT -63.625 -204.620 -60.695 -204.020 ;
        RECT -58.840 -204.620 -55.910 -204.020 ;
        RECT -63.680 -205.395 -60.680 -204.635 ;
        RECT -58.895 -205.395 -55.895 -204.635 ;
        RECT -54.705 -205.145 -50.725 -204.385 ;
        RECT -50.125 -204.620 -47.195 -204.020 ;
        RECT -45.715 -204.620 -42.785 -204.020 ;
        RECT -33.010 -204.055 -30.080 -203.455 ;
        RECT -28.825 -204.055 -25.895 -203.455 ;
        RECT -25.295 -203.690 -21.315 -202.930 ;
        RECT -19.525 -203.440 -16.525 -202.680 ;
        RECT -15.340 -203.440 -12.340 -202.680 ;
        RECT -19.510 -204.055 -16.580 -203.455 ;
        RECT -15.325 -204.055 -12.395 -203.455 ;
        RECT -11.795 -203.690 -7.815 -202.930 ;
        RECT -1.750 -203.045 4.880 -202.460 ;
        RECT 23.060 -203.090 29.690 -202.505 ;
        RECT -50.180 -205.395 -47.180 -204.635 ;
        RECT -45.770 -205.395 -42.770 -204.635 ;
        RECT -40.525 -205.850 -39.485 -204.090 ;
        RECT -38.825 -205.850 -37.295 -204.090 ;
        RECT -1.750 -205.005 -0.710 -203.745 ;
        RECT -32.970 -205.955 -30.040 -205.355 ;
        RECT -40.905 -206.805 -36.910 -206.135 ;
        RECT -33.025 -206.730 -30.025 -205.970 ;
        RECT -28.835 -206.480 -24.855 -205.720 ;
        RECT -24.255 -205.955 -21.325 -205.355 ;
        RECT -19.470 -205.955 -16.540 -205.355 ;
        RECT -24.310 -206.730 -21.310 -205.970 ;
        RECT -19.525 -206.730 -16.525 -205.970 ;
        RECT -15.335 -206.480 -11.355 -205.720 ;
        RECT -10.755 -205.955 -7.825 -205.355 ;
        RECT -6.345 -205.955 -3.415 -205.355 ;
        RECT 0.315 -205.505 1.845 -203.745 ;
        RECT 1.860 -205.505 3.390 -203.745 ;
        RECT 3.410 -205.510 4.940 -203.750 ;
        RECT 10.495 -204.010 13.000 -203.445 ;
        RECT 18.520 -204.000 21.025 -203.435 ;
        RECT 10.450 -205.790 12.960 -204.030 ;
        RECT 18.475 -205.780 20.985 -204.020 ;
        RECT 23.060 -205.050 24.100 -203.790 ;
        RECT 25.125 -205.550 26.655 -203.790 ;
        RECT 26.670 -205.550 28.200 -203.790 ;
        RECT 28.220 -205.555 29.750 -203.795 ;
        RECT 37.170 -204.100 40.590 -203.360 ;
        RECT 90.660 -203.865 92.190 -202.605 ;
        RECT 95.390 -203.865 96.920 -202.605 ;
        RECT 31.125 -205.505 32.165 -204.245 ;
        RECT 33.195 -205.505 34.235 -204.245 ;
        RECT 35.005 -205.505 36.045 -204.245 ;
        RECT 36.475 -205.505 37.515 -204.245 ;
        RECT 38.025 -205.505 39.065 -204.245 ;
        RECT 39.570 -205.505 40.610 -204.245 ;
        RECT 99.480 -204.460 101.010 -202.700 ;
        RECT 101.030 -204.455 102.560 -202.695 ;
        RECT 102.575 -204.455 104.105 -202.695 ;
        RECT 105.130 -203.955 106.170 -202.695 ;
        RECT 109.025 -203.225 110.065 -201.965 ;
        RECT 110.075 -203.225 111.115 -201.965 ;
        RECT 113.175 -202.680 114.215 -198.920 ;
        RECT 115.175 -202.680 116.215 -198.920 ;
        RECT 118.175 -202.680 119.215 -198.920 ;
        RECT 120.175 -202.680 121.215 -198.920 ;
        RECT 123.175 -202.680 124.215 -198.920 ;
        RECT 125.175 -202.680 126.215 -198.920 ;
        RECT 142.875 -201.285 145.380 -200.720 ;
        RECT 138.180 -202.185 141.085 -201.530 ;
        RECT 138.540 -203.455 140.560 -202.195 ;
        RECT 142.915 -203.065 145.425 -201.305 ;
        RECT 161.215 -201.440 163.720 -200.875 ;
        RECT 185.075 -201.340 187.580 -200.775 ;
        RECT 156.520 -202.340 159.425 -201.685 ;
        RECT 108.920 -204.170 111.575 -203.505 ;
        RECT 146.090 -203.830 148.995 -203.175 ;
        RECT 156.880 -203.610 158.900 -202.350 ;
        RECT 161.255 -203.220 163.765 -201.460 ;
        RECT 180.380 -202.240 183.285 -201.585 ;
        RECT 108.790 -204.785 111.720 -204.185 ;
        RECT 146.450 -204.600 148.470 -203.840 ;
        RECT 164.430 -203.985 167.335 -203.330 ;
        RECT 180.740 -203.510 182.760 -202.250 ;
        RECT 185.115 -203.120 187.625 -201.360 ;
        RECT 203.415 -201.495 205.920 -200.930 ;
        RECT 198.720 -202.395 201.625 -201.740 ;
        RECT 188.290 -203.885 191.195 -203.230 ;
        RECT 199.080 -203.665 201.100 -202.405 ;
        RECT 203.455 -203.275 205.965 -201.515 ;
        RECT 229.390 -201.535 231.895 -200.970 ;
        RECT 224.695 -202.435 227.600 -201.780 ;
        RECT 164.790 -204.755 166.810 -203.995 ;
        RECT 188.650 -204.655 190.670 -203.895 ;
        RECT 206.630 -204.040 209.535 -203.385 ;
        RECT 225.055 -203.705 227.075 -202.445 ;
        RECT 229.430 -203.315 231.940 -201.555 ;
        RECT 247.730 -201.690 250.235 -201.125 ;
        RECT 275.380 -201.365 277.885 -200.800 ;
        RECT 243.035 -202.590 245.940 -201.935 ;
        RECT 108.775 -205.560 111.775 -204.800 ;
        RECT 206.990 -204.810 209.010 -204.050 ;
        RECT 232.605 -204.080 235.510 -203.425 ;
        RECT 243.395 -203.860 245.415 -202.600 ;
        RECT 247.770 -203.470 250.280 -201.710 ;
        RECT 270.685 -202.265 273.590 -201.610 ;
        RECT 271.045 -203.535 273.065 -202.275 ;
        RECT 275.420 -203.145 277.930 -201.385 ;
        RECT 293.720 -201.520 296.225 -200.955 ;
        RECT 319.150 -201.035 321.655 -200.470 ;
        RECT 289.025 -202.420 291.930 -201.765 ;
        RECT 232.965 -204.850 234.985 -204.090 ;
        RECT 250.945 -204.235 253.850 -203.580 ;
        RECT 278.595 -203.910 281.500 -203.255 ;
        RECT 289.385 -203.690 291.405 -202.430 ;
        RECT 293.760 -203.300 296.270 -201.540 ;
        RECT 314.455 -201.935 317.360 -201.280 ;
        RECT 314.815 -203.205 316.835 -201.945 ;
        RECT 319.190 -202.815 321.700 -201.055 ;
        RECT 337.490 -201.190 339.995 -200.625 ;
        RECT 364.915 -200.950 367.420 -200.385 ;
        RECT 332.795 -202.090 335.700 -201.435 ;
        RECT 251.305 -205.005 253.325 -204.245 ;
        RECT 278.955 -204.680 280.975 -203.920 ;
        RECT 296.935 -204.065 299.840 -203.410 ;
        RECT 322.365 -203.580 325.270 -202.925 ;
        RECT 333.155 -203.360 335.175 -202.100 ;
        RECT 337.530 -202.970 340.040 -201.210 ;
        RECT 360.220 -201.850 363.125 -201.195 ;
        RECT 297.295 -204.835 299.315 -204.075 ;
        RECT 322.725 -204.350 324.745 -203.590 ;
        RECT 340.705 -203.735 343.610 -203.080 ;
        RECT 360.580 -203.120 362.600 -201.860 ;
        RECT 364.955 -202.730 367.465 -200.970 ;
        RECT 383.255 -201.105 385.760 -200.540 ;
        RECT 411.735 -200.760 414.240 -200.195 ;
        RECT 378.560 -202.005 381.465 -201.350 ;
        RECT 368.130 -203.495 371.035 -202.840 ;
        RECT 378.920 -203.275 380.940 -202.015 ;
        RECT 383.295 -202.885 385.805 -201.125 ;
        RECT 407.040 -201.660 409.945 -201.005 ;
        RECT 407.400 -202.930 409.420 -201.670 ;
        RECT 411.775 -202.540 414.285 -200.780 ;
        RECT 430.075 -200.915 432.580 -200.350 ;
        RECT 425.380 -201.815 428.285 -201.160 ;
        RECT 341.065 -204.505 343.085 -203.745 ;
        RECT 368.490 -204.265 370.510 -203.505 ;
        RECT 386.470 -203.650 389.375 -202.995 ;
        RECT 414.950 -203.305 417.855 -202.650 ;
        RECT 425.740 -203.085 427.760 -201.825 ;
        RECT 430.115 -202.695 432.625 -200.935 ;
        RECT 386.830 -204.420 388.850 -203.660 ;
        RECT 415.310 -204.075 417.330 -203.315 ;
        RECT 433.290 -203.460 436.195 -202.805 ;
        RECT 433.650 -204.230 435.670 -203.470 ;
        RECT -10.810 -206.730 -7.810 -205.970 ;
        RECT -6.400 -206.730 -3.400 -205.970 ;
        RECT 6.880 -206.555 9.785 -205.900 ;
        RECT 14.905 -206.545 17.810 -205.890 ;
        RECT 7.405 -207.325 9.425 -206.565 ;
        RECT 15.430 -207.315 17.450 -206.555 ;
        RECT -89.040 -209.005 -86.135 -208.350 ;
        RECT -109.290 -210.950 -107.270 -209.690 ;
        RECT -103.865 -210.215 -100.620 -209.510 ;
        RECT -99.340 -210.220 -96.095 -209.515 ;
        RECT -88.680 -209.775 -86.660 -209.015 ;
        RECT 141.455 -210.400 143.475 -209.640 ;
        RECT 141.095 -211.065 144.000 -210.410 ;
        RECT 159.795 -210.555 161.815 -209.795 ;
        RECT 183.655 -210.455 185.675 -209.695 ;
        RECT -109.775 -212.045 -105.230 -211.255 ;
        RECT 137.920 -212.935 140.430 -211.175 ;
        RECT 159.435 -211.220 162.340 -210.565 ;
        RECT 183.295 -211.120 186.200 -210.465 ;
        RECT 201.995 -210.610 204.015 -209.850 ;
        RECT 56.160 -213.785 59.160 -213.025 ;
        RECT 60.570 -213.785 63.570 -213.025 ;
        RECT -110.975 -214.720 -104.345 -214.135 ;
        RECT 56.175 -214.400 59.105 -213.800 ;
        RECT 60.585 -214.400 63.515 -213.800 ;
        RECT 64.115 -214.035 68.095 -213.275 ;
        RECT 69.285 -213.785 72.285 -213.025 ;
        RECT 74.070 -213.785 77.070 -213.025 ;
        RECT 69.300 -214.400 72.230 -213.800 ;
        RECT 74.085 -214.400 77.015 -213.800 ;
        RECT 77.615 -214.035 81.595 -213.275 ;
        RECT 82.785 -213.785 85.785 -213.025 ;
        RECT 137.880 -213.520 140.385 -212.955 ;
        RECT 82.800 -214.400 85.730 -213.800 ;
        RECT 145.645 -214.365 147.175 -212.605 ;
        RECT 147.835 -214.365 148.875 -212.605 ;
        RECT 156.260 -213.090 158.770 -211.330 ;
        RECT 156.220 -213.675 158.725 -213.110 ;
        RECT 163.985 -214.520 165.515 -212.760 ;
        RECT 166.175 -214.520 167.215 -212.760 ;
        RECT 180.120 -212.990 182.630 -211.230 ;
        RECT 201.635 -211.275 204.540 -210.620 ;
        RECT 227.970 -210.650 229.990 -209.890 ;
        RECT 227.610 -211.315 230.515 -210.660 ;
        RECT 246.310 -210.805 248.330 -210.045 ;
        RECT 273.960 -210.480 275.980 -209.720 ;
        RECT 180.080 -213.575 182.585 -213.010 ;
        RECT 187.845 -214.420 189.375 -212.660 ;
        RECT 190.035 -214.420 191.075 -212.660 ;
        RECT 198.460 -213.145 200.970 -211.385 ;
        RECT 198.420 -213.730 200.925 -213.165 ;
        RECT 206.185 -214.575 207.715 -212.815 ;
        RECT 208.375 -214.575 209.415 -212.815 ;
        RECT 224.435 -213.185 226.945 -211.425 ;
        RECT 245.950 -211.470 248.855 -210.815 ;
        RECT 273.600 -211.145 276.505 -210.490 ;
        RECT 292.300 -210.635 294.320 -209.875 ;
        RECT 317.730 -210.150 319.750 -209.390 ;
        RECT 224.395 -213.770 226.900 -213.205 ;
        RECT 232.160 -214.615 233.690 -212.855 ;
        RECT 234.350 -214.615 235.390 -212.855 ;
        RECT 242.775 -213.340 245.285 -211.580 ;
        RECT 242.735 -213.925 245.240 -213.360 ;
        RECT -110.975 -216.680 -109.935 -215.420 ;
        RECT -108.910 -217.180 -107.380 -215.420 ;
        RECT -107.365 -217.180 -105.835 -215.420 ;
        RECT -105.815 -217.185 -104.285 -215.425 ;
        RECT -83.685 -215.575 -81.665 -214.815 ;
        RECT -27.880 -215.355 -24.460 -214.615 ;
        RECT -15.380 -215.355 -11.960 -214.615 ;
        RECT -2.880 -215.355 0.540 -214.615 ;
        RECT 9.620 -215.355 13.040 -214.615 ;
        RECT 22.120 -215.355 25.540 -214.615 ;
        RECT 37.120 -215.355 40.540 -214.615 ;
        RECT 145.260 -215.320 149.255 -214.650 ;
        RECT 163.600 -215.475 167.595 -214.805 ;
        RECT 187.460 -215.375 191.455 -214.705 ;
        RECT 250.500 -214.770 252.030 -213.010 ;
        RECT 252.690 -214.770 253.730 -213.010 ;
        RECT 270.425 -213.015 272.935 -211.255 ;
        RECT 291.940 -211.300 294.845 -210.645 ;
        RECT 317.370 -210.815 320.275 -210.160 ;
        RECT 336.070 -210.305 338.090 -209.545 ;
        RECT 363.495 -210.065 365.515 -209.305 ;
        RECT 270.385 -213.600 272.890 -213.035 ;
        RECT 278.150 -214.445 279.680 -212.685 ;
        RECT 280.340 -214.445 281.380 -212.685 ;
        RECT 288.765 -213.170 291.275 -211.410 ;
        RECT 314.195 -212.685 316.705 -210.925 ;
        RECT 335.710 -210.970 338.615 -210.315 ;
        RECT 363.135 -210.730 366.040 -210.075 ;
        RECT 381.835 -210.220 383.855 -209.460 ;
        RECT 410.315 -209.875 412.335 -209.115 ;
        RECT 288.725 -213.755 291.230 -213.190 ;
        RECT 296.490 -214.600 298.020 -212.840 ;
        RECT 298.680 -214.600 299.720 -212.840 ;
        RECT 314.155 -213.270 316.660 -212.705 ;
        RECT 321.920 -214.115 323.450 -212.355 ;
        RECT 324.110 -214.115 325.150 -212.355 ;
        RECT 332.535 -212.840 335.045 -211.080 ;
        RECT 332.495 -213.425 335.000 -212.860 ;
        RECT 340.260 -214.270 341.790 -212.510 ;
        RECT 342.450 -214.270 343.490 -212.510 ;
        RECT 359.960 -212.600 362.470 -210.840 ;
        RECT 381.475 -210.885 384.380 -210.230 ;
        RECT 409.955 -210.540 412.860 -209.885 ;
        RECT 428.655 -210.030 430.675 -209.270 ;
        RECT 359.920 -213.185 362.425 -212.620 ;
        RECT 367.685 -214.030 369.215 -212.270 ;
        RECT 369.875 -214.030 370.915 -212.270 ;
        RECT 378.300 -212.755 380.810 -210.995 ;
        RECT 406.780 -212.410 409.290 -210.650 ;
        RECT 428.295 -210.695 431.200 -210.040 ;
        RECT 378.260 -213.340 380.765 -212.775 ;
        RECT 386.025 -214.185 387.555 -212.425 ;
        RECT 388.215 -214.185 389.255 -212.425 ;
        RECT 406.740 -212.995 409.245 -212.430 ;
        RECT 414.505 -213.840 416.035 -212.080 ;
        RECT 416.695 -213.840 417.735 -212.080 ;
        RECT 425.120 -212.565 427.630 -210.805 ;
        RECT 425.080 -213.150 427.585 -212.585 ;
        RECT 432.845 -213.995 434.375 -212.235 ;
        RECT 435.035 -213.995 436.075 -212.235 ;
        RECT -91.595 -217.220 -89.575 -215.960 ;
        RECT -84.045 -216.240 -81.140 -215.585 ;
        RECT -91.955 -217.885 -89.050 -217.230 ;
        RECT -87.220 -218.110 -84.710 -216.350 ;
        RECT -33.925 -216.760 -32.885 -215.500 ;
        RECT -31.855 -216.760 -30.815 -215.500 ;
        RECT -30.045 -216.760 -29.005 -215.500 ;
        RECT -28.575 -216.760 -27.535 -215.500 ;
        RECT -27.025 -216.760 -25.985 -215.500 ;
        RECT -25.480 -216.760 -24.440 -215.500 ;
        RECT -21.425 -216.760 -20.385 -215.500 ;
        RECT -19.355 -216.760 -18.315 -215.500 ;
        RECT -17.545 -216.760 -16.505 -215.500 ;
        RECT -16.075 -216.760 -15.035 -215.500 ;
        RECT -14.525 -216.760 -13.485 -215.500 ;
        RECT -12.980 -216.760 -11.940 -215.500 ;
        RECT -8.925 -216.760 -7.885 -215.500 ;
        RECT -6.855 -216.760 -5.815 -215.500 ;
        RECT -5.045 -216.760 -4.005 -215.500 ;
        RECT -3.575 -216.760 -2.535 -215.500 ;
        RECT -2.025 -216.760 -0.985 -215.500 ;
        RECT -0.480 -216.760 0.560 -215.500 ;
        RECT 3.575 -216.760 4.615 -215.500 ;
        RECT 5.645 -216.760 6.685 -215.500 ;
        RECT 7.455 -216.760 8.495 -215.500 ;
        RECT 8.925 -216.760 9.965 -215.500 ;
        RECT 10.475 -216.760 11.515 -215.500 ;
        RECT 12.020 -216.760 13.060 -215.500 ;
        RECT 16.075 -216.760 17.115 -215.500 ;
        RECT 18.145 -216.760 19.185 -215.500 ;
        RECT 19.955 -216.760 20.995 -215.500 ;
        RECT 21.425 -216.760 22.465 -215.500 ;
        RECT 22.975 -216.760 24.015 -215.500 ;
        RECT 24.520 -216.760 25.560 -215.500 ;
        RECT 31.075 -216.760 32.115 -215.500 ;
        RECT 33.145 -216.760 34.185 -215.500 ;
        RECT 34.955 -216.760 35.995 -215.500 ;
        RECT 36.425 -216.760 37.465 -215.500 ;
        RECT 37.975 -216.760 39.015 -215.500 ;
        RECT 39.520 -216.760 40.560 -215.500 ;
        RECT 205.800 -215.530 209.795 -214.860 ;
        RECT 231.775 -215.570 235.770 -214.900 ;
        RECT 60.575 -216.825 64.555 -216.065 ;
        RECT 65.155 -216.300 68.085 -215.700 ;
        RECT 69.340 -216.300 72.270 -215.700 ;
        RECT 65.100 -217.075 68.100 -216.315 ;
        RECT 69.285 -217.075 72.285 -216.315 ;
        RECT 74.075 -216.825 78.055 -216.065 ;
        RECT 78.655 -216.300 81.585 -215.700 ;
        RECT 82.840 -216.300 85.770 -215.700 ;
        RECT 250.115 -215.725 254.110 -215.055 ;
        RECT 277.765 -215.400 281.760 -214.730 ;
        RECT 296.105 -215.555 300.100 -214.885 ;
        RECT 321.535 -215.070 325.530 -214.400 ;
        RECT 339.875 -215.225 343.870 -214.555 ;
        RECT 367.300 -214.985 371.295 -214.315 ;
        RECT 385.640 -215.140 389.635 -214.470 ;
        RECT 414.120 -214.795 418.115 -214.125 ;
        RECT 432.460 -214.950 436.455 -214.280 ;
        RECT 78.600 -217.075 81.600 -216.315 ;
        RECT 82.785 -217.075 85.785 -216.315 ;
        RECT -87.260 -218.695 -84.755 -218.130 ;
        RECT -144.380 -297.250 -143.490 -260.985 ;
        RECT -143.330 -297.070 -141.070 -261.120 ;
        RECT -68.880 -268.025 -65.880 -267.265 ;
        RECT -64.695 -268.025 -61.695 -267.265 ;
        RECT -68.865 -268.640 -65.935 -268.040 ;
        RECT -64.680 -268.640 -61.750 -268.040 ;
        RECT -61.150 -268.275 -57.170 -267.515 ;
        RECT -55.380 -268.025 -52.380 -267.265 ;
        RECT -51.195 -268.025 -48.195 -267.265 ;
        RECT -55.365 -268.640 -52.435 -268.040 ;
        RECT -51.180 -268.640 -48.250 -268.040 ;
        RECT -47.650 -268.275 -43.670 -267.515 ;
        RECT -81.360 -270.320 -77.365 -269.650 ;
        RECT -68.825 -270.540 -65.895 -269.940 ;
        RECT -93.345 -271.820 -91.325 -271.060 ;
        RECT -106.875 -274.095 -105.345 -272.335 ;
        RECT -105.325 -274.100 -103.795 -272.340 ;
        RECT -103.780 -274.100 -102.250 -272.340 ;
        RECT -93.705 -272.485 -90.800 -271.830 ;
        RECT -88.740 -272.015 -86.235 -271.450 ;
        RECT -101.225 -274.100 -100.185 -272.840 ;
        RECT -96.880 -274.355 -94.370 -272.595 ;
        RECT -88.700 -273.795 -86.190 -272.035 ;
        RECT -80.975 -272.365 -79.445 -270.605 ;
        RECT -78.785 -272.365 -77.745 -270.605 ;
        RECT -68.880 -271.315 -65.880 -270.555 ;
        RECT -64.690 -271.065 -60.710 -270.305 ;
        RECT -60.110 -270.540 -57.180 -269.940 ;
        RECT -55.325 -270.540 -52.395 -269.940 ;
        RECT -60.165 -271.315 -57.165 -270.555 ;
        RECT -55.380 -271.315 -52.380 -270.555 ;
        RECT -51.190 -271.065 -47.210 -270.305 ;
        RECT -46.610 -270.540 -43.680 -269.940 ;
        RECT -42.200 -270.540 -39.270 -269.940 ;
        RECT -46.665 -271.315 -43.665 -270.555 ;
        RECT -42.255 -271.315 -39.255 -270.555 ;
        RECT -37.145 -271.735 -36.105 -269.975 ;
        RECT -35.445 -271.735 -33.915 -269.975 ;
        RECT -30.410 -270.685 -29.370 -269.425 ;
        RECT -28.340 -270.685 -27.300 -269.425 ;
        RECT -26.530 -270.685 -25.490 -269.425 ;
        RECT -25.060 -270.685 -24.020 -269.425 ;
        RECT -23.510 -270.685 -22.470 -269.425 ;
        RECT -21.965 -270.685 -20.925 -269.425 ;
        RECT -17.910 -270.685 -16.870 -269.425 ;
        RECT -15.840 -270.685 -14.800 -269.425 ;
        RECT -14.030 -270.685 -12.990 -269.425 ;
        RECT -12.560 -270.685 -11.520 -269.425 ;
        RECT -11.010 -270.685 -9.970 -269.425 ;
        RECT -9.465 -270.685 -8.425 -269.425 ;
        RECT -5.410 -270.685 -4.370 -269.425 ;
        RECT -3.340 -270.685 -2.300 -269.425 ;
        RECT -1.530 -270.685 -0.490 -269.425 ;
        RECT -0.060 -270.685 0.980 -269.425 ;
        RECT 1.490 -270.685 2.530 -269.425 ;
        RECT 3.035 -270.685 4.075 -269.425 ;
        RECT 7.090 -270.685 8.130 -269.425 ;
        RECT 9.160 -270.685 10.200 -269.425 ;
        RECT 10.970 -270.685 12.010 -269.425 ;
        RECT 12.440 -270.685 13.480 -269.425 ;
        RECT 13.990 -270.685 15.030 -269.425 ;
        RECT 15.535 -270.685 16.575 -269.425 ;
        RECT 19.590 -270.685 20.630 -269.425 ;
        RECT 21.660 -270.685 22.700 -269.425 ;
        RECT 23.470 -270.685 24.510 -269.425 ;
        RECT 24.940 -270.685 25.980 -269.425 ;
        RECT 26.490 -270.685 27.530 -269.425 ;
        RECT 28.035 -270.685 29.075 -269.425 ;
        RECT 34.590 -270.685 35.630 -269.425 ;
        RECT 36.660 -270.685 37.700 -269.425 ;
        RECT 38.470 -270.685 39.510 -269.425 ;
        RECT 39.940 -270.685 40.980 -269.425 ;
        RECT 41.490 -270.685 42.530 -269.425 ;
        RECT 43.035 -270.685 44.075 -269.425 ;
        RECT -28.210 -271.625 -25.280 -271.025 ;
        RECT -24.365 -271.570 -20.945 -270.830 ;
        RECT -11.865 -271.570 -8.445 -270.830 ;
        RECT 0.635 -271.570 4.055 -270.830 ;
        RECT 13.135 -271.570 16.555 -270.830 ;
        RECT 25.635 -271.570 29.055 -270.830 ;
        RECT 40.635 -271.570 44.055 -270.830 ;
        RECT -37.525 -272.690 -33.530 -272.020 ;
        RECT -28.225 -272.400 -25.225 -271.640 ;
        RECT -106.815 -275.385 -100.185 -274.800 ;
        RECT -96.920 -274.940 -94.415 -274.375 ;
        RECT -85.525 -274.560 -82.620 -273.905 ;
        RECT -85.165 -275.330 -83.145 -274.570 ;
        RECT -56.415 -275.200 -52.420 -274.530 ;
        RECT 146.430 -274.575 148.935 -274.010 ;
        RECT 141.735 -275.475 144.640 -274.820 ;
        RECT -63.795 -276.895 -61.290 -276.330 ;
        RECT -63.755 -278.675 -61.245 -276.915 ;
        RECT -56.030 -277.245 -54.500 -275.485 ;
        RECT -53.840 -277.245 -52.800 -275.485 ;
        RECT 142.095 -276.745 144.115 -275.485 ;
        RECT 146.470 -276.355 148.980 -274.595 ;
        RECT 188.630 -274.630 191.135 -274.065 ;
        RECT 183.935 -275.530 186.840 -274.875 ;
        RECT 149.645 -277.120 152.550 -276.465 ;
        RECT 184.295 -276.800 186.315 -275.540 ;
        RECT 188.670 -276.410 191.180 -274.650 ;
        RECT 232.945 -274.825 235.450 -274.260 ;
        RECT 278.935 -274.655 281.440 -274.090 ;
        RECT 322.705 -274.325 325.210 -273.760 ;
        RECT 368.470 -274.240 370.975 -273.675 ;
        RECT 415.290 -274.050 417.795 -273.485 ;
        RECT 228.250 -275.725 231.155 -275.070 ;
        RECT 150.005 -277.890 152.025 -277.130 ;
        RECT 191.845 -277.175 194.750 -276.520 ;
        RECT 228.610 -276.995 230.630 -275.735 ;
        RECT 232.985 -276.605 235.495 -274.845 ;
        RECT 274.240 -275.555 277.145 -274.900 ;
        RECT 192.205 -277.945 194.225 -277.185 ;
        RECT 236.160 -277.370 239.065 -276.715 ;
        RECT 274.600 -276.825 276.620 -275.565 ;
        RECT 278.975 -276.435 281.485 -274.675 ;
        RECT 318.010 -275.225 320.915 -274.570 ;
        RECT 318.370 -276.495 320.390 -275.235 ;
        RECT 322.745 -276.105 325.255 -274.345 ;
        RECT 363.775 -275.140 366.680 -274.485 ;
        RECT 282.150 -277.200 285.055 -276.545 ;
        RECT 325.920 -276.870 328.825 -276.215 ;
        RECT 364.135 -276.410 366.155 -275.150 ;
        RECT 368.510 -276.020 371.020 -274.260 ;
        RECT 410.595 -274.950 413.500 -274.295 ;
        RECT 371.685 -276.785 374.590 -276.130 ;
        RECT 410.955 -276.220 412.975 -274.960 ;
        RECT 415.330 -275.830 417.840 -274.070 ;
        RECT 418.505 -276.595 421.410 -275.940 ;
        RECT 236.520 -278.140 238.540 -277.380 ;
        RECT 282.510 -277.970 284.530 -277.210 ;
        RECT 326.280 -277.640 328.300 -276.880 ;
        RECT 372.045 -277.555 374.065 -276.795 ;
        RECT 418.865 -277.365 420.885 -276.605 ;
        RECT -60.580 -279.440 -57.675 -278.785 ;
        RECT -60.220 -280.210 -58.200 -279.450 ;
        RECT -29.510 -280.215 -26.510 -279.455 ;
        RECT -103.055 -281.365 -101.035 -280.605 ;
        RECT -80.170 -281.130 -78.150 -280.370 ;
        RECT -29.455 -280.830 -26.525 -280.230 ;
        RECT -25.320 -280.465 -21.340 -279.705 ;
        RECT -20.795 -280.215 -17.795 -279.455 ;
        RECT -16.010 -280.215 -13.010 -279.455 ;
        RECT -20.740 -280.830 -17.810 -280.230 ;
        RECT -15.955 -280.830 -13.025 -280.230 ;
        RECT -11.820 -280.465 -7.840 -279.705 ;
        RECT -7.295 -280.215 -4.295 -279.455 ;
        RECT -2.885 -280.215 0.115 -279.455 ;
        RECT 10.920 -279.620 12.940 -278.860 ;
        RECT 18.945 -279.630 20.965 -278.870 ;
        RECT -7.240 -280.830 -4.310 -280.230 ;
        RECT -2.830 -280.830 0.100 -280.230 ;
        RECT 10.395 -280.285 13.300 -279.630 ;
        RECT 18.420 -280.295 21.325 -279.640 ;
        RECT 93.715 -279.765 98.260 -278.975 ;
        RECT -103.415 -282.030 -100.510 -281.375 ;
        RECT -106.590 -283.900 -104.080 -282.140 ;
        RECT -97.725 -283.775 -96.195 -282.015 ;
        RECT -96.175 -283.780 -94.645 -282.020 ;
        RECT -94.630 -283.780 -93.100 -282.020 ;
        RECT -92.075 -283.780 -91.035 -282.520 ;
        RECT -88.080 -282.775 -86.060 -281.515 ;
        RECT -80.530 -281.795 -77.625 -281.140 ;
        RECT -88.440 -283.440 -85.535 -282.785 ;
        RECT -83.705 -283.665 -81.195 -281.905 ;
        RECT -29.495 -282.730 -26.565 -282.130 ;
        RECT -25.310 -282.730 -22.380 -282.130 ;
        RECT -29.510 -283.505 -26.510 -282.745 ;
        RECT -25.325 -283.505 -22.325 -282.745 ;
        RECT -21.780 -283.255 -17.800 -282.495 ;
        RECT -15.995 -282.730 -13.065 -282.130 ;
        RECT -11.810 -282.730 -8.880 -282.130 ;
        RECT 1.765 -282.440 2.805 -281.180 ;
        RECT 3.830 -282.440 5.360 -280.680 ;
        RECT 5.375 -282.440 6.905 -280.680 ;
        RECT 6.925 -282.435 8.455 -280.675 ;
        RECT 13.965 -282.155 16.475 -280.395 ;
        RECT 21.990 -282.165 24.500 -280.405 ;
        RECT -16.010 -283.505 -13.010 -282.745 ;
        RECT -11.825 -283.505 -8.825 -282.745 ;
        RECT -8.280 -283.255 -4.300 -282.495 ;
        RECT 14.010 -282.740 16.515 -282.175 ;
        RECT 22.035 -282.750 24.540 -282.185 ;
        RECT 26.575 -282.395 27.615 -281.135 ;
        RECT 28.640 -282.395 30.170 -280.635 ;
        RECT 30.185 -282.395 31.715 -280.635 ;
        RECT 31.735 -282.390 33.265 -280.630 ;
        RECT 34.640 -281.940 35.680 -280.680 ;
        RECT 36.710 -281.940 37.750 -280.680 ;
        RECT 38.520 -281.940 39.560 -280.680 ;
        RECT 39.990 -281.940 41.030 -280.680 ;
        RECT 41.540 -281.940 42.580 -280.680 ;
        RECT 43.085 -281.940 44.125 -280.680 ;
        RECT 94.200 -281.330 96.220 -280.070 ;
        RECT 104.730 -281.810 108.710 -281.050 ;
        RECT 109.255 -281.560 112.255 -280.800 ;
        RECT 113.440 -281.560 116.440 -280.800 ;
        RECT 40.685 -282.825 44.105 -282.085 ;
        RECT 109.310 -282.175 112.240 -281.575 ;
        RECT 113.495 -282.175 116.425 -281.575 ;
        RECT 118.230 -281.810 122.210 -281.050 ;
        RECT 122.755 -281.560 125.755 -280.800 ;
        RECT 126.940 -281.560 129.940 -280.800 ;
        RECT 122.810 -282.175 125.740 -281.575 ;
        RECT 126.995 -282.175 129.925 -281.575 ;
        RECT -106.630 -284.485 -104.125 -283.920 ;
        RECT -83.745 -284.250 -81.240 -283.685 ;
        RECT 1.765 -283.725 8.395 -283.140 ;
        RECT 26.575 -283.680 33.205 -283.095 ;
        RECT 100.330 -284.075 103.260 -283.475 ;
        RECT 104.740 -284.075 107.670 -283.475 ;
        RECT -97.665 -285.065 -91.035 -284.480 ;
        RECT 100.315 -284.850 103.315 -284.090 ;
        RECT 104.725 -284.850 107.725 -284.090 ;
        RECT 108.270 -284.600 112.250 -283.840 ;
        RECT 113.455 -284.075 116.385 -283.475 ;
        RECT 118.240 -284.075 121.170 -283.475 ;
        RECT 113.440 -284.850 116.440 -284.090 ;
        RECT 118.225 -284.850 121.225 -284.090 ;
        RECT 121.770 -284.600 125.750 -283.840 ;
        RECT 126.955 -284.075 129.885 -283.475 ;
        RECT 145.010 -283.690 147.030 -282.930 ;
        RECT 126.940 -284.850 129.940 -284.090 ;
        RECT 144.650 -284.355 147.555 -283.700 ;
        RECT 187.210 -283.745 189.230 -282.985 ;
        RECT 186.850 -284.410 189.755 -283.755 ;
        RECT 231.525 -283.940 233.545 -283.180 ;
        RECT 277.515 -283.770 279.535 -283.010 ;
        RECT 321.285 -283.440 323.305 -282.680 ;
        RECT 367.050 -283.355 369.070 -282.595 ;
        RECT 413.870 -283.165 415.890 -282.405 ;
        RECT -55.225 -286.010 -53.205 -285.250 ;
        RECT -63.135 -287.655 -61.115 -286.395 ;
        RECT -55.585 -286.675 -52.680 -286.020 ;
        RECT 141.475 -286.225 143.985 -284.465 ;
        RECT -63.495 -288.320 -60.590 -287.665 ;
        RECT -58.760 -288.545 -56.250 -286.785 ;
        RECT 141.435 -286.810 143.940 -286.245 ;
        RECT 149.200 -287.655 150.730 -285.895 ;
        RECT 151.390 -287.655 152.430 -285.895 ;
        RECT 158.670 -287.365 159.710 -285.605 ;
        RECT 161.020 -287.365 162.060 -284.605 ;
        RECT 162.135 -287.365 163.175 -284.605 ;
        RECT 163.275 -287.365 164.805 -284.605 ;
        RECT 164.905 -287.365 165.945 -285.605 ;
        RECT 183.675 -286.280 186.185 -284.520 ;
        RECT 231.165 -284.605 234.070 -283.950 ;
        RECT 277.155 -284.435 280.060 -283.780 ;
        RECT 320.925 -284.105 323.830 -283.450 ;
        RECT 366.690 -284.020 369.595 -283.365 ;
        RECT 413.510 -283.830 416.415 -283.175 ;
        RECT 183.635 -286.865 186.140 -286.300 ;
        RECT -58.800 -289.130 -56.295 -288.565 ;
        RECT 116.265 -289.150 130.160 -288.405 ;
        RECT 148.815 -288.610 152.810 -287.940 ;
        RECT 158.340 -288.680 165.965 -287.615 ;
        RECT 191.400 -287.710 192.930 -285.950 ;
        RECT 193.590 -287.710 194.630 -285.950 ;
        RECT 200.870 -287.420 201.910 -285.660 ;
        RECT 203.220 -287.420 204.260 -284.660 ;
        RECT 204.335 -287.420 205.375 -284.660 ;
        RECT 205.475 -287.420 207.005 -284.660 ;
        RECT 207.105 -287.420 208.145 -285.660 ;
        RECT 227.990 -286.475 230.500 -284.715 ;
        RECT 227.950 -287.060 230.455 -286.495 ;
        RECT 191.015 -288.665 195.010 -287.995 ;
        RECT 200.540 -288.735 208.165 -287.670 ;
        RECT 235.715 -287.905 237.245 -286.145 ;
        RECT 237.905 -287.905 238.945 -286.145 ;
        RECT 245.185 -287.615 246.225 -285.855 ;
        RECT 247.535 -287.615 248.575 -284.855 ;
        RECT 248.650 -287.615 249.690 -284.855 ;
        RECT 249.790 -287.615 251.320 -284.855 ;
        RECT 251.420 -287.615 252.460 -285.855 ;
        RECT 273.980 -286.305 276.490 -284.545 ;
        RECT 273.940 -286.890 276.445 -286.325 ;
        RECT 281.705 -287.735 283.235 -285.975 ;
        RECT 283.895 -287.735 284.935 -285.975 ;
        RECT 291.175 -287.445 292.215 -285.685 ;
        RECT 293.525 -287.445 294.565 -284.685 ;
        RECT 294.640 -287.445 295.680 -284.685 ;
        RECT 295.780 -287.445 297.310 -284.685 ;
        RECT 297.410 -287.445 298.450 -285.685 ;
        RECT 317.750 -285.975 320.260 -284.215 ;
        RECT 317.710 -286.560 320.215 -285.995 ;
        RECT 325.475 -287.405 327.005 -285.645 ;
        RECT 327.665 -287.405 328.705 -285.645 ;
        RECT 334.945 -287.115 335.985 -285.355 ;
        RECT 337.295 -287.115 338.335 -284.355 ;
        RECT 338.410 -287.115 339.450 -284.355 ;
        RECT 339.550 -287.115 341.080 -284.355 ;
        RECT 341.180 -287.115 342.220 -285.355 ;
        RECT 363.515 -285.890 366.025 -284.130 ;
        RECT 363.475 -286.475 365.980 -285.910 ;
        RECT 371.240 -287.320 372.770 -285.560 ;
        RECT 373.430 -287.320 374.470 -285.560 ;
        RECT 380.710 -287.030 381.750 -285.270 ;
        RECT 383.060 -287.030 384.100 -284.270 ;
        RECT 384.175 -287.030 385.215 -284.270 ;
        RECT 385.315 -287.030 386.845 -284.270 ;
        RECT 386.945 -287.030 387.985 -285.270 ;
        RECT 410.335 -285.700 412.845 -283.940 ;
        RECT 410.295 -286.285 412.800 -285.720 ;
        RECT 418.060 -287.130 419.590 -285.370 ;
        RECT 420.250 -287.130 421.290 -285.370 ;
        RECT 427.530 -286.840 428.570 -285.080 ;
        RECT 429.880 -286.840 430.920 -284.080 ;
        RECT 430.995 -286.840 432.035 -284.080 ;
        RECT 432.135 -286.840 433.665 -284.080 ;
        RECT 433.765 -286.840 434.805 -285.080 ;
        RECT 235.330 -288.860 239.325 -288.190 ;
        RECT 244.855 -288.930 252.480 -287.865 ;
        RECT 281.320 -288.690 285.315 -288.020 ;
        RECT 290.845 -288.760 298.470 -287.695 ;
        RECT 325.090 -288.360 329.085 -287.690 ;
        RECT 334.615 -288.430 342.240 -287.365 ;
        RECT 370.855 -288.275 374.850 -287.605 ;
        RECT 380.380 -288.345 388.005 -287.280 ;
        RECT 417.675 -288.085 421.670 -287.415 ;
        RECT 427.200 -288.155 434.825 -287.090 ;
        RECT -68.880 -292.660 -65.880 -291.900 ;
        RECT -64.695 -292.660 -61.695 -291.900 ;
        RECT -68.865 -293.275 -65.935 -292.675 ;
        RECT -64.680 -293.275 -61.750 -292.675 ;
        RECT -61.150 -292.910 -57.170 -292.150 ;
        RECT -55.380 -292.660 -52.380 -291.900 ;
        RECT -51.195 -292.660 -48.195 -291.900 ;
        RECT -55.365 -293.275 -52.435 -292.675 ;
        RECT -51.180 -293.275 -48.250 -292.675 ;
        RECT -47.650 -292.910 -43.670 -292.150 ;
        RECT 93.570 -292.885 96.815 -292.180 ;
        RECT 98.300 -292.885 101.545 -292.180 ;
        RECT 103.055 -292.550 109.685 -291.965 ;
        RECT -29.510 -293.995 -26.510 -293.235 ;
        RECT -25.325 -293.995 -22.325 -293.235 ;
        RECT -81.360 -295.320 -77.365 -294.650 ;
        RECT -68.825 -295.175 -65.895 -294.575 ;
        RECT -88.740 -297.015 -86.235 -296.450 ;
        RECT -99.745 -299.790 -98.215 -298.530 ;
        RECT -95.220 -299.795 -93.690 -298.535 ;
        RECT -88.700 -298.795 -86.190 -297.035 ;
        RECT -80.975 -297.365 -79.445 -295.605 ;
        RECT -78.785 -297.365 -77.745 -295.605 ;
        RECT -68.880 -295.950 -65.880 -295.190 ;
        RECT -64.690 -295.700 -60.710 -294.940 ;
        RECT -60.110 -295.175 -57.180 -294.575 ;
        RECT -55.325 -295.175 -52.395 -294.575 ;
        RECT -60.165 -295.950 -57.165 -295.190 ;
        RECT -55.380 -295.950 -52.380 -295.190 ;
        RECT -51.190 -295.700 -47.210 -294.940 ;
        RECT -46.610 -295.175 -43.680 -294.575 ;
        RECT -42.200 -295.175 -39.270 -294.575 ;
        RECT -29.495 -294.610 -26.565 -294.010 ;
        RECT -25.310 -294.610 -22.380 -294.010 ;
        RECT -21.780 -294.245 -17.800 -293.485 ;
        RECT -16.010 -293.995 -13.010 -293.235 ;
        RECT -11.825 -293.995 -8.825 -293.235 ;
        RECT -15.995 -294.610 -13.065 -294.010 ;
        RECT -11.810 -294.610 -8.880 -294.010 ;
        RECT -8.280 -294.245 -4.300 -293.485 ;
        RECT 1.765 -293.600 8.395 -293.015 ;
        RECT 26.575 -293.645 33.205 -293.060 ;
        RECT -46.665 -295.950 -43.665 -295.190 ;
        RECT -42.255 -295.950 -39.255 -295.190 ;
        RECT -37.010 -296.405 -35.970 -294.645 ;
        RECT -35.310 -296.405 -33.780 -294.645 ;
        RECT 1.765 -295.560 2.805 -294.300 ;
        RECT -29.455 -296.510 -26.525 -295.910 ;
        RECT -37.390 -297.360 -33.395 -296.690 ;
        RECT -29.510 -297.285 -26.510 -296.525 ;
        RECT -25.320 -297.035 -21.340 -296.275 ;
        RECT -20.740 -296.510 -17.810 -295.910 ;
        RECT -15.955 -296.510 -13.025 -295.910 ;
        RECT -20.795 -297.285 -17.795 -296.525 ;
        RECT -16.010 -297.285 -13.010 -296.525 ;
        RECT -11.820 -297.035 -7.840 -296.275 ;
        RECT -7.240 -296.510 -4.310 -295.910 ;
        RECT -2.830 -296.510 0.100 -295.910 ;
        RECT 3.830 -296.060 5.360 -294.300 ;
        RECT 5.375 -296.060 6.905 -294.300 ;
        RECT 6.925 -296.065 8.455 -294.305 ;
        RECT 14.010 -294.565 16.515 -294.000 ;
        RECT 22.035 -294.555 24.540 -293.990 ;
        RECT 13.965 -296.345 16.475 -294.585 ;
        RECT 21.990 -296.335 24.500 -294.575 ;
        RECT 26.575 -295.605 27.615 -294.345 ;
        RECT 28.640 -296.105 30.170 -294.345 ;
        RECT 30.185 -296.105 31.715 -294.345 ;
        RECT 31.735 -296.110 33.265 -294.350 ;
        RECT 40.685 -294.655 44.105 -293.915 ;
        RECT 94.175 -294.420 95.705 -293.160 ;
        RECT 98.905 -294.420 100.435 -293.160 ;
        RECT 34.640 -296.060 35.680 -294.800 ;
        RECT 36.710 -296.060 37.750 -294.800 ;
        RECT 38.520 -296.060 39.560 -294.800 ;
        RECT 39.990 -296.060 41.030 -294.800 ;
        RECT 41.540 -296.060 42.580 -294.800 ;
        RECT 43.085 -296.060 44.125 -294.800 ;
        RECT 102.995 -295.015 104.525 -293.255 ;
        RECT 104.545 -295.010 106.075 -293.250 ;
        RECT 106.090 -295.010 107.620 -293.250 ;
        RECT 108.645 -294.510 109.685 -293.250 ;
        RECT 112.540 -293.780 113.580 -292.520 ;
        RECT 113.590 -293.780 114.630 -292.520 ;
        RECT 116.690 -293.235 117.730 -289.475 ;
        RECT 118.690 -293.235 119.730 -289.475 ;
        RECT 121.690 -293.235 122.730 -289.475 ;
        RECT 123.690 -293.235 124.730 -289.475 ;
        RECT 126.690 -293.235 127.730 -289.475 ;
        RECT 128.690 -293.235 129.730 -289.475 ;
        RECT 146.390 -291.840 148.895 -291.275 ;
        RECT 141.695 -292.740 144.600 -292.085 ;
        RECT 142.055 -294.010 144.075 -292.750 ;
        RECT 146.430 -293.620 148.940 -291.860 ;
        RECT 164.730 -291.995 167.235 -291.430 ;
        RECT 188.590 -291.895 191.095 -291.330 ;
        RECT 160.035 -292.895 162.940 -292.240 ;
        RECT 112.435 -294.725 115.090 -294.060 ;
        RECT 149.605 -294.385 152.510 -293.730 ;
        RECT 160.395 -294.165 162.415 -292.905 ;
        RECT 164.770 -293.775 167.280 -292.015 ;
        RECT 183.895 -292.795 186.800 -292.140 ;
        RECT 112.305 -295.340 115.235 -294.740 ;
        RECT 149.965 -295.155 151.985 -294.395 ;
        RECT 167.945 -294.540 170.850 -293.885 ;
        RECT 184.255 -294.065 186.275 -292.805 ;
        RECT 188.630 -293.675 191.140 -291.915 ;
        RECT 206.930 -292.050 209.435 -291.485 ;
        RECT 202.235 -292.950 205.140 -292.295 ;
        RECT 191.805 -294.440 194.710 -293.785 ;
        RECT 202.595 -294.220 204.615 -292.960 ;
        RECT 206.970 -293.830 209.480 -292.070 ;
        RECT 232.905 -292.090 235.410 -291.525 ;
        RECT 228.210 -292.990 231.115 -292.335 ;
        RECT 168.305 -295.310 170.325 -294.550 ;
        RECT 192.165 -295.210 194.185 -294.450 ;
        RECT 210.145 -294.595 213.050 -293.940 ;
        RECT 228.570 -294.260 230.590 -293.000 ;
        RECT 232.945 -293.870 235.455 -292.110 ;
        RECT 251.245 -292.245 253.750 -291.680 ;
        RECT 278.895 -291.920 281.400 -291.355 ;
        RECT 246.550 -293.145 249.455 -292.490 ;
        RECT 112.290 -296.115 115.290 -295.355 ;
        RECT 210.505 -295.365 212.525 -294.605 ;
        RECT 236.120 -294.635 239.025 -293.980 ;
        RECT 246.910 -294.415 248.930 -293.155 ;
        RECT 251.285 -294.025 253.795 -292.265 ;
        RECT 274.200 -292.820 277.105 -292.165 ;
        RECT 274.560 -294.090 276.580 -292.830 ;
        RECT 278.935 -293.700 281.445 -291.940 ;
        RECT 297.235 -292.075 299.740 -291.510 ;
        RECT 322.665 -291.590 325.170 -291.025 ;
        RECT 292.540 -292.975 295.445 -292.320 ;
        RECT 236.480 -295.405 238.500 -294.645 ;
        RECT 254.460 -294.790 257.365 -294.135 ;
        RECT 282.110 -294.465 285.015 -293.810 ;
        RECT 292.900 -294.245 294.920 -292.985 ;
        RECT 297.275 -293.855 299.785 -292.095 ;
        RECT 317.970 -292.490 320.875 -291.835 ;
        RECT 318.330 -293.760 320.350 -292.500 ;
        RECT 322.705 -293.370 325.215 -291.610 ;
        RECT 341.005 -291.745 343.510 -291.180 ;
        RECT 368.430 -291.505 370.935 -290.940 ;
        RECT 336.310 -292.645 339.215 -291.990 ;
        RECT 254.820 -295.560 256.840 -294.800 ;
        RECT 282.470 -295.235 284.490 -294.475 ;
        RECT 300.450 -294.620 303.355 -293.965 ;
        RECT 325.880 -294.135 328.785 -293.480 ;
        RECT 336.670 -293.915 338.690 -292.655 ;
        RECT 341.045 -293.525 343.555 -291.765 ;
        RECT 363.735 -292.405 366.640 -291.750 ;
        RECT 300.810 -295.390 302.830 -294.630 ;
        RECT 326.240 -294.905 328.260 -294.145 ;
        RECT 344.220 -294.290 347.125 -293.635 ;
        RECT 364.095 -293.675 366.115 -292.415 ;
        RECT 368.470 -293.285 370.980 -291.525 ;
        RECT 386.770 -291.660 389.275 -291.095 ;
        RECT 415.250 -291.315 417.755 -290.750 ;
        RECT 382.075 -292.560 384.980 -291.905 ;
        RECT 371.645 -294.050 374.550 -293.395 ;
        RECT 382.435 -293.830 384.455 -292.570 ;
        RECT 386.810 -293.440 389.320 -291.680 ;
        RECT 410.555 -292.215 413.460 -291.560 ;
        RECT 410.915 -293.485 412.935 -292.225 ;
        RECT 415.290 -293.095 417.800 -291.335 ;
        RECT 433.590 -291.470 436.095 -290.905 ;
        RECT 428.895 -292.370 431.800 -291.715 ;
        RECT 344.580 -295.060 346.600 -294.300 ;
        RECT 372.005 -294.820 374.025 -294.060 ;
        RECT 389.985 -294.205 392.890 -293.550 ;
        RECT 418.465 -293.860 421.370 -293.205 ;
        RECT 429.255 -293.640 431.275 -292.380 ;
        RECT 433.630 -293.250 436.140 -291.490 ;
        RECT 390.345 -294.975 392.365 -294.215 ;
        RECT 418.825 -294.630 420.845 -293.870 ;
        RECT 436.805 -294.015 439.710 -293.360 ;
        RECT 437.165 -294.785 439.185 -294.025 ;
        RECT -7.295 -297.285 -4.295 -296.525 ;
        RECT -2.885 -297.285 0.115 -296.525 ;
        RECT 10.395 -297.110 13.300 -296.455 ;
        RECT 18.420 -297.100 21.325 -296.445 ;
        RECT 10.920 -297.880 12.940 -297.120 ;
        RECT 18.945 -297.870 20.965 -297.110 ;
        RECT -85.525 -299.560 -82.620 -298.905 ;
        RECT -105.775 -301.505 -103.755 -300.245 ;
        RECT -100.350 -300.770 -97.105 -300.065 ;
        RECT -95.825 -300.775 -92.580 -300.070 ;
        RECT -85.165 -300.330 -83.145 -299.570 ;
        RECT 144.970 -300.955 146.990 -300.195 ;
        RECT 144.610 -301.620 147.515 -300.965 ;
        RECT 163.310 -301.110 165.330 -300.350 ;
        RECT 187.170 -301.010 189.190 -300.250 ;
        RECT -106.260 -302.600 -101.715 -301.810 ;
        RECT 141.435 -303.490 143.945 -301.730 ;
        RECT 162.950 -301.775 165.855 -301.120 ;
        RECT 186.810 -301.675 189.715 -301.020 ;
        RECT 205.510 -301.165 207.530 -300.405 ;
        RECT 59.675 -304.340 62.675 -303.580 ;
        RECT 64.085 -304.340 67.085 -303.580 ;
        RECT -107.460 -305.275 -100.830 -304.690 ;
        RECT 59.690 -304.955 62.620 -304.355 ;
        RECT 64.100 -304.955 67.030 -304.355 ;
        RECT 67.630 -304.590 71.610 -303.830 ;
        RECT 72.800 -304.340 75.800 -303.580 ;
        RECT 77.585 -304.340 80.585 -303.580 ;
        RECT 72.815 -304.955 75.745 -304.355 ;
        RECT 77.600 -304.955 80.530 -304.355 ;
        RECT 81.130 -304.590 85.110 -303.830 ;
        RECT 86.300 -304.340 89.300 -303.580 ;
        RECT 141.395 -304.075 143.900 -303.510 ;
        RECT 86.315 -304.955 89.245 -304.355 ;
        RECT 149.160 -304.920 150.690 -303.160 ;
        RECT 151.350 -304.920 152.390 -303.160 ;
        RECT 159.775 -303.645 162.285 -301.885 ;
        RECT 159.735 -304.230 162.240 -303.665 ;
        RECT 167.500 -305.075 169.030 -303.315 ;
        RECT 169.690 -305.075 170.730 -303.315 ;
        RECT 183.635 -303.545 186.145 -301.785 ;
        RECT 205.150 -301.830 208.055 -301.175 ;
        RECT 231.485 -301.205 233.505 -300.445 ;
        RECT 231.125 -301.870 234.030 -301.215 ;
        RECT 249.825 -301.360 251.845 -300.600 ;
        RECT 277.475 -301.035 279.495 -300.275 ;
        RECT 183.595 -304.130 186.100 -303.565 ;
        RECT 191.360 -304.975 192.890 -303.215 ;
        RECT 193.550 -304.975 194.590 -303.215 ;
        RECT 201.975 -303.700 204.485 -301.940 ;
        RECT 201.935 -304.285 204.440 -303.720 ;
        RECT 209.700 -305.130 211.230 -303.370 ;
        RECT 211.890 -305.130 212.930 -303.370 ;
        RECT 227.950 -303.740 230.460 -301.980 ;
        RECT 249.465 -302.025 252.370 -301.370 ;
        RECT 277.115 -301.700 280.020 -301.045 ;
        RECT 295.815 -301.190 297.835 -300.430 ;
        RECT 321.245 -300.705 323.265 -299.945 ;
        RECT 227.910 -304.325 230.415 -303.760 ;
        RECT 235.675 -305.170 237.205 -303.410 ;
        RECT 237.865 -305.170 238.905 -303.410 ;
        RECT 246.290 -303.895 248.800 -302.135 ;
        RECT 246.250 -304.480 248.755 -303.915 ;
        RECT -107.460 -307.235 -106.420 -305.975 ;
        RECT -105.395 -307.735 -103.865 -305.975 ;
        RECT -103.850 -307.735 -102.320 -305.975 ;
        RECT -102.300 -307.740 -100.770 -305.980 ;
        RECT -80.170 -306.130 -78.150 -305.370 ;
        RECT -24.365 -305.910 -20.945 -305.170 ;
        RECT -11.865 -305.910 -8.445 -305.170 ;
        RECT 0.635 -305.910 4.055 -305.170 ;
        RECT 13.135 -305.910 16.555 -305.170 ;
        RECT 25.635 -305.910 29.055 -305.170 ;
        RECT 40.635 -305.910 44.055 -305.170 ;
        RECT 148.775 -305.875 152.770 -305.205 ;
        RECT 167.115 -306.030 171.110 -305.360 ;
        RECT 190.975 -305.930 194.970 -305.260 ;
        RECT 254.015 -305.325 255.545 -303.565 ;
        RECT 256.205 -305.325 257.245 -303.565 ;
        RECT 273.940 -303.570 276.450 -301.810 ;
        RECT 295.455 -301.855 298.360 -301.200 ;
        RECT 320.885 -301.370 323.790 -300.715 ;
        RECT 339.585 -300.860 341.605 -300.100 ;
        RECT 367.010 -300.620 369.030 -299.860 ;
        RECT 273.900 -304.155 276.405 -303.590 ;
        RECT 281.665 -305.000 283.195 -303.240 ;
        RECT 283.855 -305.000 284.895 -303.240 ;
        RECT 292.280 -303.725 294.790 -301.965 ;
        RECT 317.710 -303.240 320.220 -301.480 ;
        RECT 339.225 -301.525 342.130 -300.870 ;
        RECT 366.650 -301.285 369.555 -300.630 ;
        RECT 385.350 -300.775 387.370 -300.015 ;
        RECT 413.830 -300.430 415.850 -299.670 ;
        RECT 292.240 -304.310 294.745 -303.745 ;
        RECT 300.005 -305.155 301.535 -303.395 ;
        RECT 302.195 -305.155 303.235 -303.395 ;
        RECT 317.670 -303.825 320.175 -303.260 ;
        RECT 325.435 -304.670 326.965 -302.910 ;
        RECT 327.625 -304.670 328.665 -302.910 ;
        RECT 336.050 -303.395 338.560 -301.635 ;
        RECT 336.010 -303.980 338.515 -303.415 ;
        RECT 343.775 -304.825 345.305 -303.065 ;
        RECT 345.965 -304.825 347.005 -303.065 ;
        RECT 363.475 -303.155 365.985 -301.395 ;
        RECT 384.990 -301.440 387.895 -300.785 ;
        RECT 413.470 -301.095 416.375 -300.440 ;
        RECT 432.170 -300.585 434.190 -299.825 ;
        RECT 363.435 -303.740 365.940 -303.175 ;
        RECT 371.200 -304.585 372.730 -302.825 ;
        RECT 373.390 -304.585 374.430 -302.825 ;
        RECT 381.815 -303.310 384.325 -301.550 ;
        RECT 410.295 -302.965 412.805 -301.205 ;
        RECT 431.810 -301.250 434.715 -300.595 ;
        RECT 381.775 -303.895 384.280 -303.330 ;
        RECT 389.540 -304.740 391.070 -302.980 ;
        RECT 391.730 -304.740 392.770 -302.980 ;
        RECT 410.255 -303.550 412.760 -302.985 ;
        RECT 418.020 -304.395 419.550 -302.635 ;
        RECT 420.210 -304.395 421.250 -302.635 ;
        RECT 428.635 -303.120 431.145 -301.360 ;
        RECT 428.595 -303.705 431.100 -303.140 ;
        RECT 436.360 -304.550 437.890 -302.790 ;
        RECT 438.550 -304.550 439.590 -302.790 ;
        RECT -88.080 -307.775 -86.060 -306.515 ;
        RECT -80.530 -306.795 -77.625 -306.140 ;
        RECT -88.440 -308.440 -85.535 -307.785 ;
        RECT -83.705 -308.665 -81.195 -306.905 ;
        RECT -30.410 -307.315 -29.370 -306.055 ;
        RECT -28.340 -307.315 -27.300 -306.055 ;
        RECT -26.530 -307.315 -25.490 -306.055 ;
        RECT -25.060 -307.315 -24.020 -306.055 ;
        RECT -23.510 -307.315 -22.470 -306.055 ;
        RECT -21.965 -307.315 -20.925 -306.055 ;
        RECT -17.910 -307.315 -16.870 -306.055 ;
        RECT -15.840 -307.315 -14.800 -306.055 ;
        RECT -14.030 -307.315 -12.990 -306.055 ;
        RECT -12.560 -307.315 -11.520 -306.055 ;
        RECT -11.010 -307.315 -9.970 -306.055 ;
        RECT -9.465 -307.315 -8.425 -306.055 ;
        RECT -5.410 -307.315 -4.370 -306.055 ;
        RECT -3.340 -307.315 -2.300 -306.055 ;
        RECT -1.530 -307.315 -0.490 -306.055 ;
        RECT -0.060 -307.315 0.980 -306.055 ;
        RECT 1.490 -307.315 2.530 -306.055 ;
        RECT 3.035 -307.315 4.075 -306.055 ;
        RECT 7.090 -307.315 8.130 -306.055 ;
        RECT 9.160 -307.315 10.200 -306.055 ;
        RECT 10.970 -307.315 12.010 -306.055 ;
        RECT 12.440 -307.315 13.480 -306.055 ;
        RECT 13.990 -307.315 15.030 -306.055 ;
        RECT 15.535 -307.315 16.575 -306.055 ;
        RECT 19.590 -307.315 20.630 -306.055 ;
        RECT 21.660 -307.315 22.700 -306.055 ;
        RECT 23.470 -307.315 24.510 -306.055 ;
        RECT 24.940 -307.315 25.980 -306.055 ;
        RECT 26.490 -307.315 27.530 -306.055 ;
        RECT 28.035 -307.315 29.075 -306.055 ;
        RECT 34.590 -307.315 35.630 -306.055 ;
        RECT 36.660 -307.315 37.700 -306.055 ;
        RECT 38.470 -307.315 39.510 -306.055 ;
        RECT 39.940 -307.315 40.980 -306.055 ;
        RECT 41.490 -307.315 42.530 -306.055 ;
        RECT 43.035 -307.315 44.075 -306.055 ;
        RECT 209.315 -306.085 213.310 -305.415 ;
        RECT 235.290 -306.125 239.285 -305.455 ;
        RECT 64.090 -307.380 68.070 -306.620 ;
        RECT 68.670 -306.855 71.600 -306.255 ;
        RECT 72.855 -306.855 75.785 -306.255 ;
        RECT 68.615 -307.630 71.615 -306.870 ;
        RECT 72.800 -307.630 75.800 -306.870 ;
        RECT 77.590 -307.380 81.570 -306.620 ;
        RECT 82.170 -306.855 85.100 -306.255 ;
        RECT 86.355 -306.855 89.285 -306.255 ;
        RECT 253.630 -306.280 257.625 -305.610 ;
        RECT 281.280 -305.955 285.275 -305.285 ;
        RECT 299.620 -306.110 303.615 -305.440 ;
        RECT 325.050 -305.625 329.045 -304.955 ;
        RECT 343.390 -305.780 347.385 -305.110 ;
        RECT 370.815 -305.540 374.810 -304.870 ;
        RECT 389.155 -305.695 393.150 -305.025 ;
        RECT 417.635 -305.350 421.630 -304.680 ;
        RECT 435.975 -305.505 439.970 -304.835 ;
        RECT 82.115 -307.630 85.115 -306.870 ;
        RECT 86.300 -307.630 89.300 -306.870 ;
        RECT -83.745 -309.250 -81.240 -308.685 ;
      LAYER li1 ;
        RECT -62.330 603.475 -60.615 605.270 ;
        RECT -61.580 599.415 -61.365 603.475 ;
        RECT -60.850 600.735 -60.490 600.855 ;
        RECT -60.850 600.385 -53.455 600.735 ;
        RECT -60.850 600.330 -60.490 600.385 ;
        RECT -61.580 599.375 -60.145 599.415 ;
        RECT -61.580 599.205 -57.175 599.375 ;
        RECT -61.580 599.200 -60.145 599.205 ;
        RECT -61.580 598.990 -61.365 599.200 ;
        RECT -53.805 599.045 -53.455 600.385 ;
        RECT -61.780 598.960 -61.365 598.990 ;
        RECT -63.275 598.790 -61.365 598.960 ;
        RECT -61.780 598.770 -61.365 598.790 ;
        RECT -61.565 598.530 -61.365 598.770 ;
        RECT -60.915 598.340 -60.640 599.030 ;
        RECT -54.665 598.875 -53.455 599.045 ;
        RECT -53.510 598.385 -52.970 598.555 ;
        RECT -61.465 598.125 -60.385 598.340 ;
        RECT -57.225 598.315 -56.835 598.345 ;
        RECT -60.215 598.145 -56.835 598.315 ;
        RECT -57.225 598.135 -56.835 598.145 ;
        RECT -61.465 596.795 -61.265 598.125 ;
        RECT -60.580 597.845 -60.385 598.125 ;
        RECT -60.580 597.825 -60.115 597.845 ;
        RECT -61.025 596.915 -60.750 597.690 ;
        RECT -60.580 597.655 -57.175 597.825 ;
        RECT -60.580 597.635 -60.115 597.655 ;
        RECT -60.570 597.335 -60.125 597.360 ;
        RECT -57.005 597.355 -56.835 598.135 ;
        RECT -54.665 597.895 -54.125 598.065 ;
        RECT -53.510 597.405 -52.970 597.575 ;
        RECT -57.215 597.335 -56.835 597.355 ;
        RECT -60.570 597.165 -56.835 597.335 ;
        RECT -60.570 597.150 -60.125 597.165 ;
        RECT -61.815 596.770 -61.265 596.795 ;
        RECT -63.275 596.600 -61.265 596.770 ;
        RECT -61.815 596.570 -61.265 596.600 ;
        RECT -61.565 595.565 -61.290 596.340 ;
        RECT -61.505 595.380 -61.335 595.565 ;
        RECT -60.980 595.240 -60.800 596.915 ;
        RECT -60.570 596.300 -60.390 597.150 ;
        RECT -57.215 597.145 -56.835 597.165 ;
        RECT -54.665 596.915 -54.125 597.085 ;
        RECT -53.955 596.325 -53.655 596.690 ;
        RECT -60.570 596.280 -60.095 596.300 ;
        RECT -60.570 596.110 -57.175 596.280 ;
        RECT -60.570 596.090 -60.095 596.110 ;
        RECT -53.890 596.020 -53.685 596.325 ;
        RECT -53.890 595.965 -52.790 596.020 ;
        RECT -53.890 595.825 -52.750 595.965 ;
        RECT -53.750 595.715 -52.750 595.825 ;
        RECT -58.825 595.240 -58.475 595.270 ;
        RECT -60.990 594.890 -58.475 595.240 ;
        RECT -52.940 595.020 -52.750 595.715 ;
        RECT -52.515 595.280 -52.160 595.650 ;
        RECT -51.975 595.340 -50.435 595.510 ;
        RECT -58.825 594.050 -58.475 594.890 ;
        RECT -54.660 594.850 -52.750 595.020 ;
        RECT -58.825 593.880 -57.615 594.050 ;
        RECT -52.940 594.040 -52.750 594.850 ;
        RECT -54.660 593.870 -52.750 594.040 ;
        RECT -59.310 593.390 -58.770 593.560 ;
        RECT -58.155 592.900 -57.615 593.070 ;
        RECT -52.905 592.955 -52.635 593.630 ;
        RECT -52.385 593.575 -52.190 595.280 ;
        RECT -48.465 595.275 -43.610 595.465 ;
        RECT -51.975 594.850 -50.435 595.020 ;
        RECT -51.975 594.360 -50.435 594.530 ;
        RECT -52.385 593.225 -52.185 593.575 ;
        RECT -51.975 593.380 -50.435 593.550 ;
        RECT -52.395 593.220 -52.185 593.225 ;
        RECT -52.875 592.855 -52.675 592.955 ;
        RECT -59.310 592.410 -58.770 592.580 ;
        RECT -58.155 591.920 -57.615 592.090 ;
        RECT -52.865 591.820 -52.685 592.855 ;
        RECT -58.625 591.330 -58.325 591.695 ;
        RECT -58.595 591.025 -58.390 591.330 ;
        RECT -59.490 590.970 -58.390 591.025 ;
        RECT -59.530 590.830 -58.390 590.970 ;
        RECT -54.015 590.965 -52.975 591.135 ;
        RECT -59.530 590.720 -58.530 590.830 ;
        RECT -61.845 590.345 -60.305 590.515 ;
        RECT -60.120 590.285 -59.765 590.655 ;
        RECT -61.845 589.855 -60.305 590.025 ;
        RECT -61.845 589.365 -60.305 589.535 ;
        RECT -60.090 588.580 -59.895 590.285 ;
        RECT -59.530 590.025 -59.340 590.720 ;
        RECT -52.395 590.645 -52.195 593.220 ;
        RECT -52.395 590.480 -51.325 590.645 ;
        RECT -52.365 590.475 -51.325 590.480 ;
        RECT -59.530 589.855 -57.620 590.025 ;
        RECT -54.015 589.985 -52.975 590.155 ;
        RECT -59.530 589.045 -59.340 589.855 ;
        RECT -52.365 589.495 -51.325 589.665 ;
        RECT -59.530 588.875 -57.620 589.045 ;
        RECT -54.015 589.005 -52.975 589.175 ;
        RECT -61.845 588.385 -60.305 588.555 ;
        RECT -60.095 588.230 -59.895 588.580 ;
        RECT -52.805 588.415 -52.505 588.780 ;
        RECT -60.095 588.225 -59.885 588.230 ;
        RECT -60.085 587.095 -59.885 588.225 ;
        RECT -52.740 588.195 -52.535 588.415 ;
        RECT -52.825 588.060 -52.075 588.195 ;
        RECT -53.075 587.680 -52.075 588.060 ;
        RECT -52.825 587.545 -52.075 587.680 ;
        RECT -52.585 585.400 -52.205 587.545 ;
        RECT -50.625 586.720 -50.355 586.780 ;
        RECT -48.465 586.720 -48.275 595.275 ;
        RECT -43.800 594.195 -43.610 595.275 ;
        RECT -44.050 594.175 -40.960 594.195 ;
        RECT -45.565 594.005 -40.960 594.175 ;
        RECT -43.060 593.430 -42.765 593.700 ;
        RECT -43.020 593.170 -42.850 593.430 ;
        RECT -42.275 593.170 -42.005 593.830 ;
        RECT -41.145 593.695 -40.960 594.005 ;
        RECT -41.145 593.685 -40.495 593.695 ;
        RECT -41.145 593.515 -39.045 593.685 ;
        RECT -41.145 593.510 -40.495 593.515 ;
        RECT -43.045 593.035 -41.615 593.170 ;
        RECT -45.565 593.000 -41.615 593.035 ;
        RECT -45.565 592.865 -42.875 593.000 ;
        RECT -43.045 592.860 -42.875 592.865 ;
        RECT -45.565 592.375 -43.025 592.545 ;
        RECT -42.690 592.540 -42.000 592.810 ;
        RECT -41.785 592.545 -41.615 593.000 ;
        RECT -41.785 592.375 -39.045 592.545 ;
        RECT -42.180 591.490 -41.910 592.180 ;
        RECT -45.565 590.745 -42.870 590.915 ;
        RECT -43.045 590.290 -42.870 590.745 ;
        RECT -42.615 590.615 -42.345 591.305 ;
        RECT -42.135 590.915 -41.965 591.490 ;
        RECT -42.135 590.745 -39.045 590.915 ;
        RECT -45.565 590.120 -42.870 590.290 ;
        RECT -42.135 590.285 -41.965 590.745 ;
        RECT -42.700 590.115 -41.965 590.285 ;
        RECT -39.060 590.265 -38.695 590.270 ;
        RECT -42.700 589.800 -42.530 590.115 ;
        RECT -41.585 590.095 -38.695 590.265 ;
        RECT -45.565 589.630 -42.530 589.800 ;
        RECT -42.340 589.775 -41.550 589.780 ;
        RECT -42.340 589.605 -39.045 589.775 ;
        RECT -42.340 589.590 -41.550 589.605 ;
        RECT -43.380 589.105 -42.690 589.135 ;
        RECT -42.340 589.105 -42.150 589.590 ;
        RECT -38.865 589.285 -38.695 590.095 ;
        RECT -41.585 589.115 -38.695 589.285 ;
        RECT -39.065 589.110 -38.695 589.115 ;
        RECT -43.380 588.915 -42.150 589.105 ;
        RECT -43.380 588.865 -42.690 588.915 ;
        RECT -42.340 587.940 -42.150 588.915 ;
        RECT -38.865 588.865 -38.695 589.110 ;
        RECT -45.565 587.770 -42.150 587.940 ;
        RECT -41.975 588.665 -38.695 588.865 ;
        RECT -41.975 587.940 -41.775 588.665 ;
        RECT -41.975 587.770 -39.045 587.940 ;
        RECT -41.975 587.765 -41.545 587.770 ;
        RECT -43.295 586.865 -43.025 587.555 ;
        RECT -50.625 586.530 -48.275 586.720 ;
        RECT -50.625 586.415 -50.355 586.530 ;
        RECT -44.270 586.175 -43.875 586.235 ;
        RECT -43.240 586.175 -43.070 586.865 ;
        RECT -42.615 586.585 -42.345 587.275 ;
        RECT -44.270 585.840 -43.070 586.175 ;
        RECT -43.920 585.815 -43.070 585.840 ;
        RECT -52.585 585.020 -48.305 585.400 ;
        RECT -61.425 584.595 -59.965 584.810 ;
        RECT -61.425 581.075 -61.210 584.595 ;
        RECT -60.180 583.600 -59.965 584.595 ;
        RECT -50.090 583.600 -49.665 583.730 ;
        RECT -60.180 583.385 -49.665 583.600 ;
        RECT -50.090 583.270 -49.665 583.385 ;
        RECT -60.695 582.395 -60.335 582.515 ;
        RECT -60.695 582.045 -53.300 582.395 ;
        RECT -60.695 581.990 -60.335 582.045 ;
        RECT -61.425 581.035 -59.990 581.075 ;
        RECT -61.425 580.865 -57.020 581.035 ;
        RECT -61.425 580.860 -59.990 580.865 ;
        RECT -61.425 580.650 -61.210 580.860 ;
        RECT -53.650 580.705 -53.300 582.045 ;
        RECT -61.625 580.620 -61.210 580.650 ;
        RECT -63.120 580.450 -61.210 580.620 ;
        RECT -61.625 580.430 -61.210 580.450 ;
        RECT -61.410 580.190 -61.210 580.430 ;
        RECT -60.760 580.000 -60.485 580.690 ;
        RECT -54.510 580.535 -53.300 580.705 ;
        RECT -53.355 580.045 -52.815 580.215 ;
        RECT -61.310 579.785 -60.230 580.000 ;
        RECT -57.070 579.975 -56.680 580.005 ;
        RECT -60.060 579.805 -56.680 579.975 ;
        RECT -57.070 579.795 -56.680 579.805 ;
        RECT -61.310 578.455 -61.110 579.785 ;
        RECT -60.425 579.505 -60.230 579.785 ;
        RECT -60.425 579.485 -59.960 579.505 ;
        RECT -60.870 578.575 -60.595 579.350 ;
        RECT -60.425 579.315 -57.020 579.485 ;
        RECT -60.425 579.295 -59.960 579.315 ;
        RECT -60.415 578.995 -59.970 579.020 ;
        RECT -56.850 579.015 -56.680 579.795 ;
        RECT -54.510 579.555 -53.970 579.725 ;
        RECT -53.355 579.065 -52.815 579.235 ;
        RECT -57.060 578.995 -56.680 579.015 ;
        RECT -60.415 578.825 -56.680 578.995 ;
        RECT -60.415 578.810 -59.970 578.825 ;
        RECT -61.660 578.430 -61.110 578.455 ;
        RECT -63.120 578.260 -61.110 578.430 ;
        RECT -61.660 578.230 -61.110 578.260 ;
        RECT -61.410 577.225 -61.135 578.000 ;
        RECT -61.350 577.040 -61.180 577.225 ;
        RECT -60.825 576.900 -60.645 578.575 ;
        RECT -60.415 577.960 -60.235 578.810 ;
        RECT -57.060 578.805 -56.680 578.825 ;
        RECT -54.510 578.575 -53.970 578.745 ;
        RECT -53.800 577.985 -53.500 578.350 ;
        RECT -60.415 577.940 -59.940 577.960 ;
        RECT -60.415 577.770 -57.020 577.940 ;
        RECT -60.415 577.750 -59.940 577.770 ;
        RECT -53.735 577.680 -53.530 577.985 ;
        RECT -53.735 577.625 -52.635 577.680 ;
        RECT -53.735 577.485 -52.595 577.625 ;
        RECT -53.595 577.375 -52.595 577.485 ;
        RECT -58.670 576.900 -58.320 576.930 ;
        RECT -60.835 576.550 -58.320 576.900 ;
        RECT -52.785 576.680 -52.595 577.375 ;
        RECT -52.360 576.940 -52.005 577.310 ;
        RECT -51.820 577.000 -50.280 577.170 ;
        RECT -58.670 575.710 -58.320 576.550 ;
        RECT -54.505 576.510 -52.595 576.680 ;
        RECT -58.670 575.540 -57.460 575.710 ;
        RECT -52.785 575.700 -52.595 576.510 ;
        RECT -54.505 575.530 -52.595 575.700 ;
        RECT -59.155 575.050 -58.615 575.220 ;
        RECT -58.000 574.560 -57.460 574.730 ;
        RECT -52.750 574.615 -52.480 575.290 ;
        RECT -52.230 575.235 -52.035 576.940 ;
        RECT -51.820 576.510 -50.280 576.680 ;
        RECT -51.820 576.020 -50.280 576.190 ;
        RECT -52.230 574.885 -52.030 575.235 ;
        RECT -51.820 575.040 -50.280 575.210 ;
        RECT -52.240 574.880 -52.030 574.885 ;
        RECT -52.720 574.515 -52.520 574.615 ;
        RECT -59.155 574.070 -58.615 574.240 ;
        RECT -58.000 573.580 -57.460 573.750 ;
        RECT -52.710 573.480 -52.530 574.515 ;
        RECT -58.470 572.990 -58.170 573.355 ;
        RECT -58.440 572.685 -58.235 572.990 ;
        RECT -59.335 572.630 -58.235 572.685 ;
        RECT -59.375 572.490 -58.235 572.630 ;
        RECT -53.860 572.625 -52.820 572.795 ;
        RECT -59.375 572.380 -58.375 572.490 ;
        RECT -61.690 572.005 -60.150 572.175 ;
        RECT -59.965 571.945 -59.610 572.315 ;
        RECT -61.690 571.515 -60.150 571.685 ;
        RECT -61.690 571.025 -60.150 571.195 ;
        RECT -59.935 570.240 -59.740 571.945 ;
        RECT -59.375 571.685 -59.185 572.380 ;
        RECT -52.240 572.305 -52.040 574.880 ;
        RECT -52.240 572.140 -51.170 572.305 ;
        RECT -52.210 572.135 -51.170 572.140 ;
        RECT -59.375 571.515 -57.465 571.685 ;
        RECT -53.860 571.645 -52.820 571.815 ;
        RECT -59.375 570.705 -59.185 571.515 ;
        RECT -52.210 571.155 -51.170 571.325 ;
        RECT -59.375 570.535 -57.465 570.705 ;
        RECT -53.860 570.665 -52.820 570.835 ;
        RECT -61.690 570.045 -60.150 570.215 ;
        RECT -59.940 569.890 -59.740 570.240 ;
        RECT -52.650 570.075 -52.350 570.440 ;
        RECT -59.940 569.885 -59.730 569.890 ;
        RECT -59.930 568.755 -59.730 569.885 ;
        RECT -52.585 569.855 -52.380 570.075 ;
        RECT -52.670 569.560 -51.920 569.855 ;
        RECT -52.670 569.230 -49.595 569.560 ;
        RECT -48.685 569.440 -48.305 585.020 ;
        RECT -42.565 584.850 -42.395 586.585 ;
        RECT -44.160 584.635 -42.395 584.850 ;
        RECT -44.160 581.115 -43.945 584.635 ;
        RECT -43.430 582.435 -43.070 582.555 ;
        RECT -43.430 582.085 -36.035 582.435 ;
        RECT -43.430 582.030 -43.070 582.085 ;
        RECT -44.160 581.075 -42.725 581.115 ;
        RECT -44.160 580.905 -39.755 581.075 ;
        RECT -44.160 580.900 -42.725 580.905 ;
        RECT -44.160 580.690 -43.945 580.900 ;
        RECT -36.385 580.745 -36.035 582.085 ;
        RECT -44.360 580.660 -43.945 580.690 ;
        RECT -45.855 580.490 -43.945 580.660 ;
        RECT -44.360 580.470 -43.945 580.490 ;
        RECT -44.145 580.230 -43.945 580.470 ;
        RECT -43.495 580.040 -43.220 580.730 ;
        RECT -37.245 580.575 -36.035 580.745 ;
        RECT -36.090 580.085 -35.550 580.255 ;
        RECT -44.045 579.825 -42.965 580.040 ;
        RECT -39.805 580.015 -39.415 580.045 ;
        RECT -42.795 579.845 -39.415 580.015 ;
        RECT -39.805 579.835 -39.415 579.845 ;
        RECT -44.045 578.495 -43.845 579.825 ;
        RECT -43.160 579.545 -42.965 579.825 ;
        RECT -43.160 579.525 -42.695 579.545 ;
        RECT -43.605 578.615 -43.330 579.390 ;
        RECT -43.160 579.355 -39.755 579.525 ;
        RECT -43.160 579.335 -42.695 579.355 ;
        RECT -43.150 579.035 -42.705 579.060 ;
        RECT -39.585 579.055 -39.415 579.835 ;
        RECT -37.245 579.595 -36.705 579.765 ;
        RECT -36.090 579.105 -35.550 579.275 ;
        RECT -39.795 579.035 -39.415 579.055 ;
        RECT -43.150 578.865 -39.415 579.035 ;
        RECT -43.150 578.850 -42.705 578.865 ;
        RECT -44.395 578.470 -43.845 578.495 ;
        RECT -45.855 578.300 -43.845 578.470 ;
        RECT -44.395 578.270 -43.845 578.300 ;
        RECT -44.145 577.265 -43.870 578.040 ;
        RECT -44.085 577.080 -43.915 577.265 ;
        RECT -43.560 576.940 -43.380 578.615 ;
        RECT -43.150 578.000 -42.970 578.850 ;
        RECT -39.795 578.845 -39.415 578.865 ;
        RECT -37.245 578.615 -36.705 578.785 ;
        RECT -36.535 578.025 -36.235 578.390 ;
        RECT -43.150 577.980 -42.675 578.000 ;
        RECT -43.150 577.810 -39.755 577.980 ;
        RECT -43.150 577.790 -42.675 577.810 ;
        RECT -36.470 577.720 -36.265 578.025 ;
        RECT -36.470 577.665 -35.370 577.720 ;
        RECT -36.470 577.525 -35.330 577.665 ;
        RECT -36.330 577.415 -35.330 577.525 ;
        RECT -41.405 576.940 -41.055 576.970 ;
        RECT -43.570 576.590 -41.055 576.940 ;
        RECT -35.520 576.720 -35.330 577.415 ;
        RECT -35.095 576.980 -34.740 577.350 ;
        RECT -34.555 577.040 -33.015 577.210 ;
        RECT -41.405 575.750 -41.055 576.590 ;
        RECT -37.240 576.550 -35.330 576.720 ;
        RECT -41.405 575.580 -40.195 575.750 ;
        RECT -35.520 575.740 -35.330 576.550 ;
        RECT -37.240 575.570 -35.330 575.740 ;
        RECT -41.890 575.090 -41.350 575.260 ;
        RECT -40.735 574.600 -40.195 574.770 ;
        RECT -35.485 574.655 -35.215 575.330 ;
        RECT -34.965 575.275 -34.770 576.980 ;
        RECT -34.555 576.550 -33.015 576.720 ;
        RECT -34.555 576.060 -33.015 576.230 ;
        RECT -34.965 574.925 -34.765 575.275 ;
        RECT -34.555 575.080 -33.015 575.250 ;
        RECT -34.975 574.920 -34.765 574.925 ;
        RECT -35.455 574.555 -35.255 574.655 ;
        RECT -41.890 574.110 -41.350 574.280 ;
        RECT -40.735 573.620 -40.195 573.790 ;
        RECT -35.445 573.520 -35.265 574.555 ;
        RECT -41.205 573.030 -40.905 573.395 ;
        RECT -41.175 572.725 -40.970 573.030 ;
        RECT -42.070 572.670 -40.970 572.725 ;
        RECT -42.110 572.530 -40.970 572.670 ;
        RECT -36.595 572.665 -35.555 572.835 ;
        RECT -42.110 572.420 -41.110 572.530 ;
        RECT -44.425 572.045 -42.885 572.215 ;
        RECT -42.700 571.985 -42.345 572.355 ;
        RECT -44.425 571.555 -42.885 571.725 ;
        RECT -44.425 571.065 -42.885 571.235 ;
        RECT -42.670 570.280 -42.475 571.985 ;
        RECT -42.110 571.725 -41.920 572.420 ;
        RECT -34.975 572.345 -34.775 574.920 ;
        RECT -34.975 572.180 -33.905 572.345 ;
        RECT -34.945 572.175 -33.905 572.180 ;
        RECT -42.110 571.555 -40.200 571.725 ;
        RECT -36.595 571.685 -35.555 571.855 ;
        RECT -42.110 570.745 -41.920 571.555 ;
        RECT -34.945 571.195 -33.905 571.365 ;
        RECT -42.110 570.575 -40.200 570.745 ;
        RECT -36.595 570.705 -35.555 570.875 ;
        RECT -44.425 570.085 -42.885 570.255 ;
        RECT -42.675 569.930 -42.475 570.280 ;
        RECT -35.385 570.115 -35.085 570.480 ;
        RECT -42.675 569.925 -42.465 569.930 ;
        RECT -48.700 569.230 -47.570 569.440 ;
        RECT -42.665 569.230 -42.465 569.925 ;
        RECT -35.320 569.895 -35.115 570.115 ;
        RECT -35.405 569.245 -34.655 569.895 ;
        RECT -52.670 569.205 -42.465 569.230 ;
        RECT -52.465 569.180 -42.465 569.205 ;
        RECT -49.975 568.850 -42.465 569.180 ;
        RECT -73.090 566.165 -71.710 566.525 ;
        RECT -48.700 566.165 -47.570 568.850 ;
        RECT -42.665 568.795 -42.465 568.850 ;
        RECT -73.090 565.035 -47.570 566.165 ;
        RECT -33.725 566.115 -32.360 567.590 ;
        RECT -73.090 564.590 -71.710 565.035 ;
        RECT -61.770 557.030 -61.555 557.720 ;
        RECT -33.265 557.400 -32.570 566.115 ;
        RECT -61.920 556.520 -61.365 557.030 ;
        RECT -61.770 552.595 -61.555 556.520 ;
        RECT -33.390 556.050 -31.965 557.400 ;
        RECT -61.040 553.915 -60.680 554.035 ;
        RECT -61.040 553.565 -53.645 553.915 ;
        RECT -61.040 553.510 -60.680 553.565 ;
        RECT -61.770 552.555 -60.335 552.595 ;
        RECT -61.770 552.385 -57.365 552.555 ;
        RECT -61.770 552.380 -60.335 552.385 ;
        RECT -61.770 552.170 -61.555 552.380 ;
        RECT -53.995 552.225 -53.645 553.565 ;
        RECT -61.970 552.140 -61.555 552.170 ;
        RECT -63.465 551.970 -61.555 552.140 ;
        RECT -61.970 551.950 -61.555 551.970 ;
        RECT -61.755 551.710 -61.555 551.950 ;
        RECT -61.105 551.520 -60.830 552.210 ;
        RECT -54.855 552.055 -53.645 552.225 ;
        RECT -53.700 551.565 -53.160 551.735 ;
        RECT -61.655 551.305 -60.575 551.520 ;
        RECT -57.415 551.495 -57.025 551.525 ;
        RECT -60.405 551.325 -57.025 551.495 ;
        RECT -57.415 551.315 -57.025 551.325 ;
        RECT -61.655 549.975 -61.455 551.305 ;
        RECT -60.770 551.025 -60.575 551.305 ;
        RECT -60.770 551.005 -60.305 551.025 ;
        RECT -61.215 550.095 -60.940 550.870 ;
        RECT -60.770 550.835 -57.365 551.005 ;
        RECT -60.770 550.815 -60.305 550.835 ;
        RECT -60.760 550.515 -60.315 550.540 ;
        RECT -57.195 550.535 -57.025 551.315 ;
        RECT -54.855 551.075 -54.315 551.245 ;
        RECT -53.700 550.585 -53.160 550.755 ;
        RECT -57.405 550.515 -57.025 550.535 ;
        RECT -60.760 550.345 -57.025 550.515 ;
        RECT -60.760 550.330 -60.315 550.345 ;
        RECT -62.005 549.950 -61.455 549.975 ;
        RECT -63.465 549.780 -61.455 549.950 ;
        RECT -62.005 549.750 -61.455 549.780 ;
        RECT -61.755 548.745 -61.480 549.520 ;
        RECT -61.695 548.560 -61.525 548.745 ;
        RECT -61.170 548.420 -60.990 550.095 ;
        RECT -60.760 549.480 -60.580 550.330 ;
        RECT -57.405 550.325 -57.025 550.345 ;
        RECT -54.855 550.095 -54.315 550.265 ;
        RECT -54.145 549.505 -53.845 549.870 ;
        RECT -60.760 549.460 -60.285 549.480 ;
        RECT -60.760 549.290 -57.365 549.460 ;
        RECT -60.760 549.270 -60.285 549.290 ;
        RECT -54.080 549.200 -53.875 549.505 ;
        RECT -54.080 549.145 -52.980 549.200 ;
        RECT -54.080 549.005 -52.940 549.145 ;
        RECT -53.940 548.895 -52.940 549.005 ;
        RECT -59.015 548.420 -58.665 548.450 ;
        RECT -61.180 548.070 -58.665 548.420 ;
        RECT -53.130 548.200 -52.940 548.895 ;
        RECT -52.705 548.460 -52.350 548.830 ;
        RECT -52.165 548.520 -50.625 548.690 ;
        RECT -59.015 547.230 -58.665 548.070 ;
        RECT -54.850 548.030 -52.940 548.200 ;
        RECT -59.015 547.060 -57.805 547.230 ;
        RECT -53.130 547.220 -52.940 548.030 ;
        RECT -54.850 547.050 -52.940 547.220 ;
        RECT -59.500 546.570 -58.960 546.740 ;
        RECT -58.345 546.080 -57.805 546.250 ;
        RECT -53.095 546.135 -52.825 546.810 ;
        RECT -52.575 546.755 -52.380 548.460 ;
        RECT -48.655 548.455 -43.800 548.645 ;
        RECT -52.165 548.030 -50.625 548.200 ;
        RECT -52.165 547.540 -50.625 547.710 ;
        RECT -52.575 546.405 -52.375 546.755 ;
        RECT -52.165 546.560 -50.625 546.730 ;
        RECT -52.585 546.400 -52.375 546.405 ;
        RECT -53.065 546.035 -52.865 546.135 ;
        RECT -59.500 545.590 -58.960 545.760 ;
        RECT -58.345 545.100 -57.805 545.270 ;
        RECT -53.055 545.000 -52.875 546.035 ;
        RECT -58.815 544.510 -58.515 544.875 ;
        RECT -58.785 544.205 -58.580 544.510 ;
        RECT -59.680 544.150 -58.580 544.205 ;
        RECT -59.720 544.010 -58.580 544.150 ;
        RECT -54.205 544.145 -53.165 544.315 ;
        RECT -59.720 543.900 -58.720 544.010 ;
        RECT -62.035 543.525 -60.495 543.695 ;
        RECT -60.310 543.465 -59.955 543.835 ;
        RECT -62.035 543.035 -60.495 543.205 ;
        RECT -62.035 542.545 -60.495 542.715 ;
        RECT -60.280 541.760 -60.085 543.465 ;
        RECT -59.720 543.205 -59.530 543.900 ;
        RECT -52.585 543.825 -52.385 546.400 ;
        RECT -52.585 543.660 -51.515 543.825 ;
        RECT -52.555 543.655 -51.515 543.660 ;
        RECT -59.720 543.035 -57.810 543.205 ;
        RECT -54.205 543.165 -53.165 543.335 ;
        RECT -59.720 542.225 -59.530 543.035 ;
        RECT -52.555 542.675 -51.515 542.845 ;
        RECT -59.720 542.055 -57.810 542.225 ;
        RECT -54.205 542.185 -53.165 542.355 ;
        RECT -62.035 541.565 -60.495 541.735 ;
        RECT -60.285 541.410 -60.085 541.760 ;
        RECT -52.995 541.595 -52.695 541.960 ;
        RECT -60.285 541.405 -60.075 541.410 ;
        RECT -60.275 540.275 -60.075 541.405 ;
        RECT -52.930 541.375 -52.725 541.595 ;
        RECT -53.015 541.240 -52.265 541.375 ;
        RECT -53.265 540.860 -52.265 541.240 ;
        RECT -53.015 540.725 -52.265 540.860 ;
        RECT -52.775 538.580 -52.395 540.725 ;
        RECT -50.815 539.900 -50.545 539.960 ;
        RECT -48.655 539.900 -48.465 548.455 ;
        RECT -43.990 547.375 -43.800 548.455 ;
        RECT -44.240 547.355 -41.150 547.375 ;
        RECT -45.755 547.185 -41.150 547.355 ;
        RECT -43.250 546.610 -42.955 546.880 ;
        RECT -43.210 546.350 -43.040 546.610 ;
        RECT -42.465 546.350 -42.195 547.010 ;
        RECT -41.335 546.875 -41.150 547.185 ;
        RECT -41.335 546.865 -40.685 546.875 ;
        RECT -41.335 546.695 -39.235 546.865 ;
        RECT -41.335 546.690 -40.685 546.695 ;
        RECT -43.235 546.215 -41.805 546.350 ;
        RECT -45.755 546.180 -41.805 546.215 ;
        RECT -45.755 546.045 -43.065 546.180 ;
        RECT -43.235 546.040 -43.065 546.045 ;
        RECT -45.755 545.555 -43.215 545.725 ;
        RECT -42.880 545.720 -42.190 545.990 ;
        RECT -41.975 545.725 -41.805 546.180 ;
        RECT -41.975 545.555 -39.235 545.725 ;
        RECT -42.370 544.670 -42.100 545.360 ;
        RECT -45.755 543.925 -43.060 544.095 ;
        RECT -43.235 543.470 -43.060 543.925 ;
        RECT -42.805 543.795 -42.535 544.485 ;
        RECT -42.325 544.095 -42.155 544.670 ;
        RECT -42.325 543.925 -39.235 544.095 ;
        RECT -45.755 543.300 -43.060 543.470 ;
        RECT -42.325 543.465 -42.155 543.925 ;
        RECT -42.890 543.295 -42.155 543.465 ;
        RECT -39.250 543.445 -38.885 543.450 ;
        RECT -42.890 542.980 -42.720 543.295 ;
        RECT -41.775 543.275 -38.885 543.445 ;
        RECT -45.755 542.810 -42.720 542.980 ;
        RECT -42.530 542.955 -41.740 542.960 ;
        RECT -42.530 542.785 -39.235 542.955 ;
        RECT -42.530 542.770 -41.740 542.785 ;
        RECT -43.570 542.285 -42.880 542.315 ;
        RECT -42.530 542.285 -42.340 542.770 ;
        RECT -39.055 542.465 -38.885 543.275 ;
        RECT -41.775 542.295 -38.885 542.465 ;
        RECT -39.255 542.290 -38.885 542.295 ;
        RECT -43.570 542.095 -42.340 542.285 ;
        RECT -43.570 542.045 -42.880 542.095 ;
        RECT -42.530 541.120 -42.340 542.095 ;
        RECT -39.055 542.045 -38.885 542.290 ;
        RECT -45.755 540.950 -42.340 541.120 ;
        RECT -42.165 541.845 -38.885 542.045 ;
        RECT -42.165 541.120 -41.965 541.845 ;
        RECT -42.165 540.950 -39.235 541.120 ;
        RECT -42.165 540.945 -41.735 540.950 ;
        RECT -43.485 540.045 -43.215 540.735 ;
        RECT -50.815 539.710 -48.465 539.900 ;
        RECT -50.815 539.595 -50.545 539.710 ;
        RECT -44.460 539.355 -44.065 539.415 ;
        RECT -43.430 539.355 -43.260 540.045 ;
        RECT -42.805 539.765 -42.535 540.455 ;
        RECT -44.460 539.020 -43.260 539.355 ;
        RECT -44.110 538.995 -43.260 539.020 ;
        RECT -52.775 538.200 -48.495 538.580 ;
        RECT -61.615 537.775 -60.155 537.990 ;
        RECT -61.615 534.255 -61.400 537.775 ;
        RECT -60.370 536.780 -60.155 537.775 ;
        RECT -50.280 536.780 -49.855 536.910 ;
        RECT -60.370 536.565 -49.855 536.780 ;
        RECT -50.280 536.450 -49.855 536.565 ;
        RECT -60.885 535.575 -60.525 535.695 ;
        RECT -60.885 535.225 -53.490 535.575 ;
        RECT -60.885 535.170 -60.525 535.225 ;
        RECT -61.615 534.215 -60.180 534.255 ;
        RECT -61.615 534.045 -57.210 534.215 ;
        RECT -61.615 534.040 -60.180 534.045 ;
        RECT -61.615 533.830 -61.400 534.040 ;
        RECT -53.840 533.885 -53.490 535.225 ;
        RECT -61.815 533.800 -61.400 533.830 ;
        RECT -63.310 533.630 -61.400 533.800 ;
        RECT -61.815 533.610 -61.400 533.630 ;
        RECT -61.600 533.370 -61.400 533.610 ;
        RECT -60.950 533.180 -60.675 533.870 ;
        RECT -54.700 533.715 -53.490 533.885 ;
        RECT -53.545 533.225 -53.005 533.395 ;
        RECT -61.500 532.965 -60.420 533.180 ;
        RECT -57.260 533.155 -56.870 533.185 ;
        RECT -60.250 532.985 -56.870 533.155 ;
        RECT -57.260 532.975 -56.870 532.985 ;
        RECT -61.500 531.635 -61.300 532.965 ;
        RECT -60.615 532.685 -60.420 532.965 ;
        RECT -60.615 532.665 -60.150 532.685 ;
        RECT -61.060 531.755 -60.785 532.530 ;
        RECT -60.615 532.495 -57.210 532.665 ;
        RECT -60.615 532.475 -60.150 532.495 ;
        RECT -60.605 532.175 -60.160 532.200 ;
        RECT -57.040 532.195 -56.870 532.975 ;
        RECT -54.700 532.735 -54.160 532.905 ;
        RECT -53.545 532.245 -53.005 532.415 ;
        RECT -57.250 532.175 -56.870 532.195 ;
        RECT -60.605 532.005 -56.870 532.175 ;
        RECT -60.605 531.990 -60.160 532.005 ;
        RECT -61.850 531.610 -61.300 531.635 ;
        RECT -63.310 531.440 -61.300 531.610 ;
        RECT -61.850 531.410 -61.300 531.440 ;
        RECT -61.600 530.405 -61.325 531.180 ;
        RECT -61.540 530.220 -61.370 530.405 ;
        RECT -61.015 530.080 -60.835 531.755 ;
        RECT -60.605 531.140 -60.425 531.990 ;
        RECT -57.250 531.985 -56.870 532.005 ;
        RECT -54.700 531.755 -54.160 531.925 ;
        RECT -53.990 531.165 -53.690 531.530 ;
        RECT -60.605 531.120 -60.130 531.140 ;
        RECT -60.605 530.950 -57.210 531.120 ;
        RECT -60.605 530.930 -60.130 530.950 ;
        RECT -53.925 530.860 -53.720 531.165 ;
        RECT -53.925 530.805 -52.825 530.860 ;
        RECT -53.925 530.665 -52.785 530.805 ;
        RECT -53.785 530.555 -52.785 530.665 ;
        RECT -58.860 530.080 -58.510 530.110 ;
        RECT -61.025 529.730 -58.510 530.080 ;
        RECT -52.975 529.860 -52.785 530.555 ;
        RECT -52.550 530.120 -52.195 530.490 ;
        RECT -52.010 530.180 -50.470 530.350 ;
        RECT -58.860 528.890 -58.510 529.730 ;
        RECT -54.695 529.690 -52.785 529.860 ;
        RECT -58.860 528.720 -57.650 528.890 ;
        RECT -52.975 528.880 -52.785 529.690 ;
        RECT -54.695 528.710 -52.785 528.880 ;
        RECT -59.345 528.230 -58.805 528.400 ;
        RECT -58.190 527.740 -57.650 527.910 ;
        RECT -52.940 527.795 -52.670 528.470 ;
        RECT -52.420 528.415 -52.225 530.120 ;
        RECT -52.010 529.690 -50.470 529.860 ;
        RECT -52.010 529.200 -50.470 529.370 ;
        RECT -52.420 528.065 -52.220 528.415 ;
        RECT -52.010 528.220 -50.470 528.390 ;
        RECT -52.430 528.060 -52.220 528.065 ;
        RECT -52.910 527.695 -52.710 527.795 ;
        RECT -59.345 527.250 -58.805 527.420 ;
        RECT -58.190 526.760 -57.650 526.930 ;
        RECT -52.900 526.660 -52.720 527.695 ;
        RECT -58.660 526.170 -58.360 526.535 ;
        RECT -58.630 525.865 -58.425 526.170 ;
        RECT -59.525 525.810 -58.425 525.865 ;
        RECT -59.565 525.670 -58.425 525.810 ;
        RECT -54.050 525.805 -53.010 525.975 ;
        RECT -59.565 525.560 -58.565 525.670 ;
        RECT -61.880 525.185 -60.340 525.355 ;
        RECT -60.155 525.125 -59.800 525.495 ;
        RECT -61.880 524.695 -60.340 524.865 ;
        RECT -61.880 524.205 -60.340 524.375 ;
        RECT -60.125 523.420 -59.930 525.125 ;
        RECT -59.565 524.865 -59.375 525.560 ;
        RECT -52.430 525.485 -52.230 528.060 ;
        RECT -52.430 525.320 -51.360 525.485 ;
        RECT -52.400 525.315 -51.360 525.320 ;
        RECT -59.565 524.695 -57.655 524.865 ;
        RECT -54.050 524.825 -53.010 524.995 ;
        RECT -59.565 523.885 -59.375 524.695 ;
        RECT -52.400 524.335 -51.360 524.505 ;
        RECT -59.565 523.715 -57.655 523.885 ;
        RECT -54.050 523.845 -53.010 524.015 ;
        RECT -61.880 523.225 -60.340 523.395 ;
        RECT -60.130 523.070 -59.930 523.420 ;
        RECT -52.840 523.255 -52.540 523.620 ;
        RECT -60.130 523.065 -59.920 523.070 ;
        RECT -60.120 521.935 -59.920 523.065 ;
        RECT -52.775 523.035 -52.570 523.255 ;
        RECT -52.860 522.740 -52.110 523.035 ;
        RECT -52.860 522.410 -49.785 522.740 ;
        RECT -48.875 522.410 -48.495 538.200 ;
        RECT -42.755 538.030 -42.585 539.765 ;
        RECT -44.350 537.815 -42.585 538.030 ;
        RECT -44.350 534.295 -44.135 537.815 ;
        RECT -43.620 535.615 -43.260 535.735 ;
        RECT -43.620 535.265 -36.225 535.615 ;
        RECT -43.620 535.210 -43.260 535.265 ;
        RECT -44.350 534.255 -42.915 534.295 ;
        RECT -44.350 534.085 -39.945 534.255 ;
        RECT -44.350 534.080 -42.915 534.085 ;
        RECT -44.350 533.870 -44.135 534.080 ;
        RECT -36.575 533.925 -36.225 535.265 ;
        RECT -44.550 533.840 -44.135 533.870 ;
        RECT -46.045 533.670 -44.135 533.840 ;
        RECT -44.550 533.650 -44.135 533.670 ;
        RECT -44.335 533.410 -44.135 533.650 ;
        RECT -43.685 533.220 -43.410 533.910 ;
        RECT -37.435 533.755 -36.225 533.925 ;
        RECT -36.280 533.265 -35.740 533.435 ;
        RECT -44.235 533.005 -43.155 533.220 ;
        RECT -39.995 533.195 -39.605 533.225 ;
        RECT -42.985 533.025 -39.605 533.195 ;
        RECT -39.995 533.015 -39.605 533.025 ;
        RECT -44.235 531.675 -44.035 533.005 ;
        RECT -43.350 532.725 -43.155 533.005 ;
        RECT -43.350 532.705 -42.885 532.725 ;
        RECT -43.795 531.795 -43.520 532.570 ;
        RECT -43.350 532.535 -39.945 532.705 ;
        RECT -43.350 532.515 -42.885 532.535 ;
        RECT -43.340 532.215 -42.895 532.240 ;
        RECT -39.775 532.235 -39.605 533.015 ;
        RECT -37.435 532.775 -36.895 532.945 ;
        RECT -36.280 532.285 -35.740 532.455 ;
        RECT -39.985 532.215 -39.605 532.235 ;
        RECT -43.340 532.045 -39.605 532.215 ;
        RECT -43.340 532.030 -42.895 532.045 ;
        RECT -44.585 531.650 -44.035 531.675 ;
        RECT -46.045 531.480 -44.035 531.650 ;
        RECT -44.585 531.450 -44.035 531.480 ;
        RECT -44.335 530.445 -44.060 531.220 ;
        RECT -44.275 530.260 -44.105 530.445 ;
        RECT -43.750 530.120 -43.570 531.795 ;
        RECT -43.340 531.180 -43.160 532.030 ;
        RECT -39.985 532.025 -39.605 532.045 ;
        RECT -37.435 531.795 -36.895 531.965 ;
        RECT -36.725 531.205 -36.425 531.570 ;
        RECT -43.340 531.160 -42.865 531.180 ;
        RECT -43.340 530.990 -39.945 531.160 ;
        RECT -43.340 530.970 -42.865 530.990 ;
        RECT -36.660 530.900 -36.455 531.205 ;
        RECT -36.660 530.845 -35.560 530.900 ;
        RECT -36.660 530.705 -35.520 530.845 ;
        RECT -36.520 530.595 -35.520 530.705 ;
        RECT -41.595 530.120 -41.245 530.150 ;
        RECT -43.760 529.770 -41.245 530.120 ;
        RECT -35.710 529.900 -35.520 530.595 ;
        RECT -35.285 530.160 -34.930 530.530 ;
        RECT -34.745 530.220 -33.205 530.390 ;
        RECT -41.595 528.930 -41.245 529.770 ;
        RECT -37.430 529.730 -35.520 529.900 ;
        RECT -41.595 528.760 -40.385 528.930 ;
        RECT -35.710 528.920 -35.520 529.730 ;
        RECT -37.430 528.750 -35.520 528.920 ;
        RECT -42.080 528.270 -41.540 528.440 ;
        RECT -40.925 527.780 -40.385 527.950 ;
        RECT -35.675 527.835 -35.405 528.510 ;
        RECT -35.155 528.455 -34.960 530.160 ;
        RECT -34.745 529.730 -33.205 529.900 ;
        RECT -34.745 529.240 -33.205 529.410 ;
        RECT -35.155 528.105 -34.955 528.455 ;
        RECT -34.745 528.260 -33.205 528.430 ;
        RECT -35.165 528.100 -34.955 528.105 ;
        RECT -35.645 527.735 -35.445 527.835 ;
        RECT -42.080 527.290 -41.540 527.460 ;
        RECT -40.925 526.800 -40.385 526.970 ;
        RECT -35.635 526.700 -35.455 527.735 ;
        RECT -41.395 526.210 -41.095 526.575 ;
        RECT -41.365 525.905 -41.160 526.210 ;
        RECT -42.260 525.850 -41.160 525.905 ;
        RECT -42.300 525.710 -41.160 525.850 ;
        RECT -36.785 525.845 -35.745 526.015 ;
        RECT -42.300 525.600 -41.300 525.710 ;
        RECT -44.615 525.225 -43.075 525.395 ;
        RECT -42.890 525.165 -42.535 525.535 ;
        RECT -44.615 524.735 -43.075 524.905 ;
        RECT -44.615 524.245 -43.075 524.415 ;
        RECT -42.860 523.460 -42.665 525.165 ;
        RECT -42.300 524.905 -42.110 525.600 ;
        RECT -35.165 525.525 -34.965 528.100 ;
        RECT -35.165 525.360 -34.095 525.525 ;
        RECT -35.135 525.355 -34.095 525.360 ;
        RECT -42.300 524.735 -40.390 524.905 ;
        RECT -36.785 524.865 -35.745 525.035 ;
        RECT -42.300 523.925 -42.110 524.735 ;
        RECT -35.135 524.375 -34.095 524.545 ;
        RECT -42.300 523.755 -40.390 523.925 ;
        RECT -36.785 523.885 -35.745 524.055 ;
        RECT -44.615 523.265 -43.075 523.435 ;
        RECT -42.865 523.110 -42.665 523.460 ;
        RECT -35.575 523.295 -35.275 523.660 ;
        RECT -42.865 523.105 -42.655 523.110 ;
        RECT -42.855 522.410 -42.655 523.105 ;
        RECT -35.510 523.075 -35.305 523.295 ;
        RECT -35.595 522.425 -34.845 523.075 ;
        RECT -52.860 522.385 -42.655 522.410 ;
        RECT -52.655 522.360 -42.655 522.385 ;
        RECT -50.165 522.030 -42.655 522.360 ;
        RECT -68.895 519.505 -67.995 519.690 ;
        RECT -48.815 519.505 -47.965 522.030 ;
        RECT -42.855 521.975 -42.655 522.030 ;
        RECT -33.870 519.840 -32.670 521.180 ;
        RECT -68.895 518.655 -47.965 519.505 ;
        RECT -68.895 518.460 -67.995 518.655 ;
        RECT -61.855 511.395 -61.640 511.955 ;
        RECT -33.530 511.590 -32.875 519.840 ;
        RECT -62.355 510.090 -60.835 511.395 ;
        RECT -61.855 506.830 -61.640 510.090 ;
        RECT -33.850 509.900 -32.395 511.590 ;
        RECT -61.125 508.150 -60.765 508.270 ;
        RECT -61.125 507.800 -53.730 508.150 ;
        RECT -61.125 507.745 -60.765 507.800 ;
        RECT -61.855 506.790 -60.420 506.830 ;
        RECT -61.855 506.620 -57.450 506.790 ;
        RECT -61.855 506.615 -60.420 506.620 ;
        RECT -61.855 506.405 -61.640 506.615 ;
        RECT -54.080 506.460 -53.730 507.800 ;
        RECT -62.055 506.375 -61.640 506.405 ;
        RECT -63.550 506.205 -61.640 506.375 ;
        RECT -62.055 506.185 -61.640 506.205 ;
        RECT -61.840 505.945 -61.640 506.185 ;
        RECT -61.190 505.755 -60.915 506.445 ;
        RECT -54.940 506.290 -53.730 506.460 ;
        RECT -53.785 505.800 -53.245 505.970 ;
        RECT -61.740 505.540 -60.660 505.755 ;
        RECT -57.500 505.730 -57.110 505.760 ;
        RECT -60.490 505.560 -57.110 505.730 ;
        RECT -57.500 505.550 -57.110 505.560 ;
        RECT -61.740 504.210 -61.540 505.540 ;
        RECT -60.855 505.260 -60.660 505.540 ;
        RECT -60.855 505.240 -60.390 505.260 ;
        RECT -61.300 504.330 -61.025 505.105 ;
        RECT -60.855 505.070 -57.450 505.240 ;
        RECT -60.855 505.050 -60.390 505.070 ;
        RECT -60.845 504.750 -60.400 504.775 ;
        RECT -57.280 504.770 -57.110 505.550 ;
        RECT -54.940 505.310 -54.400 505.480 ;
        RECT -53.785 504.820 -53.245 504.990 ;
        RECT -57.490 504.750 -57.110 504.770 ;
        RECT -60.845 504.580 -57.110 504.750 ;
        RECT -60.845 504.565 -60.400 504.580 ;
        RECT -62.090 504.185 -61.540 504.210 ;
        RECT -63.550 504.015 -61.540 504.185 ;
        RECT -62.090 503.985 -61.540 504.015 ;
        RECT -61.840 502.980 -61.565 503.755 ;
        RECT -61.780 502.795 -61.610 502.980 ;
        RECT -61.255 502.655 -61.075 504.330 ;
        RECT -60.845 503.715 -60.665 504.565 ;
        RECT -57.490 504.560 -57.110 504.580 ;
        RECT -54.940 504.330 -54.400 504.500 ;
        RECT -54.230 503.740 -53.930 504.105 ;
        RECT -60.845 503.695 -60.370 503.715 ;
        RECT -60.845 503.525 -57.450 503.695 ;
        RECT -60.845 503.505 -60.370 503.525 ;
        RECT -54.165 503.435 -53.960 503.740 ;
        RECT -54.165 503.380 -53.065 503.435 ;
        RECT -54.165 503.240 -53.025 503.380 ;
        RECT -54.025 503.130 -53.025 503.240 ;
        RECT -59.100 502.655 -58.750 502.685 ;
        RECT -61.265 502.305 -58.750 502.655 ;
        RECT -53.215 502.435 -53.025 503.130 ;
        RECT -52.790 502.695 -52.435 503.065 ;
        RECT -52.250 502.755 -50.710 502.925 ;
        RECT -59.100 501.465 -58.750 502.305 ;
        RECT -54.935 502.265 -53.025 502.435 ;
        RECT -59.100 501.295 -57.890 501.465 ;
        RECT -53.215 501.455 -53.025 502.265 ;
        RECT -54.935 501.285 -53.025 501.455 ;
        RECT -59.585 500.805 -59.045 500.975 ;
        RECT -58.430 500.315 -57.890 500.485 ;
        RECT -53.180 500.370 -52.910 501.045 ;
        RECT -52.660 500.990 -52.465 502.695 ;
        RECT -48.740 502.690 -43.885 502.880 ;
        RECT -52.250 502.265 -50.710 502.435 ;
        RECT -52.250 501.775 -50.710 501.945 ;
        RECT -52.660 500.640 -52.460 500.990 ;
        RECT -52.250 500.795 -50.710 500.965 ;
        RECT -52.670 500.635 -52.460 500.640 ;
        RECT -53.150 500.270 -52.950 500.370 ;
        RECT -59.585 499.825 -59.045 499.995 ;
        RECT -58.430 499.335 -57.890 499.505 ;
        RECT -53.140 499.235 -52.960 500.270 ;
        RECT -58.900 498.745 -58.600 499.110 ;
        RECT -58.870 498.440 -58.665 498.745 ;
        RECT -59.765 498.385 -58.665 498.440 ;
        RECT -59.805 498.245 -58.665 498.385 ;
        RECT -54.290 498.380 -53.250 498.550 ;
        RECT -59.805 498.135 -58.805 498.245 ;
        RECT -62.120 497.760 -60.580 497.930 ;
        RECT -60.395 497.700 -60.040 498.070 ;
        RECT -62.120 497.270 -60.580 497.440 ;
        RECT -62.120 496.780 -60.580 496.950 ;
        RECT -60.365 495.995 -60.170 497.700 ;
        RECT -59.805 497.440 -59.615 498.135 ;
        RECT -52.670 498.060 -52.470 500.635 ;
        RECT -52.670 497.895 -51.600 498.060 ;
        RECT -52.640 497.890 -51.600 497.895 ;
        RECT -59.805 497.270 -57.895 497.440 ;
        RECT -54.290 497.400 -53.250 497.570 ;
        RECT -59.805 496.460 -59.615 497.270 ;
        RECT -52.640 496.910 -51.600 497.080 ;
        RECT -59.805 496.290 -57.895 496.460 ;
        RECT -54.290 496.420 -53.250 496.590 ;
        RECT -62.120 495.800 -60.580 495.970 ;
        RECT -60.370 495.645 -60.170 495.995 ;
        RECT -53.080 495.830 -52.780 496.195 ;
        RECT -60.370 495.640 -60.160 495.645 ;
        RECT -60.360 494.510 -60.160 495.640 ;
        RECT -53.015 495.610 -52.810 495.830 ;
        RECT -53.100 495.475 -52.350 495.610 ;
        RECT -53.350 495.095 -52.350 495.475 ;
        RECT -53.100 494.960 -52.350 495.095 ;
        RECT -52.860 492.815 -52.480 494.960 ;
        RECT -50.900 494.135 -50.630 494.195 ;
        RECT -48.740 494.135 -48.550 502.690 ;
        RECT -44.075 501.610 -43.885 502.690 ;
        RECT -44.325 501.590 -41.235 501.610 ;
        RECT -45.840 501.420 -41.235 501.590 ;
        RECT -43.335 500.845 -43.040 501.115 ;
        RECT -43.295 500.585 -43.125 500.845 ;
        RECT -42.550 500.585 -42.280 501.245 ;
        RECT -41.420 501.110 -41.235 501.420 ;
        RECT -41.420 501.100 -40.770 501.110 ;
        RECT -41.420 500.930 -39.320 501.100 ;
        RECT -41.420 500.925 -40.770 500.930 ;
        RECT -43.320 500.450 -41.890 500.585 ;
        RECT -45.840 500.415 -41.890 500.450 ;
        RECT -45.840 500.280 -43.150 500.415 ;
        RECT -43.320 500.275 -43.150 500.280 ;
        RECT -45.840 499.790 -43.300 499.960 ;
        RECT -42.965 499.955 -42.275 500.225 ;
        RECT -42.060 499.960 -41.890 500.415 ;
        RECT -42.060 499.790 -39.320 499.960 ;
        RECT -42.455 498.905 -42.185 499.595 ;
        RECT -45.840 498.160 -43.145 498.330 ;
        RECT -43.320 497.705 -43.145 498.160 ;
        RECT -42.890 498.030 -42.620 498.720 ;
        RECT -42.410 498.330 -42.240 498.905 ;
        RECT -42.410 498.160 -39.320 498.330 ;
        RECT -45.840 497.535 -43.145 497.705 ;
        RECT -42.410 497.700 -42.240 498.160 ;
        RECT -42.975 497.530 -42.240 497.700 ;
        RECT -39.335 497.680 -38.970 497.685 ;
        RECT -42.975 497.215 -42.805 497.530 ;
        RECT -41.860 497.510 -38.970 497.680 ;
        RECT -45.840 497.045 -42.805 497.215 ;
        RECT -42.615 497.190 -41.825 497.195 ;
        RECT -42.615 497.020 -39.320 497.190 ;
        RECT -42.615 497.005 -41.825 497.020 ;
        RECT -43.655 496.520 -42.965 496.550 ;
        RECT -42.615 496.520 -42.425 497.005 ;
        RECT -39.140 496.700 -38.970 497.510 ;
        RECT -41.860 496.530 -38.970 496.700 ;
        RECT -39.340 496.525 -38.970 496.530 ;
        RECT -43.655 496.330 -42.425 496.520 ;
        RECT -43.655 496.280 -42.965 496.330 ;
        RECT -42.615 495.355 -42.425 496.330 ;
        RECT -39.140 496.280 -38.970 496.525 ;
        RECT -45.840 495.185 -42.425 495.355 ;
        RECT -42.250 496.080 -38.970 496.280 ;
        RECT -42.250 495.355 -42.050 496.080 ;
        RECT -42.250 495.185 -39.320 495.355 ;
        RECT -42.250 495.180 -41.820 495.185 ;
        RECT -43.570 494.280 -43.300 494.970 ;
        RECT -50.900 493.945 -48.550 494.135 ;
        RECT -50.900 493.830 -50.630 493.945 ;
        RECT -44.545 493.590 -44.150 493.650 ;
        RECT -43.515 493.590 -43.345 494.280 ;
        RECT -42.890 494.000 -42.620 494.690 ;
        RECT -44.545 493.255 -43.345 493.590 ;
        RECT -44.195 493.230 -43.345 493.255 ;
        RECT -52.860 492.435 -48.580 492.815 ;
        RECT -61.700 492.010 -60.240 492.225 ;
        RECT -61.700 488.490 -61.485 492.010 ;
        RECT -60.455 491.015 -60.240 492.010 ;
        RECT -50.365 491.015 -49.940 491.145 ;
        RECT -60.455 490.800 -49.940 491.015 ;
        RECT -50.365 490.685 -49.940 490.800 ;
        RECT -60.970 489.810 -60.610 489.930 ;
        RECT -60.970 489.460 -53.575 489.810 ;
        RECT -60.970 489.405 -60.610 489.460 ;
        RECT -61.700 488.450 -60.265 488.490 ;
        RECT -61.700 488.280 -57.295 488.450 ;
        RECT -61.700 488.275 -60.265 488.280 ;
        RECT -61.700 488.065 -61.485 488.275 ;
        RECT -53.925 488.120 -53.575 489.460 ;
        RECT -61.900 488.035 -61.485 488.065 ;
        RECT -63.395 487.865 -61.485 488.035 ;
        RECT -61.900 487.845 -61.485 487.865 ;
        RECT -61.685 487.605 -61.485 487.845 ;
        RECT -61.035 487.415 -60.760 488.105 ;
        RECT -54.785 487.950 -53.575 488.120 ;
        RECT -53.630 487.460 -53.090 487.630 ;
        RECT -61.585 487.200 -60.505 487.415 ;
        RECT -57.345 487.390 -56.955 487.420 ;
        RECT -60.335 487.220 -56.955 487.390 ;
        RECT -57.345 487.210 -56.955 487.220 ;
        RECT -61.585 485.870 -61.385 487.200 ;
        RECT -60.700 486.920 -60.505 487.200 ;
        RECT -60.700 486.900 -60.235 486.920 ;
        RECT -61.145 485.990 -60.870 486.765 ;
        RECT -60.700 486.730 -57.295 486.900 ;
        RECT -60.700 486.710 -60.235 486.730 ;
        RECT -60.690 486.410 -60.245 486.435 ;
        RECT -57.125 486.430 -56.955 487.210 ;
        RECT -54.785 486.970 -54.245 487.140 ;
        RECT -53.630 486.480 -53.090 486.650 ;
        RECT -57.335 486.410 -56.955 486.430 ;
        RECT -60.690 486.240 -56.955 486.410 ;
        RECT -60.690 486.225 -60.245 486.240 ;
        RECT -61.935 485.845 -61.385 485.870 ;
        RECT -63.395 485.675 -61.385 485.845 ;
        RECT -61.935 485.645 -61.385 485.675 ;
        RECT -61.685 484.640 -61.410 485.415 ;
        RECT -61.625 484.455 -61.455 484.640 ;
        RECT -61.100 484.315 -60.920 485.990 ;
        RECT -60.690 485.375 -60.510 486.225 ;
        RECT -57.335 486.220 -56.955 486.240 ;
        RECT -54.785 485.990 -54.245 486.160 ;
        RECT -54.075 485.400 -53.775 485.765 ;
        RECT -60.690 485.355 -60.215 485.375 ;
        RECT -60.690 485.185 -57.295 485.355 ;
        RECT -60.690 485.165 -60.215 485.185 ;
        RECT -54.010 485.095 -53.805 485.400 ;
        RECT -54.010 485.040 -52.910 485.095 ;
        RECT -54.010 484.900 -52.870 485.040 ;
        RECT -53.870 484.790 -52.870 484.900 ;
        RECT -58.945 484.315 -58.595 484.345 ;
        RECT -61.110 483.965 -58.595 484.315 ;
        RECT -53.060 484.095 -52.870 484.790 ;
        RECT -52.635 484.355 -52.280 484.725 ;
        RECT -52.095 484.415 -50.555 484.585 ;
        RECT -58.945 483.125 -58.595 483.965 ;
        RECT -54.780 483.925 -52.870 484.095 ;
        RECT -58.945 482.955 -57.735 483.125 ;
        RECT -53.060 483.115 -52.870 483.925 ;
        RECT -54.780 482.945 -52.870 483.115 ;
        RECT -59.430 482.465 -58.890 482.635 ;
        RECT -58.275 481.975 -57.735 482.145 ;
        RECT -53.025 482.030 -52.755 482.705 ;
        RECT -52.505 482.650 -52.310 484.355 ;
        RECT -52.095 483.925 -50.555 484.095 ;
        RECT -52.095 483.435 -50.555 483.605 ;
        RECT -52.505 482.300 -52.305 482.650 ;
        RECT -52.095 482.455 -50.555 482.625 ;
        RECT -52.515 482.295 -52.305 482.300 ;
        RECT -52.995 481.930 -52.795 482.030 ;
        RECT -59.430 481.485 -58.890 481.655 ;
        RECT -58.275 480.995 -57.735 481.165 ;
        RECT -52.985 480.895 -52.805 481.930 ;
        RECT -58.745 480.405 -58.445 480.770 ;
        RECT -58.715 480.100 -58.510 480.405 ;
        RECT -59.610 480.045 -58.510 480.100 ;
        RECT -59.650 479.905 -58.510 480.045 ;
        RECT -54.135 480.040 -53.095 480.210 ;
        RECT -59.650 479.795 -58.650 479.905 ;
        RECT -61.965 479.420 -60.425 479.590 ;
        RECT -60.240 479.360 -59.885 479.730 ;
        RECT -61.965 478.930 -60.425 479.100 ;
        RECT -61.965 478.440 -60.425 478.610 ;
        RECT -60.210 477.655 -60.015 479.360 ;
        RECT -59.650 479.100 -59.460 479.795 ;
        RECT -52.515 479.720 -52.315 482.295 ;
        RECT -52.515 479.555 -51.445 479.720 ;
        RECT -52.485 479.550 -51.445 479.555 ;
        RECT -59.650 478.930 -57.740 479.100 ;
        RECT -54.135 479.060 -53.095 479.230 ;
        RECT -59.650 478.120 -59.460 478.930 ;
        RECT -52.485 478.570 -51.445 478.740 ;
        RECT -59.650 477.950 -57.740 478.120 ;
        RECT -54.135 478.080 -53.095 478.250 ;
        RECT -61.965 477.460 -60.425 477.630 ;
        RECT -60.215 477.305 -60.015 477.655 ;
        RECT -52.925 477.490 -52.625 477.855 ;
        RECT -60.215 477.300 -60.005 477.305 ;
        RECT -60.205 476.170 -60.005 477.300 ;
        RECT -52.860 477.270 -52.655 477.490 ;
        RECT -52.945 476.975 -52.195 477.270 ;
        RECT -52.945 476.645 -49.870 476.975 ;
        RECT -48.960 476.645 -48.580 492.435 ;
        RECT -42.840 492.265 -42.670 494.000 ;
        RECT -44.435 492.050 -42.670 492.265 ;
        RECT -44.435 488.530 -44.220 492.050 ;
        RECT -43.705 489.850 -43.345 489.970 ;
        RECT -43.705 489.500 -36.310 489.850 ;
        RECT -43.705 489.445 -43.345 489.500 ;
        RECT -44.435 488.490 -43.000 488.530 ;
        RECT -44.435 488.320 -40.030 488.490 ;
        RECT -44.435 488.315 -43.000 488.320 ;
        RECT -44.435 488.105 -44.220 488.315 ;
        RECT -36.660 488.160 -36.310 489.500 ;
        RECT -44.635 488.075 -44.220 488.105 ;
        RECT -46.130 487.905 -44.220 488.075 ;
        RECT -44.635 487.885 -44.220 487.905 ;
        RECT -44.420 487.645 -44.220 487.885 ;
        RECT -43.770 487.455 -43.495 488.145 ;
        RECT -37.520 487.990 -36.310 488.160 ;
        RECT -36.365 487.500 -35.825 487.670 ;
        RECT -44.320 487.240 -43.240 487.455 ;
        RECT -40.080 487.430 -39.690 487.460 ;
        RECT -43.070 487.260 -39.690 487.430 ;
        RECT -40.080 487.250 -39.690 487.260 ;
        RECT -44.320 485.910 -44.120 487.240 ;
        RECT -43.435 486.960 -43.240 487.240 ;
        RECT -43.435 486.940 -42.970 486.960 ;
        RECT -43.880 486.030 -43.605 486.805 ;
        RECT -43.435 486.770 -40.030 486.940 ;
        RECT -43.435 486.750 -42.970 486.770 ;
        RECT -43.425 486.450 -42.980 486.475 ;
        RECT -39.860 486.470 -39.690 487.250 ;
        RECT -37.520 487.010 -36.980 487.180 ;
        RECT -36.365 486.520 -35.825 486.690 ;
        RECT -40.070 486.450 -39.690 486.470 ;
        RECT -43.425 486.280 -39.690 486.450 ;
        RECT -43.425 486.265 -42.980 486.280 ;
        RECT -44.670 485.885 -44.120 485.910 ;
        RECT -46.130 485.715 -44.120 485.885 ;
        RECT -44.670 485.685 -44.120 485.715 ;
        RECT -44.420 484.680 -44.145 485.455 ;
        RECT -44.360 484.495 -44.190 484.680 ;
        RECT -43.835 484.355 -43.655 486.030 ;
        RECT -43.425 485.415 -43.245 486.265 ;
        RECT -40.070 486.260 -39.690 486.280 ;
        RECT -37.520 486.030 -36.980 486.200 ;
        RECT -36.810 485.440 -36.510 485.805 ;
        RECT -43.425 485.395 -42.950 485.415 ;
        RECT -43.425 485.225 -40.030 485.395 ;
        RECT -43.425 485.205 -42.950 485.225 ;
        RECT -36.745 485.135 -36.540 485.440 ;
        RECT -36.745 485.080 -35.645 485.135 ;
        RECT -36.745 484.940 -35.605 485.080 ;
        RECT -36.605 484.830 -35.605 484.940 ;
        RECT -41.680 484.355 -41.330 484.385 ;
        RECT -43.845 484.005 -41.330 484.355 ;
        RECT -35.795 484.135 -35.605 484.830 ;
        RECT -35.370 484.395 -35.015 484.765 ;
        RECT -34.830 484.455 -33.290 484.625 ;
        RECT -41.680 483.165 -41.330 484.005 ;
        RECT -37.515 483.965 -35.605 484.135 ;
        RECT -41.680 482.995 -40.470 483.165 ;
        RECT -35.795 483.155 -35.605 483.965 ;
        RECT -37.515 482.985 -35.605 483.155 ;
        RECT -42.165 482.505 -41.625 482.675 ;
        RECT -41.010 482.015 -40.470 482.185 ;
        RECT -35.760 482.070 -35.490 482.745 ;
        RECT -35.240 482.690 -35.045 484.395 ;
        RECT -34.830 483.965 -33.290 484.135 ;
        RECT -34.830 483.475 -33.290 483.645 ;
        RECT -35.240 482.340 -35.040 482.690 ;
        RECT -34.830 482.495 -33.290 482.665 ;
        RECT -35.250 482.335 -35.040 482.340 ;
        RECT -35.730 481.970 -35.530 482.070 ;
        RECT -42.165 481.525 -41.625 481.695 ;
        RECT -41.010 481.035 -40.470 481.205 ;
        RECT -35.720 480.935 -35.540 481.970 ;
        RECT -41.480 480.445 -41.180 480.810 ;
        RECT -41.450 480.140 -41.245 480.445 ;
        RECT -42.345 480.085 -41.245 480.140 ;
        RECT -42.385 479.945 -41.245 480.085 ;
        RECT -36.870 480.080 -35.830 480.250 ;
        RECT -42.385 479.835 -41.385 479.945 ;
        RECT -44.700 479.460 -43.160 479.630 ;
        RECT -42.975 479.400 -42.620 479.770 ;
        RECT -44.700 478.970 -43.160 479.140 ;
        RECT -44.700 478.480 -43.160 478.650 ;
        RECT -42.945 477.695 -42.750 479.400 ;
        RECT -42.385 479.140 -42.195 479.835 ;
        RECT -35.250 479.760 -35.050 482.335 ;
        RECT -35.250 479.595 -34.180 479.760 ;
        RECT -35.220 479.590 -34.180 479.595 ;
        RECT -42.385 478.970 -40.475 479.140 ;
        RECT -36.870 479.100 -35.830 479.270 ;
        RECT -42.385 478.160 -42.195 478.970 ;
        RECT -35.220 478.610 -34.180 478.780 ;
        RECT -42.385 477.990 -40.475 478.160 ;
        RECT -36.870 478.120 -35.830 478.290 ;
        RECT -44.700 477.500 -43.160 477.670 ;
        RECT -42.950 477.345 -42.750 477.695 ;
        RECT -35.660 477.530 -35.360 477.895 ;
        RECT -42.950 477.340 -42.740 477.345 ;
        RECT -42.940 476.645 -42.740 477.340 ;
        RECT -35.595 477.310 -35.390 477.530 ;
        RECT -35.680 476.660 -34.930 477.310 ;
        RECT -52.945 476.620 -42.740 476.645 ;
        RECT -52.740 476.595 -42.740 476.620 ;
        RECT -50.250 476.265 -42.740 476.595 ;
        RECT -73.110 473.785 -71.695 474.135 ;
        RECT -48.845 473.785 -47.760 476.265 ;
        RECT -42.940 476.210 -42.740 476.265 ;
        RECT -33.855 474.025 -32.710 475.275 ;
        RECT -73.110 472.700 -47.760 473.785 ;
        RECT -73.110 472.415 -71.695 472.700 ;
        RECT -62.185 467.725 -61.970 468.185 ;
        RECT -33.600 467.900 -32.845 474.025 ;
        RECT -62.620 466.265 -61.125 467.725 ;
        RECT -62.185 463.060 -61.970 466.265 ;
        RECT -33.940 466.020 -32.370 467.900 ;
        RECT -61.455 464.380 -61.095 464.500 ;
        RECT -61.455 464.030 -54.060 464.380 ;
        RECT -61.455 463.975 -61.095 464.030 ;
        RECT -62.185 463.020 -60.750 463.060 ;
        RECT -62.185 462.850 -57.780 463.020 ;
        RECT -62.185 462.845 -60.750 462.850 ;
        RECT -62.185 462.635 -61.970 462.845 ;
        RECT -54.410 462.690 -54.060 464.030 ;
        RECT -62.385 462.605 -61.970 462.635 ;
        RECT -63.880 462.435 -61.970 462.605 ;
        RECT -62.385 462.415 -61.970 462.435 ;
        RECT -62.170 462.175 -61.970 462.415 ;
        RECT -61.520 461.985 -61.245 462.675 ;
        RECT -55.270 462.520 -54.060 462.690 ;
        RECT -54.115 462.030 -53.575 462.200 ;
        RECT -62.070 461.770 -60.990 461.985 ;
        RECT -57.830 461.960 -57.440 461.990 ;
        RECT -60.820 461.790 -57.440 461.960 ;
        RECT -57.830 461.780 -57.440 461.790 ;
        RECT -62.070 460.440 -61.870 461.770 ;
        RECT -61.185 461.490 -60.990 461.770 ;
        RECT -61.185 461.470 -60.720 461.490 ;
        RECT -61.630 460.560 -61.355 461.335 ;
        RECT -61.185 461.300 -57.780 461.470 ;
        RECT -61.185 461.280 -60.720 461.300 ;
        RECT -61.175 460.980 -60.730 461.005 ;
        RECT -57.610 461.000 -57.440 461.780 ;
        RECT -55.270 461.540 -54.730 461.710 ;
        RECT -54.115 461.050 -53.575 461.220 ;
        RECT -57.820 460.980 -57.440 461.000 ;
        RECT -61.175 460.810 -57.440 460.980 ;
        RECT -61.175 460.795 -60.730 460.810 ;
        RECT -62.420 460.415 -61.870 460.440 ;
        RECT -63.880 460.245 -61.870 460.415 ;
        RECT -62.420 460.215 -61.870 460.245 ;
        RECT -62.170 459.210 -61.895 459.985 ;
        RECT -62.110 459.025 -61.940 459.210 ;
        RECT -61.585 458.885 -61.405 460.560 ;
        RECT -61.175 459.945 -60.995 460.795 ;
        RECT -57.820 460.790 -57.440 460.810 ;
        RECT -55.270 460.560 -54.730 460.730 ;
        RECT -54.560 459.970 -54.260 460.335 ;
        RECT -61.175 459.925 -60.700 459.945 ;
        RECT -61.175 459.755 -57.780 459.925 ;
        RECT -61.175 459.735 -60.700 459.755 ;
        RECT -54.495 459.665 -54.290 459.970 ;
        RECT -54.495 459.610 -53.395 459.665 ;
        RECT -54.495 459.470 -53.355 459.610 ;
        RECT -54.355 459.360 -53.355 459.470 ;
        RECT -59.430 458.885 -59.080 458.915 ;
        RECT -61.595 458.535 -59.080 458.885 ;
        RECT -53.545 458.665 -53.355 459.360 ;
        RECT -53.120 458.925 -52.765 459.295 ;
        RECT -52.580 458.985 -51.040 459.155 ;
        RECT -59.430 457.695 -59.080 458.535 ;
        RECT -55.265 458.495 -53.355 458.665 ;
        RECT -59.430 457.525 -58.220 457.695 ;
        RECT -53.545 457.685 -53.355 458.495 ;
        RECT -55.265 457.515 -53.355 457.685 ;
        RECT -59.915 457.035 -59.375 457.205 ;
        RECT -58.760 456.545 -58.220 456.715 ;
        RECT -53.510 456.600 -53.240 457.275 ;
        RECT -52.990 457.220 -52.795 458.925 ;
        RECT -49.070 458.920 -44.215 459.110 ;
        RECT -52.580 458.495 -51.040 458.665 ;
        RECT -52.580 458.005 -51.040 458.175 ;
        RECT -52.990 456.870 -52.790 457.220 ;
        RECT -52.580 457.025 -51.040 457.195 ;
        RECT -53.000 456.865 -52.790 456.870 ;
        RECT -53.480 456.500 -53.280 456.600 ;
        RECT -59.915 456.055 -59.375 456.225 ;
        RECT -58.760 455.565 -58.220 455.735 ;
        RECT -53.470 455.465 -53.290 456.500 ;
        RECT -59.230 454.975 -58.930 455.340 ;
        RECT -59.200 454.670 -58.995 454.975 ;
        RECT -60.095 454.615 -58.995 454.670 ;
        RECT -60.135 454.475 -58.995 454.615 ;
        RECT -54.620 454.610 -53.580 454.780 ;
        RECT -60.135 454.365 -59.135 454.475 ;
        RECT -62.450 453.990 -60.910 454.160 ;
        RECT -60.725 453.930 -60.370 454.300 ;
        RECT -62.450 453.500 -60.910 453.670 ;
        RECT -62.450 453.010 -60.910 453.180 ;
        RECT -60.695 452.225 -60.500 453.930 ;
        RECT -60.135 453.670 -59.945 454.365 ;
        RECT -53.000 454.290 -52.800 456.865 ;
        RECT -53.000 454.125 -51.930 454.290 ;
        RECT -52.970 454.120 -51.930 454.125 ;
        RECT -60.135 453.500 -58.225 453.670 ;
        RECT -54.620 453.630 -53.580 453.800 ;
        RECT -60.135 452.690 -59.945 453.500 ;
        RECT -52.970 453.140 -51.930 453.310 ;
        RECT -60.135 452.520 -58.225 452.690 ;
        RECT -54.620 452.650 -53.580 452.820 ;
        RECT -62.450 452.030 -60.910 452.200 ;
        RECT -60.700 451.875 -60.500 452.225 ;
        RECT -53.410 452.060 -53.110 452.425 ;
        RECT -60.700 451.870 -60.490 451.875 ;
        RECT -60.690 450.740 -60.490 451.870 ;
        RECT -53.345 451.840 -53.140 452.060 ;
        RECT -53.430 451.705 -52.680 451.840 ;
        RECT -53.680 451.325 -52.680 451.705 ;
        RECT -53.430 451.190 -52.680 451.325 ;
        RECT -53.190 449.045 -52.810 451.190 ;
        RECT -51.230 450.365 -50.960 450.425 ;
        RECT -49.070 450.365 -48.880 458.920 ;
        RECT -44.405 457.840 -44.215 458.920 ;
        RECT -44.655 457.820 -41.565 457.840 ;
        RECT -46.170 457.650 -41.565 457.820 ;
        RECT -43.665 457.075 -43.370 457.345 ;
        RECT -43.625 456.815 -43.455 457.075 ;
        RECT -42.880 456.815 -42.610 457.475 ;
        RECT -41.750 457.340 -41.565 457.650 ;
        RECT -41.750 457.330 -41.100 457.340 ;
        RECT -41.750 457.160 -39.650 457.330 ;
        RECT -41.750 457.155 -41.100 457.160 ;
        RECT -43.650 456.680 -42.220 456.815 ;
        RECT -46.170 456.645 -42.220 456.680 ;
        RECT -46.170 456.510 -43.480 456.645 ;
        RECT -43.650 456.505 -43.480 456.510 ;
        RECT -46.170 456.020 -43.630 456.190 ;
        RECT -43.295 456.185 -42.605 456.455 ;
        RECT -42.390 456.190 -42.220 456.645 ;
        RECT -42.390 456.020 -39.650 456.190 ;
        RECT -42.785 455.135 -42.515 455.825 ;
        RECT -46.170 454.390 -43.475 454.560 ;
        RECT -43.650 453.935 -43.475 454.390 ;
        RECT -43.220 454.260 -42.950 454.950 ;
        RECT -42.740 454.560 -42.570 455.135 ;
        RECT -42.740 454.390 -39.650 454.560 ;
        RECT -46.170 453.765 -43.475 453.935 ;
        RECT -42.740 453.930 -42.570 454.390 ;
        RECT -43.305 453.760 -42.570 453.930 ;
        RECT -39.665 453.910 -39.300 453.915 ;
        RECT -43.305 453.445 -43.135 453.760 ;
        RECT -42.190 453.740 -39.300 453.910 ;
        RECT -46.170 453.275 -43.135 453.445 ;
        RECT -42.945 453.420 -42.155 453.425 ;
        RECT -42.945 453.250 -39.650 453.420 ;
        RECT -42.945 453.235 -42.155 453.250 ;
        RECT -43.985 452.750 -43.295 452.780 ;
        RECT -42.945 452.750 -42.755 453.235 ;
        RECT -39.470 452.930 -39.300 453.740 ;
        RECT -42.190 452.760 -39.300 452.930 ;
        RECT -39.670 452.755 -39.300 452.760 ;
        RECT -43.985 452.560 -42.755 452.750 ;
        RECT -43.985 452.510 -43.295 452.560 ;
        RECT -42.945 451.585 -42.755 452.560 ;
        RECT -39.470 452.510 -39.300 452.755 ;
        RECT -46.170 451.415 -42.755 451.585 ;
        RECT -42.580 452.310 -39.300 452.510 ;
        RECT -42.580 451.585 -42.380 452.310 ;
        RECT -42.580 451.415 -39.650 451.585 ;
        RECT -42.580 451.410 -42.150 451.415 ;
        RECT -43.900 450.510 -43.630 451.200 ;
        RECT -51.230 450.175 -48.880 450.365 ;
        RECT -51.230 450.060 -50.960 450.175 ;
        RECT -44.875 449.820 -44.480 449.880 ;
        RECT -43.845 449.820 -43.675 450.510 ;
        RECT -43.220 450.230 -42.950 450.920 ;
        RECT -44.875 449.485 -43.675 449.820 ;
        RECT -44.525 449.460 -43.675 449.485 ;
        RECT -53.190 448.665 -48.910 449.045 ;
        RECT -62.030 448.240 -60.570 448.455 ;
        RECT -62.030 444.720 -61.815 448.240 ;
        RECT -60.785 447.245 -60.570 448.240 ;
        RECT -50.695 447.245 -50.270 447.375 ;
        RECT -60.785 447.030 -50.270 447.245 ;
        RECT -50.695 446.915 -50.270 447.030 ;
        RECT -61.300 446.040 -60.940 446.160 ;
        RECT -61.300 445.690 -53.905 446.040 ;
        RECT -61.300 445.635 -60.940 445.690 ;
        RECT -62.030 444.680 -60.595 444.720 ;
        RECT -62.030 444.510 -57.625 444.680 ;
        RECT -62.030 444.505 -60.595 444.510 ;
        RECT -62.030 444.295 -61.815 444.505 ;
        RECT -54.255 444.350 -53.905 445.690 ;
        RECT -62.230 444.265 -61.815 444.295 ;
        RECT -63.725 444.095 -61.815 444.265 ;
        RECT -62.230 444.075 -61.815 444.095 ;
        RECT -62.015 443.835 -61.815 444.075 ;
        RECT -61.365 443.645 -61.090 444.335 ;
        RECT -55.115 444.180 -53.905 444.350 ;
        RECT -53.960 443.690 -53.420 443.860 ;
        RECT -61.915 443.430 -60.835 443.645 ;
        RECT -57.675 443.620 -57.285 443.650 ;
        RECT -60.665 443.450 -57.285 443.620 ;
        RECT -57.675 443.440 -57.285 443.450 ;
        RECT -61.915 442.100 -61.715 443.430 ;
        RECT -61.030 443.150 -60.835 443.430 ;
        RECT -61.030 443.130 -60.565 443.150 ;
        RECT -61.475 442.220 -61.200 442.995 ;
        RECT -61.030 442.960 -57.625 443.130 ;
        RECT -61.030 442.940 -60.565 442.960 ;
        RECT -61.020 442.640 -60.575 442.665 ;
        RECT -57.455 442.660 -57.285 443.440 ;
        RECT -55.115 443.200 -54.575 443.370 ;
        RECT -53.960 442.710 -53.420 442.880 ;
        RECT -57.665 442.640 -57.285 442.660 ;
        RECT -61.020 442.470 -57.285 442.640 ;
        RECT -61.020 442.455 -60.575 442.470 ;
        RECT -62.265 442.075 -61.715 442.100 ;
        RECT -63.725 441.905 -61.715 442.075 ;
        RECT -62.265 441.875 -61.715 441.905 ;
        RECT -62.015 440.870 -61.740 441.645 ;
        RECT -61.955 440.685 -61.785 440.870 ;
        RECT -61.430 440.545 -61.250 442.220 ;
        RECT -61.020 441.605 -60.840 442.455 ;
        RECT -57.665 442.450 -57.285 442.470 ;
        RECT -55.115 442.220 -54.575 442.390 ;
        RECT -54.405 441.630 -54.105 441.995 ;
        RECT -61.020 441.585 -60.545 441.605 ;
        RECT -61.020 441.415 -57.625 441.585 ;
        RECT -61.020 441.395 -60.545 441.415 ;
        RECT -54.340 441.325 -54.135 441.630 ;
        RECT -54.340 441.270 -53.240 441.325 ;
        RECT -54.340 441.130 -53.200 441.270 ;
        RECT -54.200 441.020 -53.200 441.130 ;
        RECT -59.275 440.545 -58.925 440.575 ;
        RECT -61.440 440.195 -58.925 440.545 ;
        RECT -53.390 440.325 -53.200 441.020 ;
        RECT -52.965 440.585 -52.610 440.955 ;
        RECT -52.425 440.645 -50.885 440.815 ;
        RECT -59.275 439.355 -58.925 440.195 ;
        RECT -55.110 440.155 -53.200 440.325 ;
        RECT -59.275 439.185 -58.065 439.355 ;
        RECT -53.390 439.345 -53.200 440.155 ;
        RECT -55.110 439.175 -53.200 439.345 ;
        RECT -59.760 438.695 -59.220 438.865 ;
        RECT -58.605 438.205 -58.065 438.375 ;
        RECT -53.355 438.260 -53.085 438.935 ;
        RECT -52.835 438.880 -52.640 440.585 ;
        RECT -52.425 440.155 -50.885 440.325 ;
        RECT -52.425 439.665 -50.885 439.835 ;
        RECT -52.835 438.530 -52.635 438.880 ;
        RECT -52.425 438.685 -50.885 438.855 ;
        RECT -52.845 438.525 -52.635 438.530 ;
        RECT -53.325 438.160 -53.125 438.260 ;
        RECT -59.760 437.715 -59.220 437.885 ;
        RECT -58.605 437.225 -58.065 437.395 ;
        RECT -53.315 437.125 -53.135 438.160 ;
        RECT -59.075 436.635 -58.775 437.000 ;
        RECT -59.045 436.330 -58.840 436.635 ;
        RECT -59.940 436.275 -58.840 436.330 ;
        RECT -59.980 436.135 -58.840 436.275 ;
        RECT -54.465 436.270 -53.425 436.440 ;
        RECT -59.980 436.025 -58.980 436.135 ;
        RECT -62.295 435.650 -60.755 435.820 ;
        RECT -60.570 435.590 -60.215 435.960 ;
        RECT -62.295 435.160 -60.755 435.330 ;
        RECT -62.295 434.670 -60.755 434.840 ;
        RECT -60.540 433.885 -60.345 435.590 ;
        RECT -59.980 435.330 -59.790 436.025 ;
        RECT -52.845 435.950 -52.645 438.525 ;
        RECT -52.845 435.785 -51.775 435.950 ;
        RECT -52.815 435.780 -51.775 435.785 ;
        RECT -59.980 435.160 -58.070 435.330 ;
        RECT -54.465 435.290 -53.425 435.460 ;
        RECT -59.980 434.350 -59.790 435.160 ;
        RECT -52.815 434.800 -51.775 434.970 ;
        RECT -59.980 434.180 -58.070 434.350 ;
        RECT -54.465 434.310 -53.425 434.480 ;
        RECT -62.295 433.690 -60.755 433.860 ;
        RECT -60.545 433.535 -60.345 433.885 ;
        RECT -53.255 433.720 -52.955 434.085 ;
        RECT -60.545 433.530 -60.335 433.535 ;
        RECT -60.535 432.400 -60.335 433.530 ;
        RECT -53.190 433.500 -52.985 433.720 ;
        RECT -53.275 433.205 -52.525 433.500 ;
        RECT -53.275 432.875 -50.200 433.205 ;
        RECT -49.290 432.875 -48.910 448.665 ;
        RECT -43.170 448.495 -43.000 450.230 ;
        RECT -44.765 448.280 -43.000 448.495 ;
        RECT -44.765 444.760 -44.550 448.280 ;
        RECT -44.035 446.080 -43.675 446.200 ;
        RECT -44.035 445.730 -36.640 446.080 ;
        RECT -44.035 445.675 -43.675 445.730 ;
        RECT -44.765 444.720 -43.330 444.760 ;
        RECT -44.765 444.550 -40.360 444.720 ;
        RECT -44.765 444.545 -43.330 444.550 ;
        RECT -44.765 444.335 -44.550 444.545 ;
        RECT -36.990 444.390 -36.640 445.730 ;
        RECT -44.965 444.305 -44.550 444.335 ;
        RECT -46.460 444.135 -44.550 444.305 ;
        RECT -44.965 444.115 -44.550 444.135 ;
        RECT -44.750 443.875 -44.550 444.115 ;
        RECT -44.100 443.685 -43.825 444.375 ;
        RECT -37.850 444.220 -36.640 444.390 ;
        RECT -36.695 443.730 -36.155 443.900 ;
        RECT -44.650 443.470 -43.570 443.685 ;
        RECT -40.410 443.660 -40.020 443.690 ;
        RECT -43.400 443.490 -40.020 443.660 ;
        RECT -40.410 443.480 -40.020 443.490 ;
        RECT -44.650 442.140 -44.450 443.470 ;
        RECT -43.765 443.190 -43.570 443.470 ;
        RECT -43.765 443.170 -43.300 443.190 ;
        RECT -44.210 442.260 -43.935 443.035 ;
        RECT -43.765 443.000 -40.360 443.170 ;
        RECT -43.765 442.980 -43.300 443.000 ;
        RECT -43.755 442.680 -43.310 442.705 ;
        RECT -40.190 442.700 -40.020 443.480 ;
        RECT -37.850 443.240 -37.310 443.410 ;
        RECT -36.695 442.750 -36.155 442.920 ;
        RECT -40.400 442.680 -40.020 442.700 ;
        RECT -43.755 442.510 -40.020 442.680 ;
        RECT -43.755 442.495 -43.310 442.510 ;
        RECT -45.000 442.115 -44.450 442.140 ;
        RECT -46.460 441.945 -44.450 442.115 ;
        RECT -45.000 441.915 -44.450 441.945 ;
        RECT -44.750 440.910 -44.475 441.685 ;
        RECT -44.690 440.725 -44.520 440.910 ;
        RECT -44.165 440.585 -43.985 442.260 ;
        RECT -43.755 441.645 -43.575 442.495 ;
        RECT -40.400 442.490 -40.020 442.510 ;
        RECT -37.850 442.260 -37.310 442.430 ;
        RECT -37.140 441.670 -36.840 442.035 ;
        RECT -43.755 441.625 -43.280 441.645 ;
        RECT -43.755 441.455 -40.360 441.625 ;
        RECT -43.755 441.435 -43.280 441.455 ;
        RECT -37.075 441.365 -36.870 441.670 ;
        RECT -37.075 441.310 -35.975 441.365 ;
        RECT -37.075 441.170 -35.935 441.310 ;
        RECT -36.935 441.060 -35.935 441.170 ;
        RECT -42.010 440.585 -41.660 440.615 ;
        RECT -44.175 440.235 -41.660 440.585 ;
        RECT -36.125 440.365 -35.935 441.060 ;
        RECT -35.700 440.625 -35.345 440.995 ;
        RECT -35.160 440.685 -33.620 440.855 ;
        RECT -42.010 439.395 -41.660 440.235 ;
        RECT -37.845 440.195 -35.935 440.365 ;
        RECT -42.010 439.225 -40.800 439.395 ;
        RECT -36.125 439.385 -35.935 440.195 ;
        RECT -37.845 439.215 -35.935 439.385 ;
        RECT -42.495 438.735 -41.955 438.905 ;
        RECT -41.340 438.245 -40.800 438.415 ;
        RECT -36.090 438.300 -35.820 438.975 ;
        RECT -35.570 438.920 -35.375 440.625 ;
        RECT -35.160 440.195 -33.620 440.365 ;
        RECT -35.160 439.705 -33.620 439.875 ;
        RECT -35.570 438.570 -35.370 438.920 ;
        RECT -35.160 438.725 -33.620 438.895 ;
        RECT -35.580 438.565 -35.370 438.570 ;
        RECT -36.060 438.200 -35.860 438.300 ;
        RECT -42.495 437.755 -41.955 437.925 ;
        RECT -41.340 437.265 -40.800 437.435 ;
        RECT -36.050 437.165 -35.870 438.200 ;
        RECT -41.810 436.675 -41.510 437.040 ;
        RECT -41.780 436.370 -41.575 436.675 ;
        RECT -42.675 436.315 -41.575 436.370 ;
        RECT -42.715 436.175 -41.575 436.315 ;
        RECT -37.200 436.310 -36.160 436.480 ;
        RECT -42.715 436.065 -41.715 436.175 ;
        RECT -45.030 435.690 -43.490 435.860 ;
        RECT -43.305 435.630 -42.950 436.000 ;
        RECT -45.030 435.200 -43.490 435.370 ;
        RECT -45.030 434.710 -43.490 434.880 ;
        RECT -43.275 433.925 -43.080 435.630 ;
        RECT -42.715 435.370 -42.525 436.065 ;
        RECT -35.580 435.990 -35.380 438.565 ;
        RECT -35.580 435.825 -34.510 435.990 ;
        RECT -35.550 435.820 -34.510 435.825 ;
        RECT -42.715 435.200 -40.805 435.370 ;
        RECT -37.200 435.330 -36.160 435.500 ;
        RECT -42.715 434.390 -42.525 435.200 ;
        RECT -35.550 434.840 -34.510 435.010 ;
        RECT -42.715 434.220 -40.805 434.390 ;
        RECT -37.200 434.350 -36.160 434.520 ;
        RECT -45.030 433.730 -43.490 433.900 ;
        RECT -43.280 433.575 -43.080 433.925 ;
        RECT -35.990 433.760 -35.690 434.125 ;
        RECT -43.280 433.570 -43.070 433.575 ;
        RECT -43.270 432.875 -43.070 433.570 ;
        RECT -35.925 433.540 -35.720 433.760 ;
        RECT -36.010 432.890 -35.260 433.540 ;
        RECT -53.275 432.850 -43.070 432.875 ;
        RECT -53.070 432.825 -43.070 432.850 ;
        RECT -50.580 432.495 -43.070 432.825 ;
        RECT -68.870 429.745 -68.035 429.820 ;
        RECT -48.430 429.745 -47.625 432.495 ;
        RECT -43.270 432.440 -43.070 432.495 ;
        RECT -68.870 428.940 -47.625 429.745 ;
        RECT -68.870 428.850 -68.035 428.940 ;
        RECT -34.160 428.830 -33.060 430.060 ;
        RECT -62.355 421.705 -62.140 422.195 ;
        RECT -62.665 420.635 -61.565 421.705 ;
        RECT -34.125 421.695 -33.460 428.830 ;
        RECT -62.355 417.070 -62.140 420.635 ;
        RECT -34.585 420.565 -33.415 421.695 ;
        RECT -61.625 418.390 -61.265 418.510 ;
        RECT -61.625 418.040 -54.230 418.390 ;
        RECT -61.625 417.985 -61.265 418.040 ;
        RECT -62.355 417.030 -60.920 417.070 ;
        RECT -62.355 416.860 -57.950 417.030 ;
        RECT -62.355 416.855 -60.920 416.860 ;
        RECT -62.355 416.645 -62.140 416.855 ;
        RECT -54.580 416.700 -54.230 418.040 ;
        RECT -62.555 416.615 -62.140 416.645 ;
        RECT -64.050 416.445 -62.140 416.615 ;
        RECT -62.555 416.425 -62.140 416.445 ;
        RECT -62.340 416.185 -62.140 416.425 ;
        RECT -61.690 415.995 -61.415 416.685 ;
        RECT -55.440 416.530 -54.230 416.700 ;
        RECT -54.285 416.040 -53.745 416.210 ;
        RECT -62.240 415.780 -61.160 415.995 ;
        RECT -58.000 415.970 -57.610 416.000 ;
        RECT -60.990 415.800 -57.610 415.970 ;
        RECT -58.000 415.790 -57.610 415.800 ;
        RECT -62.240 414.450 -62.040 415.780 ;
        RECT -61.355 415.500 -61.160 415.780 ;
        RECT -61.355 415.480 -60.890 415.500 ;
        RECT -61.800 414.570 -61.525 415.345 ;
        RECT -61.355 415.310 -57.950 415.480 ;
        RECT -61.355 415.290 -60.890 415.310 ;
        RECT -61.345 414.990 -60.900 415.015 ;
        RECT -57.780 415.010 -57.610 415.790 ;
        RECT -55.440 415.550 -54.900 415.720 ;
        RECT -54.285 415.060 -53.745 415.230 ;
        RECT -57.990 414.990 -57.610 415.010 ;
        RECT -61.345 414.820 -57.610 414.990 ;
        RECT -61.345 414.805 -60.900 414.820 ;
        RECT -62.590 414.425 -62.040 414.450 ;
        RECT -64.050 414.255 -62.040 414.425 ;
        RECT -62.590 414.225 -62.040 414.255 ;
        RECT -62.340 413.220 -62.065 413.995 ;
        RECT -62.280 413.035 -62.110 413.220 ;
        RECT -61.755 412.895 -61.575 414.570 ;
        RECT -61.345 413.955 -61.165 414.805 ;
        RECT -57.990 414.800 -57.610 414.820 ;
        RECT -55.440 414.570 -54.900 414.740 ;
        RECT -54.730 413.980 -54.430 414.345 ;
        RECT -61.345 413.935 -60.870 413.955 ;
        RECT -61.345 413.765 -57.950 413.935 ;
        RECT -61.345 413.745 -60.870 413.765 ;
        RECT -54.665 413.675 -54.460 413.980 ;
        RECT -54.665 413.620 -53.565 413.675 ;
        RECT -54.665 413.480 -53.525 413.620 ;
        RECT -54.525 413.370 -53.525 413.480 ;
        RECT -59.600 412.895 -59.250 412.925 ;
        RECT -61.765 412.545 -59.250 412.895 ;
        RECT -53.715 412.675 -53.525 413.370 ;
        RECT -53.290 412.935 -52.935 413.305 ;
        RECT -52.750 412.995 -51.210 413.165 ;
        RECT -59.600 411.705 -59.250 412.545 ;
        RECT -55.435 412.505 -53.525 412.675 ;
        RECT -59.600 411.535 -58.390 411.705 ;
        RECT -53.715 411.695 -53.525 412.505 ;
        RECT -55.435 411.525 -53.525 411.695 ;
        RECT -60.085 411.045 -59.545 411.215 ;
        RECT -58.930 410.555 -58.390 410.725 ;
        RECT -53.680 410.610 -53.410 411.285 ;
        RECT -53.160 411.230 -52.965 412.935 ;
        RECT -49.240 412.930 -44.385 413.120 ;
        RECT -52.750 412.505 -51.210 412.675 ;
        RECT -52.750 412.015 -51.210 412.185 ;
        RECT -53.160 410.880 -52.960 411.230 ;
        RECT -52.750 411.035 -51.210 411.205 ;
        RECT -53.170 410.875 -52.960 410.880 ;
        RECT -53.650 410.510 -53.450 410.610 ;
        RECT -60.085 410.065 -59.545 410.235 ;
        RECT -58.930 409.575 -58.390 409.745 ;
        RECT -53.640 409.475 -53.460 410.510 ;
        RECT -59.400 408.985 -59.100 409.350 ;
        RECT -59.370 408.680 -59.165 408.985 ;
        RECT -60.265 408.625 -59.165 408.680 ;
        RECT -60.305 408.485 -59.165 408.625 ;
        RECT -54.790 408.620 -53.750 408.790 ;
        RECT -60.305 408.375 -59.305 408.485 ;
        RECT -62.620 408.000 -61.080 408.170 ;
        RECT -60.895 407.940 -60.540 408.310 ;
        RECT -62.620 407.510 -61.080 407.680 ;
        RECT -62.620 407.020 -61.080 407.190 ;
        RECT -60.865 406.235 -60.670 407.940 ;
        RECT -60.305 407.680 -60.115 408.375 ;
        RECT -53.170 408.300 -52.970 410.875 ;
        RECT -53.170 408.135 -52.100 408.300 ;
        RECT -53.140 408.130 -52.100 408.135 ;
        RECT -60.305 407.510 -58.395 407.680 ;
        RECT -54.790 407.640 -53.750 407.810 ;
        RECT -60.305 406.700 -60.115 407.510 ;
        RECT -53.140 407.150 -52.100 407.320 ;
        RECT -60.305 406.530 -58.395 406.700 ;
        RECT -54.790 406.660 -53.750 406.830 ;
        RECT -62.620 406.040 -61.080 406.210 ;
        RECT -60.870 405.885 -60.670 406.235 ;
        RECT -53.580 406.070 -53.280 406.435 ;
        RECT -60.870 405.880 -60.660 405.885 ;
        RECT -60.860 404.750 -60.660 405.880 ;
        RECT -53.515 405.850 -53.310 406.070 ;
        RECT -53.600 405.715 -52.850 405.850 ;
        RECT -53.850 405.335 -52.850 405.715 ;
        RECT -53.600 405.200 -52.850 405.335 ;
        RECT -53.360 403.055 -52.980 405.200 ;
        RECT -51.400 404.375 -51.130 404.435 ;
        RECT -49.240 404.375 -49.050 412.930 ;
        RECT -44.575 411.850 -44.385 412.930 ;
        RECT -44.825 411.830 -41.735 411.850 ;
        RECT -46.340 411.660 -41.735 411.830 ;
        RECT -43.835 411.085 -43.540 411.355 ;
        RECT -43.795 410.825 -43.625 411.085 ;
        RECT -43.050 410.825 -42.780 411.485 ;
        RECT -41.920 411.350 -41.735 411.660 ;
        RECT -41.920 411.340 -41.270 411.350 ;
        RECT -41.920 411.170 -39.820 411.340 ;
        RECT -41.920 411.165 -41.270 411.170 ;
        RECT -43.820 410.690 -42.390 410.825 ;
        RECT -46.340 410.655 -42.390 410.690 ;
        RECT -46.340 410.520 -43.650 410.655 ;
        RECT -43.820 410.515 -43.650 410.520 ;
        RECT -46.340 410.030 -43.800 410.200 ;
        RECT -43.465 410.195 -42.775 410.465 ;
        RECT -42.560 410.200 -42.390 410.655 ;
        RECT -42.560 410.030 -39.820 410.200 ;
        RECT -42.955 409.145 -42.685 409.835 ;
        RECT -46.340 408.400 -43.645 408.570 ;
        RECT -43.820 407.945 -43.645 408.400 ;
        RECT -43.390 408.270 -43.120 408.960 ;
        RECT -42.910 408.570 -42.740 409.145 ;
        RECT -42.910 408.400 -39.820 408.570 ;
        RECT -46.340 407.775 -43.645 407.945 ;
        RECT -42.910 407.940 -42.740 408.400 ;
        RECT -43.475 407.770 -42.740 407.940 ;
        RECT -39.835 407.920 -39.470 407.925 ;
        RECT -43.475 407.455 -43.305 407.770 ;
        RECT -42.360 407.750 -39.470 407.920 ;
        RECT -46.340 407.285 -43.305 407.455 ;
        RECT -43.115 407.430 -42.325 407.435 ;
        RECT -43.115 407.260 -39.820 407.430 ;
        RECT -43.115 407.245 -42.325 407.260 ;
        RECT -44.155 406.760 -43.465 406.790 ;
        RECT -43.115 406.760 -42.925 407.245 ;
        RECT -39.640 406.940 -39.470 407.750 ;
        RECT -42.360 406.770 -39.470 406.940 ;
        RECT -39.840 406.765 -39.470 406.770 ;
        RECT -44.155 406.570 -42.925 406.760 ;
        RECT -44.155 406.520 -43.465 406.570 ;
        RECT -43.115 405.595 -42.925 406.570 ;
        RECT -39.640 406.520 -39.470 406.765 ;
        RECT -46.340 405.425 -42.925 405.595 ;
        RECT -42.750 406.320 -39.470 406.520 ;
        RECT -42.750 405.595 -42.550 406.320 ;
        RECT -42.750 405.425 -39.820 405.595 ;
        RECT -42.750 405.420 -42.320 405.425 ;
        RECT -44.070 404.520 -43.800 405.210 ;
        RECT -51.400 404.185 -49.050 404.375 ;
        RECT -51.400 404.070 -51.130 404.185 ;
        RECT -45.045 403.830 -44.650 403.890 ;
        RECT -44.015 403.830 -43.845 404.520 ;
        RECT -43.390 404.240 -43.120 404.930 ;
        RECT -45.045 403.495 -43.845 403.830 ;
        RECT -44.695 403.470 -43.845 403.495 ;
        RECT -53.360 402.675 -49.080 403.055 ;
        RECT -62.200 402.250 -60.740 402.465 ;
        RECT -62.200 398.730 -61.985 402.250 ;
        RECT -60.955 401.255 -60.740 402.250 ;
        RECT -50.865 401.255 -50.440 401.385 ;
        RECT -60.955 401.040 -50.440 401.255 ;
        RECT -50.865 400.925 -50.440 401.040 ;
        RECT -61.470 400.050 -61.110 400.170 ;
        RECT -61.470 399.700 -54.075 400.050 ;
        RECT -61.470 399.645 -61.110 399.700 ;
        RECT -62.200 398.690 -60.765 398.730 ;
        RECT -62.200 398.520 -57.795 398.690 ;
        RECT -62.200 398.515 -60.765 398.520 ;
        RECT -62.200 398.305 -61.985 398.515 ;
        RECT -54.425 398.360 -54.075 399.700 ;
        RECT -62.400 398.275 -61.985 398.305 ;
        RECT -63.895 398.105 -61.985 398.275 ;
        RECT -62.400 398.085 -61.985 398.105 ;
        RECT -62.185 397.845 -61.985 398.085 ;
        RECT -61.535 397.655 -61.260 398.345 ;
        RECT -55.285 398.190 -54.075 398.360 ;
        RECT -54.130 397.700 -53.590 397.870 ;
        RECT -62.085 397.440 -61.005 397.655 ;
        RECT -57.845 397.630 -57.455 397.660 ;
        RECT -60.835 397.460 -57.455 397.630 ;
        RECT -57.845 397.450 -57.455 397.460 ;
        RECT -62.085 396.110 -61.885 397.440 ;
        RECT -61.200 397.160 -61.005 397.440 ;
        RECT -61.200 397.140 -60.735 397.160 ;
        RECT -61.645 396.230 -61.370 397.005 ;
        RECT -61.200 396.970 -57.795 397.140 ;
        RECT -61.200 396.950 -60.735 396.970 ;
        RECT -61.190 396.650 -60.745 396.675 ;
        RECT -57.625 396.670 -57.455 397.450 ;
        RECT -55.285 397.210 -54.745 397.380 ;
        RECT -54.130 396.720 -53.590 396.890 ;
        RECT -57.835 396.650 -57.455 396.670 ;
        RECT -61.190 396.480 -57.455 396.650 ;
        RECT -61.190 396.465 -60.745 396.480 ;
        RECT -62.435 396.085 -61.885 396.110 ;
        RECT -63.895 395.915 -61.885 396.085 ;
        RECT -62.435 395.885 -61.885 395.915 ;
        RECT -62.185 394.880 -61.910 395.655 ;
        RECT -62.125 394.695 -61.955 394.880 ;
        RECT -61.600 394.555 -61.420 396.230 ;
        RECT -61.190 395.615 -61.010 396.465 ;
        RECT -57.835 396.460 -57.455 396.480 ;
        RECT -55.285 396.230 -54.745 396.400 ;
        RECT -54.575 395.640 -54.275 396.005 ;
        RECT -61.190 395.595 -60.715 395.615 ;
        RECT -61.190 395.425 -57.795 395.595 ;
        RECT -61.190 395.405 -60.715 395.425 ;
        RECT -54.510 395.335 -54.305 395.640 ;
        RECT -54.510 395.280 -53.410 395.335 ;
        RECT -54.510 395.140 -53.370 395.280 ;
        RECT -54.370 395.030 -53.370 395.140 ;
        RECT -59.445 394.555 -59.095 394.585 ;
        RECT -61.610 394.205 -59.095 394.555 ;
        RECT -53.560 394.335 -53.370 395.030 ;
        RECT -53.135 394.595 -52.780 394.965 ;
        RECT -52.595 394.655 -51.055 394.825 ;
        RECT -59.445 393.365 -59.095 394.205 ;
        RECT -55.280 394.165 -53.370 394.335 ;
        RECT -59.445 393.195 -58.235 393.365 ;
        RECT -53.560 393.355 -53.370 394.165 ;
        RECT -55.280 393.185 -53.370 393.355 ;
        RECT -59.930 392.705 -59.390 392.875 ;
        RECT -58.775 392.215 -58.235 392.385 ;
        RECT -53.525 392.270 -53.255 392.945 ;
        RECT -53.005 392.890 -52.810 394.595 ;
        RECT -52.595 394.165 -51.055 394.335 ;
        RECT -52.595 393.675 -51.055 393.845 ;
        RECT -53.005 392.540 -52.805 392.890 ;
        RECT -52.595 392.695 -51.055 392.865 ;
        RECT -53.015 392.535 -52.805 392.540 ;
        RECT -53.495 392.170 -53.295 392.270 ;
        RECT -59.930 391.725 -59.390 391.895 ;
        RECT -58.775 391.235 -58.235 391.405 ;
        RECT -53.485 391.135 -53.305 392.170 ;
        RECT -59.245 390.645 -58.945 391.010 ;
        RECT -59.215 390.340 -59.010 390.645 ;
        RECT -60.110 390.285 -59.010 390.340 ;
        RECT -60.150 390.145 -59.010 390.285 ;
        RECT -54.635 390.280 -53.595 390.450 ;
        RECT -60.150 390.035 -59.150 390.145 ;
        RECT -62.465 389.660 -60.925 389.830 ;
        RECT -60.740 389.600 -60.385 389.970 ;
        RECT -62.465 389.170 -60.925 389.340 ;
        RECT -62.465 388.680 -60.925 388.850 ;
        RECT -60.710 387.895 -60.515 389.600 ;
        RECT -60.150 389.340 -59.960 390.035 ;
        RECT -53.015 389.960 -52.815 392.535 ;
        RECT -53.015 389.795 -51.945 389.960 ;
        RECT -52.985 389.790 -51.945 389.795 ;
        RECT -60.150 389.170 -58.240 389.340 ;
        RECT -54.635 389.300 -53.595 389.470 ;
        RECT -60.150 388.360 -59.960 389.170 ;
        RECT -52.985 388.810 -51.945 388.980 ;
        RECT -60.150 388.190 -58.240 388.360 ;
        RECT -54.635 388.320 -53.595 388.490 ;
        RECT -62.465 387.700 -60.925 387.870 ;
        RECT -60.715 387.545 -60.515 387.895 ;
        RECT -53.425 387.730 -53.125 388.095 ;
        RECT -60.715 387.540 -60.505 387.545 ;
        RECT -60.705 386.410 -60.505 387.540 ;
        RECT -53.360 387.510 -53.155 387.730 ;
        RECT -53.445 387.215 -52.695 387.510 ;
        RECT -53.445 386.885 -50.370 387.215 ;
        RECT -49.460 386.885 -49.080 402.675 ;
        RECT -43.340 402.505 -43.170 404.240 ;
        RECT -44.935 402.290 -43.170 402.505 ;
        RECT -44.935 398.770 -44.720 402.290 ;
        RECT -44.205 400.090 -43.845 400.210 ;
        RECT -44.205 399.740 -36.810 400.090 ;
        RECT -44.205 399.685 -43.845 399.740 ;
        RECT -44.935 398.730 -43.500 398.770 ;
        RECT -44.935 398.560 -40.530 398.730 ;
        RECT -44.935 398.555 -43.500 398.560 ;
        RECT -44.935 398.345 -44.720 398.555 ;
        RECT -37.160 398.400 -36.810 399.740 ;
        RECT -45.135 398.315 -44.720 398.345 ;
        RECT -46.630 398.145 -44.720 398.315 ;
        RECT -45.135 398.125 -44.720 398.145 ;
        RECT -44.920 397.885 -44.720 398.125 ;
        RECT -44.270 397.695 -43.995 398.385 ;
        RECT -38.020 398.230 -36.810 398.400 ;
        RECT -36.865 397.740 -36.325 397.910 ;
        RECT -44.820 397.480 -43.740 397.695 ;
        RECT -40.580 397.670 -40.190 397.700 ;
        RECT -43.570 397.500 -40.190 397.670 ;
        RECT -40.580 397.490 -40.190 397.500 ;
        RECT -44.820 396.150 -44.620 397.480 ;
        RECT -43.935 397.200 -43.740 397.480 ;
        RECT -43.935 397.180 -43.470 397.200 ;
        RECT -44.380 396.270 -44.105 397.045 ;
        RECT -43.935 397.010 -40.530 397.180 ;
        RECT -43.935 396.990 -43.470 397.010 ;
        RECT -43.925 396.690 -43.480 396.715 ;
        RECT -40.360 396.710 -40.190 397.490 ;
        RECT -38.020 397.250 -37.480 397.420 ;
        RECT -36.865 396.760 -36.325 396.930 ;
        RECT -40.570 396.690 -40.190 396.710 ;
        RECT -43.925 396.520 -40.190 396.690 ;
        RECT -43.925 396.505 -43.480 396.520 ;
        RECT -45.170 396.125 -44.620 396.150 ;
        RECT -46.630 395.955 -44.620 396.125 ;
        RECT -45.170 395.925 -44.620 395.955 ;
        RECT -44.920 394.920 -44.645 395.695 ;
        RECT -44.860 394.735 -44.690 394.920 ;
        RECT -44.335 394.595 -44.155 396.270 ;
        RECT -43.925 395.655 -43.745 396.505 ;
        RECT -40.570 396.500 -40.190 396.520 ;
        RECT -38.020 396.270 -37.480 396.440 ;
        RECT -37.310 395.680 -37.010 396.045 ;
        RECT -43.925 395.635 -43.450 395.655 ;
        RECT -43.925 395.465 -40.530 395.635 ;
        RECT -43.925 395.445 -43.450 395.465 ;
        RECT -37.245 395.375 -37.040 395.680 ;
        RECT -37.245 395.320 -36.145 395.375 ;
        RECT -37.245 395.180 -36.105 395.320 ;
        RECT -37.105 395.070 -36.105 395.180 ;
        RECT -42.180 394.595 -41.830 394.625 ;
        RECT -44.345 394.245 -41.830 394.595 ;
        RECT -36.295 394.375 -36.105 395.070 ;
        RECT -35.870 394.635 -35.515 395.005 ;
        RECT -35.330 394.695 -33.790 394.865 ;
        RECT -42.180 393.405 -41.830 394.245 ;
        RECT -38.015 394.205 -36.105 394.375 ;
        RECT -42.180 393.235 -40.970 393.405 ;
        RECT -36.295 393.395 -36.105 394.205 ;
        RECT -38.015 393.225 -36.105 393.395 ;
        RECT -42.665 392.745 -42.125 392.915 ;
        RECT -41.510 392.255 -40.970 392.425 ;
        RECT -36.260 392.310 -35.990 392.985 ;
        RECT -35.740 392.930 -35.545 394.635 ;
        RECT -35.330 394.205 -33.790 394.375 ;
        RECT -35.330 393.715 -33.790 393.885 ;
        RECT -35.740 392.580 -35.540 392.930 ;
        RECT -35.330 392.735 -33.790 392.905 ;
        RECT -35.750 392.575 -35.540 392.580 ;
        RECT -36.230 392.210 -36.030 392.310 ;
        RECT -42.665 391.765 -42.125 391.935 ;
        RECT -41.510 391.275 -40.970 391.445 ;
        RECT -36.220 391.175 -36.040 392.210 ;
        RECT -41.980 390.685 -41.680 391.050 ;
        RECT -41.950 390.380 -41.745 390.685 ;
        RECT -42.845 390.325 -41.745 390.380 ;
        RECT -42.885 390.185 -41.745 390.325 ;
        RECT -37.370 390.320 -36.330 390.490 ;
        RECT -42.885 390.075 -41.885 390.185 ;
        RECT -45.200 389.700 -43.660 389.870 ;
        RECT -43.475 389.640 -43.120 390.010 ;
        RECT -45.200 389.210 -43.660 389.380 ;
        RECT -45.200 388.720 -43.660 388.890 ;
        RECT -43.445 387.935 -43.250 389.640 ;
        RECT -42.885 389.380 -42.695 390.075 ;
        RECT -35.750 390.000 -35.550 392.575 ;
        RECT -35.750 389.835 -34.680 390.000 ;
        RECT -35.720 389.830 -34.680 389.835 ;
        RECT -42.885 389.210 -40.975 389.380 ;
        RECT -37.370 389.340 -36.330 389.510 ;
        RECT -42.885 388.400 -42.695 389.210 ;
        RECT -35.720 388.850 -34.680 389.020 ;
        RECT -42.885 388.230 -40.975 388.400 ;
        RECT -37.370 388.360 -36.330 388.530 ;
        RECT -45.200 387.740 -43.660 387.910 ;
        RECT -43.450 387.585 -43.250 387.935 ;
        RECT -36.160 387.770 -35.860 388.135 ;
        RECT -43.450 387.580 -43.240 387.585 ;
        RECT -43.440 386.885 -43.240 387.580 ;
        RECT -36.095 387.550 -35.890 387.770 ;
        RECT -36.180 386.900 -35.430 387.550 ;
        RECT -53.445 386.860 -43.240 386.885 ;
        RECT -53.240 386.835 -43.240 386.860 ;
        RECT -50.750 386.505 -43.240 386.835 ;
        RECT -48.860 383.985 -48.130 386.505 ;
        RECT -43.440 386.450 -43.240 386.505 ;
        RECT -68.865 383.255 -48.130 383.985 ;
        RECT -34.390 383.875 -33.280 385.360 ;
        RECT -62.785 376.245 -61.130 377.930 ;
        RECT -34.280 377.570 -33.445 383.875 ;
        RECT -34.615 376.245 -33.290 377.570 ;
        RECT -69.045 375.865 -67.590 376.035 ;
        RECT -72.945 375.820 -67.590 375.865 ;
        RECT -72.990 374.620 -67.590 375.820 ;
        RECT -72.945 374.535 -67.590 374.620 ;
        RECT -69.045 374.450 -67.590 374.535 ;
        RECT -62.160 372.755 -61.945 376.245 ;
        RECT -61.430 374.075 -61.070 374.195 ;
        RECT -61.430 373.725 -54.035 374.075 ;
        RECT -61.430 373.670 -61.070 373.725 ;
        RECT -62.160 372.715 -60.725 372.755 ;
        RECT -62.160 372.545 -57.755 372.715 ;
        RECT -62.160 372.540 -60.725 372.545 ;
        RECT -62.160 372.330 -61.945 372.540 ;
        RECT -54.385 372.385 -54.035 373.725 ;
        RECT -62.360 372.300 -61.945 372.330 ;
        RECT -63.855 372.130 -61.945 372.300 ;
        RECT -62.360 372.110 -61.945 372.130 ;
        RECT -62.145 371.870 -61.945 372.110 ;
        RECT -61.495 371.680 -61.220 372.370 ;
        RECT -55.245 372.215 -54.035 372.385 ;
        RECT -54.090 371.725 -53.550 371.895 ;
        RECT -62.045 371.465 -60.965 371.680 ;
        RECT -57.805 371.655 -57.415 371.685 ;
        RECT -60.795 371.485 -57.415 371.655 ;
        RECT -57.805 371.475 -57.415 371.485 ;
        RECT -62.045 370.135 -61.845 371.465 ;
        RECT -61.160 371.185 -60.965 371.465 ;
        RECT -61.160 371.165 -60.695 371.185 ;
        RECT -61.605 370.255 -61.330 371.030 ;
        RECT -61.160 370.995 -57.755 371.165 ;
        RECT -61.160 370.975 -60.695 370.995 ;
        RECT -61.150 370.675 -60.705 370.700 ;
        RECT -57.585 370.695 -57.415 371.475 ;
        RECT -55.245 371.235 -54.705 371.405 ;
        RECT -54.090 370.745 -53.550 370.915 ;
        RECT -57.795 370.675 -57.415 370.695 ;
        RECT -61.150 370.505 -57.415 370.675 ;
        RECT -61.150 370.490 -60.705 370.505 ;
        RECT -62.395 370.110 -61.845 370.135 ;
        RECT -63.855 369.940 -61.845 370.110 ;
        RECT -62.395 369.910 -61.845 369.940 ;
        RECT -62.145 368.905 -61.870 369.680 ;
        RECT -62.085 368.720 -61.915 368.905 ;
        RECT -61.560 368.580 -61.380 370.255 ;
        RECT -61.150 369.640 -60.970 370.490 ;
        RECT -57.795 370.485 -57.415 370.505 ;
        RECT -55.245 370.255 -54.705 370.425 ;
        RECT -54.535 369.665 -54.235 370.030 ;
        RECT -61.150 369.620 -60.675 369.640 ;
        RECT -61.150 369.450 -57.755 369.620 ;
        RECT -61.150 369.430 -60.675 369.450 ;
        RECT -54.470 369.360 -54.265 369.665 ;
        RECT -54.470 369.305 -53.370 369.360 ;
        RECT -54.470 369.165 -53.330 369.305 ;
        RECT -54.330 369.055 -53.330 369.165 ;
        RECT -59.405 368.580 -59.055 368.610 ;
        RECT -61.570 368.230 -59.055 368.580 ;
        RECT -53.520 368.360 -53.330 369.055 ;
        RECT -53.095 368.620 -52.740 368.990 ;
        RECT -52.555 368.680 -51.015 368.850 ;
        RECT -59.405 367.390 -59.055 368.230 ;
        RECT -55.240 368.190 -53.330 368.360 ;
        RECT -59.405 367.220 -58.195 367.390 ;
        RECT -53.520 367.380 -53.330 368.190 ;
        RECT -55.240 367.210 -53.330 367.380 ;
        RECT -59.890 366.730 -59.350 366.900 ;
        RECT -58.735 366.240 -58.195 366.410 ;
        RECT -53.485 366.295 -53.215 366.970 ;
        RECT -52.965 366.915 -52.770 368.620 ;
        RECT -49.045 368.615 -44.190 368.805 ;
        RECT -52.555 368.190 -51.015 368.360 ;
        RECT -52.555 367.700 -51.015 367.870 ;
        RECT -52.965 366.565 -52.765 366.915 ;
        RECT -52.555 366.720 -51.015 366.890 ;
        RECT -52.975 366.560 -52.765 366.565 ;
        RECT -53.455 366.195 -53.255 366.295 ;
        RECT -59.890 365.750 -59.350 365.920 ;
        RECT -58.735 365.260 -58.195 365.430 ;
        RECT -53.445 365.160 -53.265 366.195 ;
        RECT -59.205 364.670 -58.905 365.035 ;
        RECT -59.175 364.365 -58.970 364.670 ;
        RECT -60.070 364.310 -58.970 364.365 ;
        RECT -60.110 364.170 -58.970 364.310 ;
        RECT -54.595 364.305 -53.555 364.475 ;
        RECT -60.110 364.060 -59.110 364.170 ;
        RECT -62.425 363.685 -60.885 363.855 ;
        RECT -60.700 363.625 -60.345 363.995 ;
        RECT -62.425 363.195 -60.885 363.365 ;
        RECT -62.425 362.705 -60.885 362.875 ;
        RECT -60.670 361.920 -60.475 363.625 ;
        RECT -60.110 363.365 -59.920 364.060 ;
        RECT -52.975 363.985 -52.775 366.560 ;
        RECT -52.975 363.820 -51.905 363.985 ;
        RECT -52.945 363.815 -51.905 363.820 ;
        RECT -60.110 363.195 -58.200 363.365 ;
        RECT -54.595 363.325 -53.555 363.495 ;
        RECT -60.110 362.385 -59.920 363.195 ;
        RECT -52.945 362.835 -51.905 363.005 ;
        RECT -60.110 362.215 -58.200 362.385 ;
        RECT -54.595 362.345 -53.555 362.515 ;
        RECT -62.425 361.725 -60.885 361.895 ;
        RECT -60.675 361.570 -60.475 361.920 ;
        RECT -53.385 361.755 -53.085 362.120 ;
        RECT -60.675 361.565 -60.465 361.570 ;
        RECT -60.665 360.435 -60.465 361.565 ;
        RECT -53.320 361.535 -53.115 361.755 ;
        RECT -53.405 361.400 -52.655 361.535 ;
        RECT -53.655 361.020 -52.655 361.400 ;
        RECT -53.405 360.885 -52.655 361.020 ;
        RECT -53.165 358.740 -52.785 360.885 ;
        RECT -51.205 360.060 -50.935 360.120 ;
        RECT -49.045 360.060 -48.855 368.615 ;
        RECT -44.380 367.535 -44.190 368.615 ;
        RECT -44.630 367.515 -41.540 367.535 ;
        RECT -46.145 367.345 -41.540 367.515 ;
        RECT -43.640 366.770 -43.345 367.040 ;
        RECT -43.600 366.510 -43.430 366.770 ;
        RECT -42.855 366.510 -42.585 367.170 ;
        RECT -41.725 367.035 -41.540 367.345 ;
        RECT -41.725 367.025 -41.075 367.035 ;
        RECT -41.725 366.855 -39.625 367.025 ;
        RECT -41.725 366.850 -41.075 366.855 ;
        RECT -43.625 366.375 -42.195 366.510 ;
        RECT -46.145 366.340 -42.195 366.375 ;
        RECT -46.145 366.205 -43.455 366.340 ;
        RECT -43.625 366.200 -43.455 366.205 ;
        RECT -46.145 365.715 -43.605 365.885 ;
        RECT -43.270 365.880 -42.580 366.150 ;
        RECT -42.365 365.885 -42.195 366.340 ;
        RECT -42.365 365.715 -39.625 365.885 ;
        RECT -42.760 364.830 -42.490 365.520 ;
        RECT -46.145 364.085 -43.450 364.255 ;
        RECT -43.625 363.630 -43.450 364.085 ;
        RECT -43.195 363.955 -42.925 364.645 ;
        RECT -42.715 364.255 -42.545 364.830 ;
        RECT -42.715 364.085 -39.625 364.255 ;
        RECT -46.145 363.460 -43.450 363.630 ;
        RECT -42.715 363.625 -42.545 364.085 ;
        RECT -43.280 363.455 -42.545 363.625 ;
        RECT -39.640 363.605 -39.275 363.610 ;
        RECT -43.280 363.140 -43.110 363.455 ;
        RECT -42.165 363.435 -39.275 363.605 ;
        RECT -46.145 362.970 -43.110 363.140 ;
        RECT -42.920 363.115 -42.130 363.120 ;
        RECT -42.920 362.945 -39.625 363.115 ;
        RECT -42.920 362.930 -42.130 362.945 ;
        RECT -43.960 362.445 -43.270 362.475 ;
        RECT -42.920 362.445 -42.730 362.930 ;
        RECT -39.445 362.625 -39.275 363.435 ;
        RECT -42.165 362.455 -39.275 362.625 ;
        RECT -39.645 362.450 -39.275 362.455 ;
        RECT -43.960 362.255 -42.730 362.445 ;
        RECT -43.960 362.205 -43.270 362.255 ;
        RECT -42.920 361.280 -42.730 362.255 ;
        RECT -39.445 362.205 -39.275 362.450 ;
        RECT -46.145 361.110 -42.730 361.280 ;
        RECT -42.555 362.005 -39.275 362.205 ;
        RECT -42.555 361.280 -42.355 362.005 ;
        RECT -42.555 361.110 -39.625 361.280 ;
        RECT -42.555 361.105 -42.125 361.110 ;
        RECT -43.875 360.205 -43.605 360.895 ;
        RECT -51.205 359.870 -48.855 360.060 ;
        RECT -51.205 359.755 -50.935 359.870 ;
        RECT -44.850 359.515 -44.455 359.575 ;
        RECT -43.820 359.515 -43.650 360.205 ;
        RECT -43.195 359.925 -42.925 360.615 ;
        RECT -44.850 359.180 -43.650 359.515 ;
        RECT -44.500 359.155 -43.650 359.180 ;
        RECT -53.165 358.360 -48.885 358.740 ;
        RECT -62.005 357.935 -60.545 358.150 ;
        RECT -62.005 354.415 -61.790 357.935 ;
        RECT -60.760 356.940 -60.545 357.935 ;
        RECT -50.670 356.940 -50.245 357.070 ;
        RECT -60.760 356.725 -50.245 356.940 ;
        RECT -50.670 356.610 -50.245 356.725 ;
        RECT -61.275 355.735 -60.915 355.855 ;
        RECT -61.275 355.385 -53.880 355.735 ;
        RECT -61.275 355.330 -60.915 355.385 ;
        RECT -62.005 354.375 -60.570 354.415 ;
        RECT -62.005 354.205 -57.600 354.375 ;
        RECT -62.005 354.200 -60.570 354.205 ;
        RECT -62.005 353.990 -61.790 354.200 ;
        RECT -54.230 354.045 -53.880 355.385 ;
        RECT -62.205 353.960 -61.790 353.990 ;
        RECT -63.700 353.790 -61.790 353.960 ;
        RECT -62.205 353.770 -61.790 353.790 ;
        RECT -61.990 353.530 -61.790 353.770 ;
        RECT -61.340 353.340 -61.065 354.030 ;
        RECT -55.090 353.875 -53.880 354.045 ;
        RECT -53.935 353.385 -53.395 353.555 ;
        RECT -61.890 353.125 -60.810 353.340 ;
        RECT -57.650 353.315 -57.260 353.345 ;
        RECT -60.640 353.145 -57.260 353.315 ;
        RECT -57.650 353.135 -57.260 353.145 ;
        RECT -61.890 351.795 -61.690 353.125 ;
        RECT -61.005 352.845 -60.810 353.125 ;
        RECT -61.005 352.825 -60.540 352.845 ;
        RECT -61.450 351.915 -61.175 352.690 ;
        RECT -61.005 352.655 -57.600 352.825 ;
        RECT -61.005 352.635 -60.540 352.655 ;
        RECT -60.995 352.335 -60.550 352.360 ;
        RECT -57.430 352.355 -57.260 353.135 ;
        RECT -55.090 352.895 -54.550 353.065 ;
        RECT -53.935 352.405 -53.395 352.575 ;
        RECT -57.640 352.335 -57.260 352.355 ;
        RECT -60.995 352.165 -57.260 352.335 ;
        RECT -60.995 352.150 -60.550 352.165 ;
        RECT -62.240 351.770 -61.690 351.795 ;
        RECT -63.700 351.600 -61.690 351.770 ;
        RECT -62.240 351.570 -61.690 351.600 ;
        RECT -61.990 350.565 -61.715 351.340 ;
        RECT -61.930 350.380 -61.760 350.565 ;
        RECT -61.405 350.240 -61.225 351.915 ;
        RECT -60.995 351.300 -60.815 352.150 ;
        RECT -57.640 352.145 -57.260 352.165 ;
        RECT -55.090 351.915 -54.550 352.085 ;
        RECT -54.380 351.325 -54.080 351.690 ;
        RECT -60.995 351.280 -60.520 351.300 ;
        RECT -60.995 351.110 -57.600 351.280 ;
        RECT -60.995 351.090 -60.520 351.110 ;
        RECT -54.315 351.020 -54.110 351.325 ;
        RECT -54.315 350.965 -53.215 351.020 ;
        RECT -54.315 350.825 -53.175 350.965 ;
        RECT -54.175 350.715 -53.175 350.825 ;
        RECT -59.250 350.240 -58.900 350.270 ;
        RECT -61.415 349.890 -58.900 350.240 ;
        RECT -53.365 350.020 -53.175 350.715 ;
        RECT -52.940 350.280 -52.585 350.650 ;
        RECT -52.400 350.340 -50.860 350.510 ;
        RECT -59.250 349.050 -58.900 349.890 ;
        RECT -55.085 349.850 -53.175 350.020 ;
        RECT -59.250 348.880 -58.040 349.050 ;
        RECT -53.365 349.040 -53.175 349.850 ;
        RECT -55.085 348.870 -53.175 349.040 ;
        RECT -59.735 348.390 -59.195 348.560 ;
        RECT -58.580 347.900 -58.040 348.070 ;
        RECT -53.330 347.955 -53.060 348.630 ;
        RECT -52.810 348.575 -52.615 350.280 ;
        RECT -52.400 349.850 -50.860 350.020 ;
        RECT -52.400 349.360 -50.860 349.530 ;
        RECT -52.810 348.225 -52.610 348.575 ;
        RECT -52.400 348.380 -50.860 348.550 ;
        RECT -52.820 348.220 -52.610 348.225 ;
        RECT -53.300 347.855 -53.100 347.955 ;
        RECT -59.735 347.410 -59.195 347.580 ;
        RECT -58.580 346.920 -58.040 347.090 ;
        RECT -53.290 346.820 -53.110 347.855 ;
        RECT -59.050 346.330 -58.750 346.695 ;
        RECT -59.020 346.025 -58.815 346.330 ;
        RECT -59.915 345.970 -58.815 346.025 ;
        RECT -59.955 345.830 -58.815 345.970 ;
        RECT -54.440 345.965 -53.400 346.135 ;
        RECT -59.955 345.720 -58.955 345.830 ;
        RECT -62.270 345.345 -60.730 345.515 ;
        RECT -60.545 345.285 -60.190 345.655 ;
        RECT -62.270 344.855 -60.730 345.025 ;
        RECT -62.270 344.365 -60.730 344.535 ;
        RECT -60.515 343.580 -60.320 345.285 ;
        RECT -59.955 345.025 -59.765 345.720 ;
        RECT -52.820 345.645 -52.620 348.220 ;
        RECT -52.820 345.480 -51.750 345.645 ;
        RECT -52.790 345.475 -51.750 345.480 ;
        RECT -59.955 344.855 -58.045 345.025 ;
        RECT -54.440 344.985 -53.400 345.155 ;
        RECT -59.955 344.045 -59.765 344.855 ;
        RECT -52.790 344.495 -51.750 344.665 ;
        RECT -59.955 343.875 -58.045 344.045 ;
        RECT -54.440 344.005 -53.400 344.175 ;
        RECT -62.270 343.385 -60.730 343.555 ;
        RECT -60.520 343.230 -60.320 343.580 ;
        RECT -53.230 343.415 -52.930 343.780 ;
        RECT -60.520 343.225 -60.310 343.230 ;
        RECT -60.510 342.095 -60.310 343.225 ;
        RECT -53.165 343.195 -52.960 343.415 ;
        RECT -53.250 342.900 -52.500 343.195 ;
        RECT -53.250 342.570 -50.175 342.900 ;
        RECT -49.265 342.570 -48.885 358.360 ;
        RECT -43.145 358.190 -42.975 359.925 ;
        RECT -44.740 357.975 -42.975 358.190 ;
        RECT -44.740 354.455 -44.525 357.975 ;
        RECT -44.010 355.775 -43.650 355.895 ;
        RECT -44.010 355.425 -36.615 355.775 ;
        RECT -44.010 355.370 -43.650 355.425 ;
        RECT -44.740 354.415 -43.305 354.455 ;
        RECT -44.740 354.245 -40.335 354.415 ;
        RECT -44.740 354.240 -43.305 354.245 ;
        RECT -44.740 354.030 -44.525 354.240 ;
        RECT -36.965 354.085 -36.615 355.425 ;
        RECT -44.940 354.000 -44.525 354.030 ;
        RECT -46.435 353.830 -44.525 354.000 ;
        RECT -44.940 353.810 -44.525 353.830 ;
        RECT -44.725 353.570 -44.525 353.810 ;
        RECT -44.075 353.380 -43.800 354.070 ;
        RECT -37.825 353.915 -36.615 354.085 ;
        RECT -36.670 353.425 -36.130 353.595 ;
        RECT -44.625 353.165 -43.545 353.380 ;
        RECT -40.385 353.355 -39.995 353.385 ;
        RECT -43.375 353.185 -39.995 353.355 ;
        RECT -40.385 353.175 -39.995 353.185 ;
        RECT -44.625 351.835 -44.425 353.165 ;
        RECT -43.740 352.885 -43.545 353.165 ;
        RECT -43.740 352.865 -43.275 352.885 ;
        RECT -44.185 351.955 -43.910 352.730 ;
        RECT -43.740 352.695 -40.335 352.865 ;
        RECT -43.740 352.675 -43.275 352.695 ;
        RECT -43.730 352.375 -43.285 352.400 ;
        RECT -40.165 352.395 -39.995 353.175 ;
        RECT -37.825 352.935 -37.285 353.105 ;
        RECT -36.670 352.445 -36.130 352.615 ;
        RECT -40.375 352.375 -39.995 352.395 ;
        RECT -43.730 352.205 -39.995 352.375 ;
        RECT -43.730 352.190 -43.285 352.205 ;
        RECT -44.975 351.810 -44.425 351.835 ;
        RECT -46.435 351.640 -44.425 351.810 ;
        RECT -44.975 351.610 -44.425 351.640 ;
        RECT -44.725 350.605 -44.450 351.380 ;
        RECT -44.665 350.420 -44.495 350.605 ;
        RECT -44.140 350.280 -43.960 351.955 ;
        RECT -43.730 351.340 -43.550 352.190 ;
        RECT -40.375 352.185 -39.995 352.205 ;
        RECT -37.825 351.955 -37.285 352.125 ;
        RECT -37.115 351.365 -36.815 351.730 ;
        RECT -43.730 351.320 -43.255 351.340 ;
        RECT -43.730 351.150 -40.335 351.320 ;
        RECT -43.730 351.130 -43.255 351.150 ;
        RECT -37.050 351.060 -36.845 351.365 ;
        RECT -37.050 351.005 -35.950 351.060 ;
        RECT -37.050 350.865 -35.910 351.005 ;
        RECT -36.910 350.755 -35.910 350.865 ;
        RECT -41.985 350.280 -41.635 350.310 ;
        RECT -44.150 349.930 -41.635 350.280 ;
        RECT -36.100 350.060 -35.910 350.755 ;
        RECT -35.675 350.320 -35.320 350.690 ;
        RECT -35.135 350.380 -33.595 350.550 ;
        RECT -41.985 349.090 -41.635 349.930 ;
        RECT -37.820 349.890 -35.910 350.060 ;
        RECT -41.985 348.920 -40.775 349.090 ;
        RECT -36.100 349.080 -35.910 349.890 ;
        RECT -37.820 348.910 -35.910 349.080 ;
        RECT -42.470 348.430 -41.930 348.600 ;
        RECT -41.315 347.940 -40.775 348.110 ;
        RECT -36.065 347.995 -35.795 348.670 ;
        RECT -35.545 348.615 -35.350 350.320 ;
        RECT -35.135 349.890 -33.595 350.060 ;
        RECT -35.135 349.400 -33.595 349.570 ;
        RECT -35.545 348.265 -35.345 348.615 ;
        RECT -35.135 348.420 -33.595 348.590 ;
        RECT -35.555 348.260 -35.345 348.265 ;
        RECT -36.035 347.895 -35.835 347.995 ;
        RECT -42.470 347.450 -41.930 347.620 ;
        RECT -41.315 346.960 -40.775 347.130 ;
        RECT -36.025 346.860 -35.845 347.895 ;
        RECT -41.785 346.370 -41.485 346.735 ;
        RECT -41.755 346.065 -41.550 346.370 ;
        RECT -42.650 346.010 -41.550 346.065 ;
        RECT -42.690 345.870 -41.550 346.010 ;
        RECT -37.175 346.005 -36.135 346.175 ;
        RECT -42.690 345.760 -41.690 345.870 ;
        RECT -45.005 345.385 -43.465 345.555 ;
        RECT -43.280 345.325 -42.925 345.695 ;
        RECT -45.005 344.895 -43.465 345.065 ;
        RECT -45.005 344.405 -43.465 344.575 ;
        RECT -43.250 343.620 -43.055 345.325 ;
        RECT -42.690 345.065 -42.500 345.760 ;
        RECT -35.555 345.685 -35.355 348.260 ;
        RECT -35.555 345.520 -34.485 345.685 ;
        RECT -35.525 345.515 -34.485 345.520 ;
        RECT -42.690 344.895 -40.780 345.065 ;
        RECT -37.175 345.025 -36.135 345.195 ;
        RECT -42.690 344.085 -42.500 344.895 ;
        RECT -35.525 344.535 -34.485 344.705 ;
        RECT -42.690 343.915 -40.780 344.085 ;
        RECT -37.175 344.045 -36.135 344.215 ;
        RECT -45.005 343.425 -43.465 343.595 ;
        RECT -43.255 343.270 -43.055 343.620 ;
        RECT -35.965 343.455 -35.665 343.820 ;
        RECT -43.255 343.265 -43.045 343.270 ;
        RECT -43.245 342.570 -43.045 343.265 ;
        RECT -35.900 343.235 -35.695 343.455 ;
        RECT -35.985 342.585 -35.235 343.235 ;
        RECT -53.250 342.545 -43.045 342.570 ;
        RECT -53.045 342.520 -43.045 342.545 ;
        RECT -50.555 342.190 -43.045 342.520 ;
        RECT -68.875 339.640 -68.140 339.810 ;
        RECT -48.225 339.640 -47.495 342.190 ;
        RECT -43.245 342.135 -43.045 342.190 ;
        RECT -68.875 338.910 -47.495 339.640 ;
        RECT -34.170 339.355 -32.835 341.140 ;
        RECT -68.875 338.795 -68.140 338.910 ;
        RECT -62.105 335.115 -61.890 335.680 ;
        RECT -33.945 335.250 -33.000 339.355 ;
        RECT -62.290 334.000 -61.440 335.115 ;
        RECT -62.105 330.555 -61.890 334.000 ;
        RECT -34.000 333.465 -32.665 335.250 ;
        RECT -61.375 331.875 -61.015 331.995 ;
        RECT -61.375 331.525 -53.980 331.875 ;
        RECT -61.375 331.470 -61.015 331.525 ;
        RECT -62.105 330.515 -60.670 330.555 ;
        RECT -62.105 330.345 -57.700 330.515 ;
        RECT -62.105 330.340 -60.670 330.345 ;
        RECT -62.105 330.130 -61.890 330.340 ;
        RECT -54.330 330.185 -53.980 331.525 ;
        RECT -62.305 330.100 -61.890 330.130 ;
        RECT -63.800 329.930 -61.890 330.100 ;
        RECT -62.305 329.910 -61.890 329.930 ;
        RECT -62.090 329.670 -61.890 329.910 ;
        RECT -61.440 329.480 -61.165 330.170 ;
        RECT -55.190 330.015 -53.980 330.185 ;
        RECT -54.035 329.525 -53.495 329.695 ;
        RECT -61.990 329.265 -60.910 329.480 ;
        RECT -57.750 329.455 -57.360 329.485 ;
        RECT -60.740 329.285 -57.360 329.455 ;
        RECT -57.750 329.275 -57.360 329.285 ;
        RECT -61.990 327.935 -61.790 329.265 ;
        RECT -61.105 328.985 -60.910 329.265 ;
        RECT -61.105 328.965 -60.640 328.985 ;
        RECT -61.550 328.055 -61.275 328.830 ;
        RECT -61.105 328.795 -57.700 328.965 ;
        RECT -61.105 328.775 -60.640 328.795 ;
        RECT -61.095 328.475 -60.650 328.500 ;
        RECT -57.530 328.495 -57.360 329.275 ;
        RECT -55.190 329.035 -54.650 329.205 ;
        RECT -54.035 328.545 -53.495 328.715 ;
        RECT -57.740 328.475 -57.360 328.495 ;
        RECT -61.095 328.305 -57.360 328.475 ;
        RECT -61.095 328.290 -60.650 328.305 ;
        RECT -62.340 327.910 -61.790 327.935 ;
        RECT -63.800 327.740 -61.790 327.910 ;
        RECT -62.340 327.710 -61.790 327.740 ;
        RECT -62.090 326.705 -61.815 327.480 ;
        RECT -62.030 326.520 -61.860 326.705 ;
        RECT -61.505 326.380 -61.325 328.055 ;
        RECT -61.095 327.440 -60.915 328.290 ;
        RECT -57.740 328.285 -57.360 328.305 ;
        RECT -55.190 328.055 -54.650 328.225 ;
        RECT -54.480 327.465 -54.180 327.830 ;
        RECT -61.095 327.420 -60.620 327.440 ;
        RECT -61.095 327.250 -57.700 327.420 ;
        RECT -61.095 327.230 -60.620 327.250 ;
        RECT -54.415 327.160 -54.210 327.465 ;
        RECT -54.415 327.105 -53.315 327.160 ;
        RECT -54.415 326.965 -53.275 327.105 ;
        RECT -54.275 326.855 -53.275 326.965 ;
        RECT -59.350 326.380 -59.000 326.410 ;
        RECT -61.515 326.030 -59.000 326.380 ;
        RECT -53.465 326.160 -53.275 326.855 ;
        RECT -53.040 326.420 -52.685 326.790 ;
        RECT -52.500 326.480 -50.960 326.650 ;
        RECT -59.350 325.190 -59.000 326.030 ;
        RECT -55.185 325.990 -53.275 326.160 ;
        RECT -59.350 325.020 -58.140 325.190 ;
        RECT -53.465 325.180 -53.275 325.990 ;
        RECT -55.185 325.010 -53.275 325.180 ;
        RECT -59.835 324.530 -59.295 324.700 ;
        RECT -58.680 324.040 -58.140 324.210 ;
        RECT -53.430 324.095 -53.160 324.770 ;
        RECT -52.910 324.715 -52.715 326.420 ;
        RECT -48.990 326.415 -44.135 326.605 ;
        RECT -52.500 325.990 -50.960 326.160 ;
        RECT -52.500 325.500 -50.960 325.670 ;
        RECT -52.910 324.365 -52.710 324.715 ;
        RECT -52.500 324.520 -50.960 324.690 ;
        RECT -52.920 324.360 -52.710 324.365 ;
        RECT -53.400 323.995 -53.200 324.095 ;
        RECT -59.835 323.550 -59.295 323.720 ;
        RECT -58.680 323.060 -58.140 323.230 ;
        RECT -53.390 322.960 -53.210 323.995 ;
        RECT -59.150 322.470 -58.850 322.835 ;
        RECT -59.120 322.165 -58.915 322.470 ;
        RECT -60.015 322.110 -58.915 322.165 ;
        RECT -60.055 321.970 -58.915 322.110 ;
        RECT -54.540 322.105 -53.500 322.275 ;
        RECT -60.055 321.860 -59.055 321.970 ;
        RECT -62.370 321.485 -60.830 321.655 ;
        RECT -60.645 321.425 -60.290 321.795 ;
        RECT -62.370 320.995 -60.830 321.165 ;
        RECT -62.370 320.505 -60.830 320.675 ;
        RECT -60.615 319.720 -60.420 321.425 ;
        RECT -60.055 321.165 -59.865 321.860 ;
        RECT -52.920 321.785 -52.720 324.360 ;
        RECT -52.920 321.620 -51.850 321.785 ;
        RECT -52.890 321.615 -51.850 321.620 ;
        RECT -60.055 320.995 -58.145 321.165 ;
        RECT -54.540 321.125 -53.500 321.295 ;
        RECT -60.055 320.185 -59.865 320.995 ;
        RECT -52.890 320.635 -51.850 320.805 ;
        RECT -60.055 320.015 -58.145 320.185 ;
        RECT -54.540 320.145 -53.500 320.315 ;
        RECT -62.370 319.525 -60.830 319.695 ;
        RECT -60.620 319.370 -60.420 319.720 ;
        RECT -53.330 319.555 -53.030 319.920 ;
        RECT -60.620 319.365 -60.410 319.370 ;
        RECT -60.610 318.235 -60.410 319.365 ;
        RECT -53.265 319.335 -53.060 319.555 ;
        RECT -53.350 319.200 -52.600 319.335 ;
        RECT -53.600 318.820 -52.600 319.200 ;
        RECT -53.350 318.685 -52.600 318.820 ;
        RECT -53.110 316.540 -52.730 318.685 ;
        RECT -51.150 317.860 -50.880 317.920 ;
        RECT -48.990 317.860 -48.800 326.415 ;
        RECT -44.325 325.335 -44.135 326.415 ;
        RECT -44.575 325.315 -41.485 325.335 ;
        RECT -46.090 325.145 -41.485 325.315 ;
        RECT -43.585 324.570 -43.290 324.840 ;
        RECT -43.545 324.310 -43.375 324.570 ;
        RECT -42.800 324.310 -42.530 324.970 ;
        RECT -41.670 324.835 -41.485 325.145 ;
        RECT -41.670 324.825 -41.020 324.835 ;
        RECT -41.670 324.655 -39.570 324.825 ;
        RECT -41.670 324.650 -41.020 324.655 ;
        RECT -43.570 324.175 -42.140 324.310 ;
        RECT -46.090 324.140 -42.140 324.175 ;
        RECT -46.090 324.005 -43.400 324.140 ;
        RECT -43.570 324.000 -43.400 324.005 ;
        RECT -46.090 323.515 -43.550 323.685 ;
        RECT -43.215 323.680 -42.525 323.950 ;
        RECT -42.310 323.685 -42.140 324.140 ;
        RECT -42.310 323.515 -39.570 323.685 ;
        RECT -42.705 322.630 -42.435 323.320 ;
        RECT -46.090 321.885 -43.395 322.055 ;
        RECT -43.570 321.430 -43.395 321.885 ;
        RECT -43.140 321.755 -42.870 322.445 ;
        RECT -42.660 322.055 -42.490 322.630 ;
        RECT -42.660 321.885 -39.570 322.055 ;
        RECT -46.090 321.260 -43.395 321.430 ;
        RECT -42.660 321.425 -42.490 321.885 ;
        RECT -43.225 321.255 -42.490 321.425 ;
        RECT -39.585 321.405 -39.220 321.410 ;
        RECT -43.225 320.940 -43.055 321.255 ;
        RECT -42.110 321.235 -39.220 321.405 ;
        RECT -46.090 320.770 -43.055 320.940 ;
        RECT -42.865 320.915 -42.075 320.920 ;
        RECT -42.865 320.745 -39.570 320.915 ;
        RECT -42.865 320.730 -42.075 320.745 ;
        RECT -43.905 320.245 -43.215 320.275 ;
        RECT -42.865 320.245 -42.675 320.730 ;
        RECT -39.390 320.425 -39.220 321.235 ;
        RECT -42.110 320.255 -39.220 320.425 ;
        RECT -39.590 320.250 -39.220 320.255 ;
        RECT -43.905 320.055 -42.675 320.245 ;
        RECT -43.905 320.005 -43.215 320.055 ;
        RECT -42.865 319.080 -42.675 320.055 ;
        RECT -39.390 320.005 -39.220 320.250 ;
        RECT -46.090 318.910 -42.675 319.080 ;
        RECT -42.500 319.805 -39.220 320.005 ;
        RECT -42.500 319.080 -42.300 319.805 ;
        RECT -42.500 318.910 -39.570 319.080 ;
        RECT -42.500 318.905 -42.070 318.910 ;
        RECT -43.820 318.005 -43.550 318.695 ;
        RECT -51.150 317.670 -48.800 317.860 ;
        RECT -51.150 317.555 -50.880 317.670 ;
        RECT -44.795 317.315 -44.400 317.375 ;
        RECT -43.765 317.315 -43.595 318.005 ;
        RECT -43.140 317.725 -42.870 318.415 ;
        RECT -44.795 316.980 -43.595 317.315 ;
        RECT -44.445 316.955 -43.595 316.980 ;
        RECT -53.110 316.160 -48.830 316.540 ;
        RECT -61.950 315.735 -60.490 315.950 ;
        RECT -61.950 312.215 -61.735 315.735 ;
        RECT -60.705 314.740 -60.490 315.735 ;
        RECT -50.615 314.740 -50.190 314.870 ;
        RECT -60.705 314.525 -50.190 314.740 ;
        RECT -50.615 314.410 -50.190 314.525 ;
        RECT -61.220 313.535 -60.860 313.655 ;
        RECT -61.220 313.185 -53.825 313.535 ;
        RECT -61.220 313.130 -60.860 313.185 ;
        RECT -61.950 312.175 -60.515 312.215 ;
        RECT -61.950 312.005 -57.545 312.175 ;
        RECT -61.950 312.000 -60.515 312.005 ;
        RECT -61.950 311.790 -61.735 312.000 ;
        RECT -54.175 311.845 -53.825 313.185 ;
        RECT -62.150 311.760 -61.735 311.790 ;
        RECT -63.645 311.590 -61.735 311.760 ;
        RECT -62.150 311.570 -61.735 311.590 ;
        RECT -61.935 311.330 -61.735 311.570 ;
        RECT -61.285 311.140 -61.010 311.830 ;
        RECT -55.035 311.675 -53.825 311.845 ;
        RECT -53.880 311.185 -53.340 311.355 ;
        RECT -61.835 310.925 -60.755 311.140 ;
        RECT -57.595 311.115 -57.205 311.145 ;
        RECT -60.585 310.945 -57.205 311.115 ;
        RECT -57.595 310.935 -57.205 310.945 ;
        RECT -61.835 309.595 -61.635 310.925 ;
        RECT -60.950 310.645 -60.755 310.925 ;
        RECT -60.950 310.625 -60.485 310.645 ;
        RECT -61.395 309.715 -61.120 310.490 ;
        RECT -60.950 310.455 -57.545 310.625 ;
        RECT -60.950 310.435 -60.485 310.455 ;
        RECT -60.940 310.135 -60.495 310.160 ;
        RECT -57.375 310.155 -57.205 310.935 ;
        RECT -55.035 310.695 -54.495 310.865 ;
        RECT -53.880 310.205 -53.340 310.375 ;
        RECT -57.585 310.135 -57.205 310.155 ;
        RECT -60.940 309.965 -57.205 310.135 ;
        RECT -60.940 309.950 -60.495 309.965 ;
        RECT -62.185 309.570 -61.635 309.595 ;
        RECT -63.645 309.400 -61.635 309.570 ;
        RECT -62.185 309.370 -61.635 309.400 ;
        RECT -61.935 308.365 -61.660 309.140 ;
        RECT -61.875 308.180 -61.705 308.365 ;
        RECT -61.350 308.040 -61.170 309.715 ;
        RECT -60.940 309.100 -60.760 309.950 ;
        RECT -57.585 309.945 -57.205 309.965 ;
        RECT -55.035 309.715 -54.495 309.885 ;
        RECT -54.325 309.125 -54.025 309.490 ;
        RECT -60.940 309.080 -60.465 309.100 ;
        RECT -60.940 308.910 -57.545 309.080 ;
        RECT -60.940 308.890 -60.465 308.910 ;
        RECT -54.260 308.820 -54.055 309.125 ;
        RECT -54.260 308.765 -53.160 308.820 ;
        RECT -54.260 308.625 -53.120 308.765 ;
        RECT -54.120 308.515 -53.120 308.625 ;
        RECT -59.195 308.040 -58.845 308.070 ;
        RECT -61.360 307.690 -58.845 308.040 ;
        RECT -53.310 307.820 -53.120 308.515 ;
        RECT -52.885 308.080 -52.530 308.450 ;
        RECT -52.345 308.140 -50.805 308.310 ;
        RECT -59.195 306.850 -58.845 307.690 ;
        RECT -55.030 307.650 -53.120 307.820 ;
        RECT -59.195 306.680 -57.985 306.850 ;
        RECT -53.310 306.840 -53.120 307.650 ;
        RECT -55.030 306.670 -53.120 306.840 ;
        RECT -59.680 306.190 -59.140 306.360 ;
        RECT -58.525 305.700 -57.985 305.870 ;
        RECT -53.275 305.755 -53.005 306.430 ;
        RECT -52.755 306.375 -52.560 308.080 ;
        RECT -52.345 307.650 -50.805 307.820 ;
        RECT -52.345 307.160 -50.805 307.330 ;
        RECT -52.755 306.025 -52.555 306.375 ;
        RECT -52.345 306.180 -50.805 306.350 ;
        RECT -52.765 306.020 -52.555 306.025 ;
        RECT -53.245 305.655 -53.045 305.755 ;
        RECT -59.680 305.210 -59.140 305.380 ;
        RECT -58.525 304.720 -57.985 304.890 ;
        RECT -53.235 304.620 -53.055 305.655 ;
        RECT -58.995 304.130 -58.695 304.495 ;
        RECT -58.965 303.825 -58.760 304.130 ;
        RECT -59.860 303.770 -58.760 303.825 ;
        RECT -59.900 303.630 -58.760 303.770 ;
        RECT -54.385 303.765 -53.345 303.935 ;
        RECT -59.900 303.520 -58.900 303.630 ;
        RECT -62.215 303.145 -60.675 303.315 ;
        RECT -60.490 303.085 -60.135 303.455 ;
        RECT -62.215 302.655 -60.675 302.825 ;
        RECT -62.215 302.165 -60.675 302.335 ;
        RECT -60.460 301.380 -60.265 303.085 ;
        RECT -59.900 302.825 -59.710 303.520 ;
        RECT -52.765 303.445 -52.565 306.020 ;
        RECT -52.765 303.280 -51.695 303.445 ;
        RECT -52.735 303.275 -51.695 303.280 ;
        RECT -59.900 302.655 -57.990 302.825 ;
        RECT -54.385 302.785 -53.345 302.955 ;
        RECT -59.900 301.845 -59.710 302.655 ;
        RECT -52.735 302.295 -51.695 302.465 ;
        RECT -59.900 301.675 -57.990 301.845 ;
        RECT -54.385 301.805 -53.345 301.975 ;
        RECT -62.215 301.185 -60.675 301.355 ;
        RECT -60.465 301.030 -60.265 301.380 ;
        RECT -53.175 301.215 -52.875 301.580 ;
        RECT -60.465 301.025 -60.255 301.030 ;
        RECT -60.455 299.895 -60.255 301.025 ;
        RECT -53.110 300.995 -52.905 301.215 ;
        RECT -53.195 300.700 -52.445 300.995 ;
        RECT -53.195 300.370 -50.120 300.700 ;
        RECT -49.210 300.370 -48.830 316.160 ;
        RECT -43.090 315.990 -42.920 317.725 ;
        RECT -44.685 315.775 -42.920 315.990 ;
        RECT -44.685 312.255 -44.470 315.775 ;
        RECT -43.955 313.575 -43.595 313.695 ;
        RECT -43.955 313.225 -36.560 313.575 ;
        RECT -43.955 313.170 -43.595 313.225 ;
        RECT -44.685 312.215 -43.250 312.255 ;
        RECT -44.685 312.045 -40.280 312.215 ;
        RECT -44.685 312.040 -43.250 312.045 ;
        RECT -44.685 311.830 -44.470 312.040 ;
        RECT -36.910 311.885 -36.560 313.225 ;
        RECT -44.885 311.800 -44.470 311.830 ;
        RECT -46.380 311.630 -44.470 311.800 ;
        RECT -44.885 311.610 -44.470 311.630 ;
        RECT -44.670 311.370 -44.470 311.610 ;
        RECT -44.020 311.180 -43.745 311.870 ;
        RECT -37.770 311.715 -36.560 311.885 ;
        RECT -36.615 311.225 -36.075 311.395 ;
        RECT -44.570 310.965 -43.490 311.180 ;
        RECT -40.330 311.155 -39.940 311.185 ;
        RECT -43.320 310.985 -39.940 311.155 ;
        RECT -40.330 310.975 -39.940 310.985 ;
        RECT -44.570 309.635 -44.370 310.965 ;
        RECT -43.685 310.685 -43.490 310.965 ;
        RECT -43.685 310.665 -43.220 310.685 ;
        RECT -44.130 309.755 -43.855 310.530 ;
        RECT -43.685 310.495 -40.280 310.665 ;
        RECT -43.685 310.475 -43.220 310.495 ;
        RECT -43.675 310.175 -43.230 310.200 ;
        RECT -40.110 310.195 -39.940 310.975 ;
        RECT -37.770 310.735 -37.230 310.905 ;
        RECT -36.615 310.245 -36.075 310.415 ;
        RECT -40.320 310.175 -39.940 310.195 ;
        RECT -43.675 310.005 -39.940 310.175 ;
        RECT -43.675 309.990 -43.230 310.005 ;
        RECT -44.920 309.610 -44.370 309.635 ;
        RECT -46.380 309.440 -44.370 309.610 ;
        RECT -44.920 309.410 -44.370 309.440 ;
        RECT -44.670 308.405 -44.395 309.180 ;
        RECT -44.610 308.220 -44.440 308.405 ;
        RECT -44.085 308.080 -43.905 309.755 ;
        RECT -43.675 309.140 -43.495 309.990 ;
        RECT -40.320 309.985 -39.940 310.005 ;
        RECT -37.770 309.755 -37.230 309.925 ;
        RECT -37.060 309.165 -36.760 309.530 ;
        RECT -43.675 309.120 -43.200 309.140 ;
        RECT -43.675 308.950 -40.280 309.120 ;
        RECT -43.675 308.930 -43.200 308.950 ;
        RECT -36.995 308.860 -36.790 309.165 ;
        RECT -36.995 308.805 -35.895 308.860 ;
        RECT -36.995 308.665 -35.855 308.805 ;
        RECT -36.855 308.555 -35.855 308.665 ;
        RECT -41.930 308.080 -41.580 308.110 ;
        RECT -44.095 307.730 -41.580 308.080 ;
        RECT -36.045 307.860 -35.855 308.555 ;
        RECT -35.620 308.120 -35.265 308.490 ;
        RECT -35.080 308.180 -33.540 308.350 ;
        RECT -41.930 306.890 -41.580 307.730 ;
        RECT -37.765 307.690 -35.855 307.860 ;
        RECT -41.930 306.720 -40.720 306.890 ;
        RECT -36.045 306.880 -35.855 307.690 ;
        RECT -37.765 306.710 -35.855 306.880 ;
        RECT -35.490 306.415 -35.295 308.120 ;
        RECT -35.080 307.690 -33.540 307.860 ;
        RECT -35.080 307.200 -33.540 307.370 ;
        RECT -42.415 306.230 -41.875 306.400 ;
        RECT -35.490 306.065 -35.290 306.415 ;
        RECT -35.080 306.220 -33.540 306.390 ;
        RECT -35.500 306.060 -35.290 306.065 ;
        RECT -41.260 305.740 -40.720 305.910 ;
        RECT -42.415 305.250 -41.875 305.420 ;
        RECT -41.260 304.760 -40.720 304.930 ;
        RECT -41.730 304.170 -41.430 304.535 ;
        RECT -41.700 303.865 -41.495 304.170 ;
        RECT -42.595 303.810 -41.495 303.865 ;
        RECT -42.635 303.670 -41.495 303.810 ;
        RECT -37.120 303.805 -36.080 303.975 ;
        RECT -42.635 303.560 -41.635 303.670 ;
        RECT -44.950 303.185 -43.410 303.355 ;
        RECT -43.225 303.125 -42.870 303.495 ;
        RECT -44.950 302.695 -43.410 302.865 ;
        RECT -44.950 302.205 -43.410 302.375 ;
        RECT -43.195 301.420 -43.000 303.125 ;
        RECT -42.635 302.865 -42.445 303.560 ;
        RECT -35.500 303.485 -35.300 306.060 ;
        RECT -35.500 303.320 -34.430 303.485 ;
        RECT -35.470 303.315 -34.430 303.320 ;
        RECT -42.635 302.695 -40.725 302.865 ;
        RECT -37.120 302.825 -36.080 302.995 ;
        RECT -42.635 301.885 -42.445 302.695 ;
        RECT -35.470 302.335 -34.430 302.505 ;
        RECT -42.635 301.715 -40.725 301.885 ;
        RECT -37.120 301.845 -36.080 302.015 ;
        RECT -44.950 301.225 -43.410 301.395 ;
        RECT -43.200 301.070 -43.000 301.420 ;
        RECT -35.910 301.255 -35.610 301.620 ;
        RECT -43.200 301.065 -42.990 301.070 ;
        RECT -43.190 300.370 -42.990 301.065 ;
        RECT -35.845 301.035 -35.640 301.255 ;
        RECT -35.930 300.385 -35.180 301.035 ;
        RECT -53.195 300.345 -42.990 300.370 ;
        RECT -52.990 300.320 -42.990 300.345 ;
        RECT -50.500 299.990 -42.990 300.320 ;
        RECT -68.880 296.740 -68.040 296.835 ;
        RECT -49.280 296.740 -48.550 299.990 ;
        RECT -43.190 299.935 -42.990 299.990 ;
        RECT -68.880 296.455 -48.550 296.740 ;
        RECT -68.885 296.010 -48.550 296.455 ;
        RECT -68.885 286.680 -68.030 296.010 ;
        RECT -52.415 289.925 -52.245 289.940 ;
        RECT -52.495 289.335 -52.205 289.925 ;
        RECT -42.120 289.905 -41.435 289.910 ;
        RECT -44.095 289.900 -39.355 289.905 ;
        RECT -44.105 289.870 -39.355 289.900 ;
        RECT -44.105 289.665 -39.205 289.870 ;
        RECT -44.105 289.490 -43.910 289.665 ;
        RECT -42.120 289.610 -41.435 289.665 ;
        RECT -44.150 289.340 -43.800 289.490 ;
        RECT -52.415 289.100 -52.245 289.335 ;
        RECT -44.515 289.310 -43.495 289.340 ;
        RECT -45.475 289.140 -43.035 289.310 ;
        RECT -44.515 289.110 -43.495 289.140 ;
        RECT -56.385 288.930 -48.420 289.100 ;
        RECT -52.530 288.055 -52.260 288.725 ;
        RECT -44.190 288.360 -43.960 289.110 ;
        RECT -39.575 289.030 -39.205 289.665 ;
        RECT -39.825 288.820 -37.865 288.850 ;
        RECT -40.285 288.650 -37.845 288.820 ;
        RECT -39.825 288.620 -37.865 288.650 ;
        RECT -44.515 288.330 -43.495 288.360 ;
        RECT -45.475 288.160 -43.035 288.330 ;
        RECT -44.515 288.130 -43.495 288.160 ;
        RECT -52.490 287.100 -52.295 288.055 ;
        RECT -44.190 287.380 -43.960 288.130 ;
        RECT -45.455 287.350 -43.495 287.380 ;
        RECT -45.475 287.180 -43.035 287.350 ;
        RECT -45.455 287.150 -43.495 287.180 ;
        RECT -56.385 286.930 -48.420 287.100 ;
        RECT -52.545 286.130 -52.275 286.695 ;
        RECT -44.115 286.130 -43.745 286.970 ;
        RECT -42.205 286.225 -42.010 288.255 ;
        RECT -39.360 287.870 -39.130 288.620 ;
        RECT -39.825 287.840 -38.805 287.870 ;
        RECT -40.285 287.670 -37.845 287.840 ;
        RECT -39.825 287.640 -38.805 287.670 ;
        RECT -39.360 286.890 -39.130 287.640 ;
        RECT -39.825 286.860 -38.805 286.890 ;
        RECT -40.285 286.690 -37.845 286.860 ;
        RECT -39.825 286.660 -38.805 286.690 ;
        RECT -39.520 286.455 -39.170 286.660 ;
        RECT -39.520 286.225 -38.275 286.455 ;
        RECT -52.545 285.780 -51.340 286.130 ;
        RECT -52.555 284.855 -52.265 285.445 ;
        RECT -44.085 285.145 -43.820 286.130 ;
        RECT -42.270 285.565 -41.970 286.225 ;
        RECT -40.295 285.860 -39.265 286.045 ;
        RECT -40.295 285.745 -39.260 285.860 ;
        RECT -39.575 285.685 -39.260 285.745 ;
        RECT -38.520 285.740 -38.275 286.225 ;
        RECT -44.900 285.140 -43.470 285.145 ;
        RECT -44.900 285.120 -43.255 285.140 ;
        RECT -45.400 284.950 -42.785 285.120 ;
        RECT -44.900 284.935 -43.255 284.950 ;
        RECT -52.495 284.100 -52.325 284.855 ;
        RECT -45.740 284.630 -45.315 284.655 ;
        RECT -45.740 284.460 -44.860 284.630 ;
        RECT -45.740 284.445 -45.315 284.460 ;
        RECT -56.385 283.930 -48.420 284.100 ;
        RECT -52.520 283.090 -52.250 283.760 ;
        RECT -45.740 283.675 -45.570 284.445 ;
        RECT -44.680 284.270 -43.505 284.935 ;
        RECT -42.845 284.630 -42.385 284.660 ;
        RECT -43.325 284.460 -42.385 284.630 ;
        RECT -42.845 284.440 -42.385 284.460 ;
        RECT -44.680 284.145 -44.510 284.270 ;
        RECT -44.950 284.140 -44.510 284.145 ;
        RECT -45.400 283.970 -44.510 284.140 ;
        RECT -44.950 283.965 -44.510 283.970 ;
        RECT -45.740 283.650 -45.290 283.675 ;
        RECT -45.740 283.480 -44.860 283.650 ;
        RECT -45.740 283.465 -45.290 283.480 ;
        RECT -52.485 282.100 -52.290 283.090 ;
        RECT -45.740 282.705 -45.570 283.465 ;
        RECT -44.680 283.175 -44.510 283.965 ;
        RECT -44.950 283.160 -44.510 283.175 ;
        RECT -45.400 282.995 -44.510 283.160 ;
        RECT -45.400 282.990 -44.860 282.995 ;
        RECT -45.740 282.670 -45.295 282.705 ;
        RECT -45.740 282.500 -44.860 282.670 ;
        RECT -45.740 282.495 -45.295 282.500 ;
        RECT -56.385 281.930 -48.420 282.100 ;
        RECT -45.740 281.695 -45.570 282.495 ;
        RECT -44.680 282.185 -44.510 282.995 ;
        RECT -43.675 284.155 -43.505 284.270 ;
        RECT -43.675 284.140 -43.260 284.155 ;
        RECT -43.675 283.970 -42.785 284.140 ;
        RECT -43.675 283.950 -43.260 283.970 ;
        RECT -43.675 283.185 -43.505 283.950 ;
        RECT -42.555 283.675 -42.385 284.440 ;
        RECT -42.900 283.650 -42.385 283.675 ;
        RECT -43.325 283.480 -42.385 283.650 ;
        RECT -42.900 283.455 -42.385 283.480 ;
        RECT -43.675 283.160 -43.260 283.185 ;
        RECT -43.675 282.990 -42.785 283.160 ;
        RECT -43.675 282.980 -43.260 282.990 ;
        RECT -44.940 282.180 -44.510 282.185 ;
        RECT -45.400 282.010 -44.510 282.180 ;
        RECT -44.940 282.005 -44.510 282.010 ;
        RECT -44.240 281.725 -43.870 282.350 ;
        RECT -43.675 282.195 -43.505 282.980 ;
        RECT -42.555 282.695 -42.385 283.455 ;
        RECT -42.900 282.670 -42.385 282.695 ;
        RECT -43.325 282.500 -42.385 282.670 ;
        RECT -42.900 282.475 -42.385 282.500 ;
        RECT -43.675 282.180 -43.300 282.195 ;
        RECT -43.675 282.010 -42.785 282.180 ;
        RECT -43.675 281.990 -43.300 282.010 ;
        RECT -52.510 281.175 -52.240 281.695 ;
        RECT -45.740 281.690 -45.345 281.695 ;
        RECT -44.975 281.690 -43.195 281.725 ;
        RECT -42.555 281.715 -42.385 282.475 ;
        RECT -42.845 281.690 -42.385 281.715 ;
        RECT -45.740 281.520 -42.385 281.690 ;
        RECT -45.740 281.515 -45.345 281.520 ;
        RECT -44.975 281.490 -43.195 281.520 ;
        RECT -42.845 281.495 -42.385 281.520 ;
        RECT -45.110 281.265 -44.270 281.270 ;
        RECT -52.510 280.825 -51.335 281.175 ;
        RECT -45.110 280.900 -43.800 281.265 ;
        RECT -44.150 280.625 -43.800 280.900 ;
        RECT -44.515 280.595 -43.495 280.625 ;
        RECT -45.475 280.425 -43.035 280.595 ;
        RECT -44.515 280.395 -43.495 280.425 ;
        RECT -52.420 279.470 -52.130 280.060 ;
        RECT -44.190 279.645 -43.960 280.395 ;
        RECT -44.515 279.615 -43.495 279.645 ;
        RECT -52.360 279.100 -52.190 279.470 ;
        RECT -45.475 279.445 -43.035 279.615 ;
        RECT -44.515 279.415 -43.495 279.445 ;
        RECT -56.385 278.930 -48.420 279.100 ;
        RECT -52.445 278.090 -52.175 278.760 ;
        RECT -44.190 278.665 -43.960 279.415 ;
        RECT -45.455 278.635 -43.495 278.665 ;
        RECT -45.475 278.465 -43.035 278.635 ;
        RECT -45.455 278.435 -43.495 278.465 ;
        RECT -52.410 277.100 -52.240 278.090 ;
        RECT -45.365 277.360 -44.545 277.645 ;
        RECT -56.385 276.930 -48.420 277.100 ;
        RECT -52.520 275.955 -52.250 276.750 ;
        RECT -44.975 276.565 -44.750 277.360 ;
        RECT -44.975 276.540 -43.855 276.565 ;
        RECT -44.975 276.340 -43.280 276.540 ;
        RECT -44.080 276.240 -43.280 276.340 ;
        RECT -44.080 275.990 -43.855 276.240 ;
        RECT -55.415 275.605 -48.580 275.955 ;
        RECT -44.150 275.840 -43.800 275.990 ;
        RECT -44.515 275.810 -43.495 275.840 ;
        RECT -45.475 275.640 -43.035 275.810 ;
        RECT -44.515 275.610 -43.495 275.640 ;
        RECT -55.415 274.690 -55.065 275.605 ;
        RECT -44.190 274.860 -43.960 275.610 ;
        RECT -44.515 274.830 -43.495 274.860 ;
        RECT -55.780 274.660 -54.760 274.690 ;
        RECT -56.740 274.490 -54.300 274.660 ;
        RECT -55.780 274.460 -54.760 274.490 ;
        RECT -51.150 274.480 -50.480 274.780 ;
        RECT -45.475 274.660 -43.035 274.830 ;
        RECT -44.515 274.630 -43.495 274.660 ;
        RECT -55.455 273.710 -55.225 274.460 ;
        RECT -51.085 274.000 -50.780 274.480 ;
        RECT -52.505 273.930 -50.420 274.000 ;
        RECT -52.505 273.830 -48.195 273.930 ;
        RECT -44.190 273.880 -43.960 274.630 ;
        RECT -45.455 273.850 -43.495 273.880 ;
        RECT -50.605 273.760 -48.195 273.830 ;
        RECT -55.780 273.680 -54.760 273.710 ;
        RECT -56.740 273.510 -54.300 273.680 ;
        RECT -55.780 273.480 -54.760 273.510 ;
        RECT -55.455 272.730 -55.225 273.480 ;
        RECT -52.780 273.340 -51.465 273.510 ;
        RECT -52.780 272.950 -52.605 273.340 ;
        RECT -51.210 272.955 -50.940 273.630 ;
        RECT -52.780 272.780 -51.465 272.950 ;
        RECT -56.720 272.700 -54.760 272.730 ;
        RECT -56.740 272.530 -54.300 272.700 ;
        RECT -56.720 272.500 -54.760 272.530 ;
        RECT -51.165 272.485 -50.970 272.955 ;
        RECT -50.605 272.950 -50.415 273.760 ;
        RECT -45.475 273.680 -43.035 273.850 ;
        RECT -45.455 273.650 -43.495 273.680 ;
        RECT -50.605 272.780 -48.195 272.950 ;
        RECT -44.115 272.630 -43.745 273.470 ;
        RECT -55.380 271.480 -55.010 272.320 ;
        RECT -51.170 272.215 -50.970 272.485 ;
        RECT -51.235 272.210 -50.945 272.215 ;
        RECT -51.240 271.415 -50.940 272.210 ;
        RECT -50.720 271.865 -50.450 272.540 ;
        RECT -50.680 271.765 -50.480 271.865 ;
        RECT -50.665 270.310 -50.485 271.765 ;
        RECT -44.070 271.645 -43.785 272.630 ;
        RECT -44.900 271.640 -43.470 271.645 ;
        RECT -44.900 271.635 -43.255 271.640 ;
        RECT -44.900 271.620 -42.645 271.635 ;
        RECT -45.400 271.450 -42.645 271.620 ;
        RECT -44.900 271.435 -42.645 271.450 ;
        RECT -45.740 271.130 -45.315 271.155 ;
        RECT -48.820 270.890 -48.160 270.965 ;
        RECT -47.245 270.890 -46.585 270.980 ;
        RECT -54.460 269.615 -54.160 270.270 ;
        RECT -50.735 269.650 -50.435 270.310 ;
        RECT -48.820 270.215 -46.585 270.890 ;
        RECT -48.820 270.165 -48.160 270.215 ;
        RECT -47.245 270.180 -46.585 270.215 ;
        RECT -45.740 270.960 -44.860 271.130 ;
        RECT -45.740 270.945 -45.315 270.960 ;
        RECT -45.740 270.175 -45.570 270.945 ;
        RECT -44.680 270.770 -43.505 271.435 ;
        RECT -43.305 271.405 -42.645 271.435 ;
        RECT -42.845 271.130 -42.385 271.160 ;
        RECT -43.325 270.960 -42.385 271.130 ;
        RECT -42.845 270.940 -42.385 270.960 ;
        RECT -44.680 270.645 -44.510 270.770 ;
        RECT -44.950 270.640 -44.510 270.645 ;
        RECT -45.400 270.470 -44.510 270.640 ;
        RECT -44.950 270.465 -44.510 270.470 ;
        RECT -45.740 270.150 -45.290 270.175 ;
        RECT -45.740 269.980 -44.860 270.150 ;
        RECT -45.740 269.965 -45.290 269.980 ;
        RECT -54.340 269.055 -54.160 269.615 ;
        RECT -45.740 269.205 -45.570 269.965 ;
        RECT -44.680 269.675 -44.510 270.465 ;
        RECT -44.950 269.660 -44.510 269.675 ;
        RECT -45.400 269.495 -44.510 269.660 ;
        RECT -45.400 269.490 -44.860 269.495 ;
        RECT -45.740 269.170 -45.295 269.205 ;
        RECT -56.775 268.885 -52.195 269.055 ;
        RECT -45.740 269.000 -44.860 269.170 ;
        RECT -45.740 268.995 -45.295 269.000 ;
        RECT -54.730 268.035 -54.460 268.710 ;
        RECT -45.740 268.195 -45.570 268.995 ;
        RECT -44.680 268.685 -44.510 269.495 ;
        RECT -43.675 270.655 -43.505 270.770 ;
        RECT -43.675 270.640 -43.260 270.655 ;
        RECT -43.675 270.470 -42.785 270.640 ;
        RECT -43.675 270.450 -43.260 270.470 ;
        RECT -43.675 269.685 -43.505 270.450 ;
        RECT -42.555 270.175 -42.385 270.940 ;
        RECT -42.900 270.150 -42.385 270.175 ;
        RECT -43.325 269.980 -42.385 270.150 ;
        RECT -42.900 269.955 -42.385 269.980 ;
        RECT -43.675 269.660 -43.260 269.685 ;
        RECT -43.675 269.490 -42.785 269.660 ;
        RECT -43.675 269.480 -43.260 269.490 ;
        RECT -44.940 268.680 -44.510 268.685 ;
        RECT -45.400 268.510 -44.510 268.680 ;
        RECT -44.940 268.505 -44.510 268.510 ;
        RECT -44.240 268.225 -43.870 268.850 ;
        RECT -43.675 268.695 -43.505 269.480 ;
        RECT -42.555 269.195 -42.385 269.955 ;
        RECT -42.900 269.170 -42.385 269.195 ;
        RECT -43.325 269.000 -42.385 269.170 ;
        RECT -42.900 268.975 -42.385 269.000 ;
        RECT -43.675 268.680 -43.300 268.695 ;
        RECT -43.675 268.510 -42.785 268.680 ;
        RECT -43.675 268.490 -43.300 268.510 ;
        RECT -45.740 268.190 -45.345 268.195 ;
        RECT -44.975 268.190 -43.195 268.225 ;
        RECT -42.555 268.215 -42.385 268.975 ;
        RECT -42.845 268.190 -42.385 268.215 ;
        RECT -54.680 266.010 -54.495 268.035 ;
        RECT -45.740 268.020 -42.385 268.190 ;
        RECT -45.740 268.015 -45.345 268.020 ;
        RECT -44.975 267.990 -43.195 268.020 ;
        RECT -42.845 267.995 -42.385 268.020 ;
        RECT -45.110 267.765 -44.270 267.770 ;
        RECT -45.110 267.400 -43.800 267.765 ;
        RECT -44.150 267.125 -43.800 267.400 ;
        RECT -44.515 267.095 -43.495 267.125 ;
        RECT -54.225 266.820 -52.195 266.990 ;
        RECT -45.475 266.925 -43.035 267.095 ;
        RECT -44.515 266.895 -43.495 266.925 ;
        RECT -54.225 266.010 -54.055 266.820 ;
        RECT -53.735 266.330 -51.535 266.500 ;
        RECT -55.555 265.840 -52.195 266.010 ;
        RECT -55.555 265.825 -54.055 265.840 ;
        RECT -55.555 265.365 -55.370 265.825 ;
        RECT -56.775 265.195 -55.370 265.365 ;
        RECT -55.555 264.385 -55.370 265.195 ;
        RECT -54.740 264.980 -54.470 265.655 ;
        RECT -51.705 265.450 -51.535 266.330 ;
        RECT -44.190 266.145 -43.960 266.895 ;
        RECT -44.515 266.115 -43.495 266.145 ;
        RECT -45.475 265.945 -43.035 266.115 ;
        RECT -44.515 265.915 -43.495 265.945 ;
        RECT -52.250 265.445 -51.535 265.450 ;
        RECT -53.735 265.275 -51.535 265.445 ;
        RECT -56.775 264.215 -55.370 264.385 ;
        RECT -55.555 263.405 -55.370 264.215 ;
        RECT -55.130 264.040 -54.860 264.715 ;
        RECT -56.775 263.235 -55.370 263.405 ;
        RECT -55.540 262.360 -55.270 263.035 ;
        RECT -55.500 262.265 -55.315 262.360 ;
        RECT -55.490 262.000 -55.315 262.265 ;
        RECT -55.975 261.700 -55.315 262.000 ;
        RECT -55.085 261.425 -54.895 264.040 ;
        RECT -54.675 262.470 -54.505 264.980 ;
        RECT -54.225 264.955 -53.735 264.960 ;
        RECT -54.225 264.785 -52.195 264.955 ;
        RECT -54.225 263.895 -54.050 264.785 ;
        RECT -51.720 264.470 -51.535 265.275 ;
        RECT -44.190 265.165 -43.960 265.915 ;
        RECT -45.455 265.135 -43.495 265.165 ;
        RECT -45.475 264.965 -43.035 265.135 ;
        RECT -45.455 264.935 -43.495 264.965 ;
        RECT -52.240 264.465 -51.535 264.470 ;
        RECT -53.735 264.295 -51.535 264.465 ;
        RECT -54.225 263.725 -52.200 263.895 ;
        RECT -45.365 263.860 -44.545 264.145 ;
        RECT -44.115 263.915 -43.745 264.755 ;
        RECT -44.060 263.740 -43.770 263.915 ;
        RECT -54.225 262.915 -54.055 263.725 ;
        RECT -44.040 263.455 -43.830 263.740 ;
        RECT -42.205 263.610 -42.010 285.565 ;
        RECT -39.575 284.845 -39.205 285.685 ;
        RECT -38.775 285.455 -37.955 285.740 ;
        RECT -39.825 284.635 -37.865 284.665 ;
        RECT -40.285 284.465 -37.845 284.635 ;
        RECT -39.825 284.435 -37.865 284.465 ;
        RECT -39.360 283.685 -39.130 284.435 ;
        RECT -39.825 283.655 -38.805 283.685 ;
        RECT -40.285 283.485 -37.845 283.655 ;
        RECT -39.825 283.455 -38.805 283.485 ;
        RECT -39.360 282.705 -39.130 283.455 ;
        RECT -39.825 282.675 -38.805 282.705 ;
        RECT -40.285 282.505 -37.845 282.675 ;
        RECT -39.825 282.475 -38.805 282.505 ;
        RECT -39.520 282.200 -39.170 282.475 ;
        RECT -39.520 281.835 -38.210 282.200 ;
        RECT -39.050 281.830 -38.210 281.835 ;
        RECT -40.935 281.580 -40.475 281.605 ;
        RECT -40.125 281.580 -38.345 281.610 ;
        RECT -37.975 281.580 -37.580 281.585 ;
        RECT -40.935 281.410 -37.580 281.580 ;
        RECT -40.935 281.385 -40.475 281.410 ;
        RECT -40.935 280.625 -40.765 281.385 ;
        RECT -40.125 281.375 -38.345 281.410 ;
        RECT -37.975 281.405 -37.580 281.410 ;
        RECT -40.020 281.090 -39.645 281.110 ;
        RECT -40.535 280.920 -39.645 281.090 ;
        RECT -40.020 280.905 -39.645 280.920 ;
        RECT -40.935 280.600 -40.420 280.625 ;
        RECT -40.935 280.430 -39.995 280.600 ;
        RECT -40.935 280.405 -40.420 280.430 ;
        RECT -40.935 279.645 -40.765 280.405 ;
        RECT -39.815 280.120 -39.645 280.905 ;
        RECT -39.450 280.750 -39.080 281.375 ;
        RECT -38.810 281.090 -38.380 281.095 ;
        RECT -38.810 280.920 -37.920 281.090 ;
        RECT -38.810 280.915 -38.380 280.920 ;
        RECT -40.060 280.110 -39.645 280.120 ;
        RECT -40.535 279.940 -39.645 280.110 ;
        RECT -40.060 279.915 -39.645 279.940 ;
        RECT -40.935 279.620 -40.420 279.645 ;
        RECT -40.935 279.450 -39.995 279.620 ;
        RECT -40.935 279.425 -40.420 279.450 ;
        RECT -40.935 278.660 -40.765 279.425 ;
        RECT -39.815 279.150 -39.645 279.915 ;
        RECT -40.060 279.130 -39.645 279.150 ;
        RECT -40.535 278.960 -39.645 279.130 ;
        RECT -40.060 278.945 -39.645 278.960 ;
        RECT -39.815 278.830 -39.645 278.945 ;
        RECT -38.810 280.105 -38.640 280.915 ;
        RECT -37.750 280.605 -37.580 281.405 ;
        RECT -38.025 280.600 -37.580 280.605 ;
        RECT -38.460 280.430 -37.580 280.600 ;
        RECT -38.025 280.395 -37.580 280.430 ;
        RECT -38.460 280.105 -37.920 280.110 ;
        RECT -38.810 279.940 -37.920 280.105 ;
        RECT -38.810 279.925 -38.370 279.940 ;
        RECT -38.810 279.135 -38.640 279.925 ;
        RECT -37.750 279.635 -37.580 280.395 ;
        RECT -38.030 279.620 -37.580 279.635 ;
        RECT -38.460 279.450 -37.580 279.620 ;
        RECT -38.030 279.425 -37.580 279.450 ;
        RECT -38.810 279.130 -38.370 279.135 ;
        RECT -38.810 278.960 -37.920 279.130 ;
        RECT -38.810 278.955 -38.370 278.960 ;
        RECT -38.810 278.830 -38.640 278.955 ;
        RECT -40.935 278.640 -40.475 278.660 ;
        RECT -40.935 278.470 -39.995 278.640 ;
        RECT -40.935 278.440 -40.475 278.470 ;
        RECT -39.815 278.165 -38.640 278.830 ;
        RECT -37.750 278.655 -37.580 279.425 ;
        RECT -38.005 278.640 -37.580 278.655 ;
        RECT -38.460 278.470 -37.580 278.640 ;
        RECT -38.005 278.445 -37.580 278.470 ;
        RECT -40.065 278.150 -38.420 278.165 ;
        RECT -40.535 277.980 -37.920 278.150 ;
        RECT -40.065 277.960 -38.420 277.980 ;
        RECT -39.850 277.955 -38.420 277.960 ;
        RECT -39.645 277.500 -39.345 277.955 ;
        RECT -39.540 276.370 -39.240 276.480 ;
        RECT -39.575 275.530 -39.205 276.370 ;
        RECT -39.825 275.320 -37.865 275.350 ;
        RECT -40.285 275.150 -37.845 275.320 ;
        RECT -39.825 275.120 -37.865 275.150 ;
        RECT -39.360 274.370 -39.130 275.120 ;
        RECT -39.825 274.340 -38.805 274.370 ;
        RECT -40.285 274.170 -37.845 274.340 ;
        RECT -39.825 274.140 -38.805 274.170 ;
        RECT -39.360 273.390 -39.130 274.140 ;
        RECT -39.825 273.360 -38.805 273.390 ;
        RECT -40.285 273.190 -37.845 273.360 ;
        RECT -39.825 273.160 -38.805 273.190 ;
        RECT -39.520 272.980 -39.170 273.160 ;
        RECT -39.520 272.670 -38.215 272.980 ;
        RECT -38.525 272.240 -38.215 272.670 ;
        RECT -38.775 271.955 -37.955 272.240 ;
        RECT -39.825 271.135 -37.865 271.165 ;
        RECT -40.285 270.965 -37.845 271.135 ;
        RECT -39.825 270.935 -37.865 270.965 ;
        RECT -39.360 270.185 -39.130 270.935 ;
        RECT -39.825 270.155 -38.805 270.185 ;
        RECT -40.285 269.985 -37.845 270.155 ;
        RECT -39.825 269.955 -38.805 269.985 ;
        RECT -39.360 269.205 -39.130 269.955 ;
        RECT -39.825 269.175 -38.805 269.205 ;
        RECT -40.285 269.005 -37.845 269.175 ;
        RECT -39.825 268.975 -38.805 269.005 ;
        RECT -39.520 268.700 -39.170 268.975 ;
        RECT -39.520 268.335 -38.210 268.700 ;
        RECT -39.050 268.330 -38.210 268.335 ;
        RECT -40.935 268.080 -40.475 268.105 ;
        RECT -40.125 268.080 -38.345 268.110 ;
        RECT -37.975 268.080 -37.580 268.085 ;
        RECT -40.935 267.910 -37.580 268.080 ;
        RECT -40.935 267.885 -40.475 267.910 ;
        RECT -40.935 267.125 -40.765 267.885 ;
        RECT -40.125 267.875 -38.345 267.910 ;
        RECT -37.975 267.905 -37.580 267.910 ;
        RECT -40.020 267.590 -39.645 267.610 ;
        RECT -40.535 267.420 -39.645 267.590 ;
        RECT -40.020 267.405 -39.645 267.420 ;
        RECT -40.935 267.100 -40.420 267.125 ;
        RECT -40.935 266.930 -39.995 267.100 ;
        RECT -40.935 266.905 -40.420 266.930 ;
        RECT -40.935 266.145 -40.765 266.905 ;
        RECT -39.815 266.620 -39.645 267.405 ;
        RECT -39.450 267.250 -39.080 267.875 ;
        RECT -38.810 267.590 -38.380 267.595 ;
        RECT -38.810 267.420 -37.920 267.590 ;
        RECT -38.810 267.415 -38.380 267.420 ;
        RECT -40.060 266.610 -39.645 266.620 ;
        RECT -40.535 266.440 -39.645 266.610 ;
        RECT -40.060 266.415 -39.645 266.440 ;
        RECT -40.935 266.120 -40.420 266.145 ;
        RECT -40.935 265.950 -39.995 266.120 ;
        RECT -40.935 265.925 -40.420 265.950 ;
        RECT -40.935 265.160 -40.765 265.925 ;
        RECT -39.815 265.650 -39.645 266.415 ;
        RECT -40.060 265.630 -39.645 265.650 ;
        RECT -40.535 265.460 -39.645 265.630 ;
        RECT -40.060 265.445 -39.645 265.460 ;
        RECT -39.815 265.330 -39.645 265.445 ;
        RECT -38.810 266.605 -38.640 267.415 ;
        RECT -37.750 267.105 -37.580 267.905 ;
        RECT -38.025 267.100 -37.580 267.105 ;
        RECT -38.460 266.930 -37.580 267.100 ;
        RECT -38.025 266.895 -37.580 266.930 ;
        RECT -38.460 266.605 -37.920 266.610 ;
        RECT -38.810 266.440 -37.920 266.605 ;
        RECT -38.810 266.425 -38.370 266.440 ;
        RECT -38.810 265.635 -38.640 266.425 ;
        RECT -37.750 266.135 -37.580 266.895 ;
        RECT -38.030 266.120 -37.580 266.135 ;
        RECT -38.460 265.950 -37.580 266.120 ;
        RECT -38.030 265.925 -37.580 265.950 ;
        RECT -38.810 265.630 -38.370 265.635 ;
        RECT -38.810 265.460 -37.920 265.630 ;
        RECT -38.810 265.455 -38.370 265.460 ;
        RECT -38.810 265.330 -38.640 265.455 ;
        RECT -40.935 265.140 -40.475 265.160 ;
        RECT -40.935 264.970 -39.995 265.140 ;
        RECT -40.935 264.940 -40.475 264.970 ;
        RECT -39.815 264.665 -38.640 265.330 ;
        RECT -37.750 265.155 -37.580 265.925 ;
        RECT -38.005 265.140 -37.580 265.155 ;
        RECT -38.460 264.970 -37.580 265.140 ;
        RECT -38.005 264.945 -37.580 264.970 ;
        RECT -40.065 264.650 -38.420 264.665 ;
        RECT -40.535 264.480 -37.920 264.650 ;
        RECT -40.065 264.460 -38.420 264.480 ;
        RECT -39.850 264.455 -38.420 264.460 ;
        RECT -39.655 264.080 -39.355 264.455 ;
        RECT -44.060 263.155 -43.400 263.455 ;
        RECT -54.225 262.745 -52.200 262.915 ;
        RECT -44.040 262.865 -43.830 263.155 ;
        RECT -42.260 262.950 -41.960 263.610 ;
        RECT -44.150 262.715 -43.800 262.865 ;
        RECT -44.515 262.685 -43.495 262.715 ;
        RECT -45.475 262.515 -43.035 262.685 ;
        RECT -44.515 262.485 -43.495 262.515 ;
        RECT -54.675 262.300 -53.345 262.470 ;
        RECT -54.675 262.275 -54.505 262.300 ;
        RECT -55.085 261.125 -54.065 261.425 ;
        RECT -53.570 260.925 -53.345 262.300 ;
        RECT -44.190 261.735 -43.960 262.485 ;
        RECT -44.515 261.705 -43.495 261.735 ;
        RECT -45.475 261.535 -43.035 261.705 ;
        RECT -44.515 261.505 -43.495 261.535 ;
        RECT -56.975 260.860 -56.465 260.895 ;
        RECT -54.795 260.860 -53.345 260.925 ;
        RECT -56.975 260.690 -53.345 260.860 ;
        RECT -44.190 260.755 -43.960 261.505 ;
        RECT -45.455 260.725 -43.495 260.755 ;
        RECT -56.975 260.665 -56.465 260.690 ;
        RECT -54.795 260.675 -53.345 260.690 ;
        RECT -56.975 259.905 -56.785 260.665 ;
        RECT -53.570 260.395 -53.345 260.675 ;
        RECT -45.475 260.555 -43.035 260.725 ;
        RECT -45.455 260.525 -43.495 260.555 ;
        RECT -54.615 260.370 -54.215 260.390 ;
        RECT -56.605 260.200 -54.215 260.370 ;
        RECT -54.615 260.165 -54.215 260.200 ;
        RECT -56.975 259.880 -56.465 259.905 ;
        RECT -56.975 259.710 -54.565 259.880 ;
        RECT -56.975 259.675 -56.465 259.710 ;
        RECT -54.395 258.830 -54.215 260.165 ;
        RECT -54.020 259.300 -53.720 260.015 ;
        RECT -53.525 259.345 -53.345 260.395 ;
        RECT -53.525 259.315 -53.100 259.345 ;
        RECT -54.590 258.825 -54.215 258.830 ;
        RECT -56.605 258.655 -54.215 258.825 ;
        RECT -54.590 258.650 -54.215 258.655 ;
        RECT -53.985 257.885 -53.805 259.300 ;
        RECT -53.525 259.145 -52.105 259.315 ;
        RECT -53.525 259.120 -53.100 259.145 ;
        RECT -53.620 258.185 -53.320 258.915 ;
        RECT -53.540 257.890 -53.360 258.185 ;
        RECT -40.525 257.865 -40.225 258.350 ;
        RECT -45.225 257.705 -44.845 257.765 ;
        RECT -45.225 257.535 -41.835 257.705 ;
        RECT -41.645 257.655 -40.225 257.865 ;
        RECT -45.225 257.485 -44.845 257.535 ;
        RECT -45.225 256.775 -45.055 257.485 ;
        RECT -41.645 257.235 -41.435 257.655 ;
        RECT -41.925 257.215 -41.435 257.235 ;
        RECT -44.875 257.045 -41.435 257.215 ;
        RECT -41.925 257.025 -41.435 257.045 ;
        RECT -45.225 256.725 -44.845 256.775 ;
        RECT -53.650 256.360 -53.350 256.605 ;
        RECT -45.225 256.555 -41.835 256.725 ;
        RECT -41.070 256.565 -40.790 256.990 ;
        RECT -45.225 256.495 -44.845 256.555 ;
        RECT -53.650 256.195 -53.345 256.360 ;
        RECT -56.975 256.130 -56.465 256.165 ;
        RECT -54.795 256.130 -53.345 256.195 ;
        RECT -56.975 255.960 -53.345 256.130 ;
        RECT -56.975 255.935 -56.465 255.960 ;
        RECT -54.795 255.945 -53.345 255.960 ;
        RECT -56.975 255.175 -56.785 255.935 ;
        RECT -53.570 255.665 -53.345 255.945 ;
        RECT -54.615 255.640 -54.215 255.660 ;
        RECT -56.605 255.470 -54.215 255.640 ;
        RECT -54.615 255.435 -54.215 255.470 ;
        RECT -56.975 255.150 -56.465 255.175 ;
        RECT -56.975 254.980 -54.565 255.150 ;
        RECT -56.975 254.945 -56.465 254.980 ;
        RECT -54.395 254.100 -54.215 255.435 ;
        RECT -54.020 254.570 -53.720 255.285 ;
        RECT -53.525 254.615 -53.345 255.665 ;
        RECT -45.225 255.715 -45.055 256.495 ;
        RECT -41.300 256.265 -40.790 256.565 ;
        RECT -41.890 256.160 -41.480 256.175 ;
        RECT -44.875 255.990 -41.480 256.160 ;
        RECT -41.890 255.965 -41.480 255.990 ;
        RECT -45.225 255.670 -44.845 255.715 ;
        RECT -45.225 255.500 -41.835 255.670 ;
        RECT -45.225 255.450 -44.845 255.500 ;
        RECT -41.665 255.195 -41.480 255.965 ;
        RECT -41.885 255.180 -41.480 255.195 ;
        RECT -44.875 255.010 -41.480 255.180 ;
        RECT -41.885 254.985 -41.480 255.010 ;
        RECT -53.525 254.585 -53.100 254.615 ;
        RECT -54.590 254.095 -54.215 254.100 ;
        RECT -56.605 253.925 -54.215 254.095 ;
        RECT -54.590 253.920 -54.215 253.925 ;
        RECT -53.985 252.460 -53.805 254.570 ;
        RECT -53.525 254.415 -52.105 254.585 ;
        RECT -53.525 254.390 -53.100 254.415 ;
        RECT -53.620 253.455 -53.320 254.185 ;
        RECT -41.665 254.135 -41.480 254.985 ;
        RECT -41.920 254.120 -41.480 254.135 ;
        RECT -44.875 253.950 -41.480 254.120 ;
        RECT -41.920 253.930 -41.480 253.950 ;
        RECT -55.060 252.280 -53.805 252.460 ;
        RECT -84.505 42.780 -83.830 218.620 ;
        RECT -83.320 126.530 -82.640 251.250 ;
        RECT -64.665 249.265 -63.980 249.270 ;
        RECT -66.745 249.260 -62.005 249.265 ;
        RECT -66.745 249.230 -61.995 249.260 ;
        RECT -66.895 249.025 -61.995 249.230 ;
        RECT -66.895 248.390 -66.525 249.025 ;
        RECT -64.665 248.970 -63.980 249.025 ;
        RECT -62.190 248.850 -61.995 249.025 ;
        RECT -62.300 248.700 -61.950 248.850 ;
        RECT -62.605 248.670 -61.585 248.700 ;
        RECT -63.065 248.500 -60.625 248.670 ;
        RECT -62.605 248.470 -61.585 248.500 ;
        RECT -68.235 248.180 -66.275 248.210 ;
        RECT -68.255 248.010 -65.815 248.180 ;
        RECT -68.235 247.980 -66.275 248.010 ;
        RECT -66.970 247.230 -66.740 247.980 ;
        RECT -62.140 247.720 -61.910 248.470 ;
        RECT -62.605 247.690 -61.585 247.720 ;
        RECT -67.295 247.200 -66.275 247.230 ;
        RECT -68.255 247.030 -65.815 247.200 ;
        RECT -67.295 247.000 -66.275 247.030 ;
        RECT -66.970 246.250 -66.740 247.000 ;
        RECT -67.295 246.220 -66.275 246.250 ;
        RECT -68.255 246.050 -65.815 246.220 ;
        RECT -67.295 246.020 -66.275 246.050 ;
        RECT -66.930 245.815 -66.580 246.020 ;
        RECT -67.825 245.585 -66.580 245.815 ;
        RECT -64.090 245.585 -63.895 247.615 ;
        RECT -63.065 247.520 -60.625 247.690 ;
        RECT -62.605 247.490 -61.585 247.520 ;
        RECT -62.140 246.740 -61.910 247.490 ;
        RECT -62.605 246.710 -60.645 246.740 ;
        RECT -63.065 246.540 -60.625 246.710 ;
        RECT -62.605 246.510 -60.645 246.540 ;
        RECT -67.825 245.100 -67.580 245.585 ;
        RECT -66.835 245.220 -65.805 245.405 ;
        RECT -66.840 245.105 -65.805 245.220 ;
        RECT -68.145 244.815 -67.325 245.100 ;
        RECT -66.840 245.045 -66.525 245.105 ;
        RECT -66.895 244.205 -66.525 245.045 ;
        RECT -64.130 244.925 -63.830 245.585 ;
        RECT -62.355 245.490 -61.985 246.330 ;
        RECT -68.235 243.995 -66.275 244.025 ;
        RECT -68.255 243.825 -65.815 243.995 ;
        RECT -68.235 243.795 -66.275 243.825 ;
        RECT -66.970 243.045 -66.740 243.795 ;
        RECT -67.295 243.015 -66.275 243.045 ;
        RECT -68.255 242.845 -65.815 243.015 ;
        RECT -67.295 242.815 -66.275 242.845 ;
        RECT -66.970 242.065 -66.740 242.815 ;
        RECT -67.295 242.035 -66.275 242.065 ;
        RECT -68.255 241.865 -65.815 242.035 ;
        RECT -67.295 241.835 -66.275 241.865 ;
        RECT -66.930 241.560 -66.580 241.835 ;
        RECT -67.890 241.195 -66.580 241.560 ;
        RECT -67.890 241.190 -67.050 241.195 ;
        RECT -68.520 240.940 -68.125 240.945 ;
        RECT -67.755 240.940 -65.975 240.970 ;
        RECT -65.625 240.940 -65.165 240.965 ;
        RECT -68.520 240.770 -65.165 240.940 ;
        RECT -68.520 240.765 -68.125 240.770 ;
        RECT -68.520 239.965 -68.350 240.765 ;
        RECT -67.755 240.735 -65.975 240.770 ;
        RECT -65.625 240.745 -65.165 240.770 ;
        RECT -67.720 240.450 -67.290 240.455 ;
        RECT -68.180 240.280 -67.290 240.450 ;
        RECT -67.720 240.275 -67.290 240.280 ;
        RECT -68.520 239.960 -68.075 239.965 ;
        RECT -68.520 239.790 -67.640 239.960 ;
        RECT -68.520 239.755 -68.075 239.790 ;
        RECT -68.520 238.995 -68.350 239.755 ;
        RECT -68.180 239.465 -67.640 239.470 ;
        RECT -67.460 239.465 -67.290 240.275 ;
        RECT -67.020 240.110 -66.650 240.735 ;
        RECT -66.455 240.450 -66.080 240.470 ;
        RECT -66.455 240.280 -65.565 240.450 ;
        RECT -66.455 240.265 -66.080 240.280 ;
        RECT -68.180 239.300 -67.290 239.465 ;
        RECT -67.730 239.285 -67.290 239.300 ;
        RECT -68.520 238.980 -68.070 238.995 ;
        RECT -68.520 238.810 -67.640 238.980 ;
        RECT -68.520 238.785 -68.070 238.810 ;
        RECT -68.520 238.015 -68.350 238.785 ;
        RECT -67.460 238.495 -67.290 239.285 ;
        RECT -67.730 238.490 -67.290 238.495 ;
        RECT -68.180 238.320 -67.290 238.490 ;
        RECT -67.730 238.315 -67.290 238.320 ;
        RECT -67.460 238.190 -67.290 238.315 ;
        RECT -66.455 239.480 -66.285 240.265 ;
        RECT -65.335 239.985 -65.165 240.745 ;
        RECT -65.680 239.960 -65.165 239.985 ;
        RECT -66.105 239.790 -65.165 239.960 ;
        RECT -65.680 239.765 -65.165 239.790 ;
        RECT -66.455 239.470 -66.040 239.480 ;
        RECT -66.455 239.300 -65.565 239.470 ;
        RECT -66.455 239.275 -66.040 239.300 ;
        RECT -66.455 238.510 -66.285 239.275 ;
        RECT -65.335 239.005 -65.165 239.765 ;
        RECT -65.680 238.980 -65.165 239.005 ;
        RECT -66.105 238.810 -65.165 238.980 ;
        RECT -65.680 238.785 -65.165 238.810 ;
        RECT -66.455 238.490 -66.040 238.510 ;
        RECT -66.455 238.320 -65.565 238.490 ;
        RECT -66.455 238.305 -66.040 238.320 ;
        RECT -66.455 238.190 -66.285 238.305 ;
        RECT -68.520 238.000 -68.095 238.015 ;
        RECT -68.520 237.830 -67.640 238.000 ;
        RECT -68.520 237.805 -68.095 237.830 ;
        RECT -67.460 237.525 -66.285 238.190 ;
        RECT -65.335 238.020 -65.165 238.785 ;
        RECT -65.625 238.000 -65.165 238.020 ;
        RECT -66.105 237.830 -65.165 238.000 ;
        RECT -65.625 237.800 -65.165 237.830 ;
        RECT -67.680 237.510 -66.035 237.525 ;
        RECT -68.180 237.340 -65.565 237.510 ;
        RECT -67.680 237.320 -66.035 237.340 ;
        RECT -67.680 237.315 -66.250 237.320 ;
        RECT -66.755 236.860 -66.455 237.315 ;
        RECT -66.860 235.730 -66.560 235.840 ;
        RECT -66.895 234.890 -66.525 235.730 ;
        RECT -68.235 234.680 -66.275 234.710 ;
        RECT -68.255 234.510 -65.815 234.680 ;
        RECT -68.235 234.480 -66.275 234.510 ;
        RECT -66.970 233.730 -66.740 234.480 ;
        RECT -67.295 233.700 -66.275 233.730 ;
        RECT -68.255 233.530 -65.815 233.700 ;
        RECT -67.295 233.500 -66.275 233.530 ;
        RECT -66.970 232.750 -66.740 233.500 ;
        RECT -67.295 232.720 -66.275 232.750 ;
        RECT -68.255 232.550 -65.815 232.720 ;
        RECT -67.295 232.520 -66.275 232.550 ;
        RECT -66.930 232.340 -66.580 232.520 ;
        RECT -67.885 232.030 -66.580 232.340 ;
        RECT -67.885 231.600 -67.575 232.030 ;
        RECT -68.145 231.315 -67.325 231.600 ;
        RECT -68.235 230.495 -66.275 230.525 ;
        RECT -68.255 230.325 -65.815 230.495 ;
        RECT -68.235 230.295 -66.275 230.325 ;
        RECT -66.970 229.545 -66.740 230.295 ;
        RECT -67.295 229.515 -66.275 229.545 ;
        RECT -68.255 229.345 -65.815 229.515 ;
        RECT -67.295 229.315 -66.275 229.345 ;
        RECT -66.970 228.565 -66.740 229.315 ;
        RECT -67.295 228.535 -66.275 228.565 ;
        RECT -68.255 228.365 -65.815 228.535 ;
        RECT -67.295 228.335 -66.275 228.365 ;
        RECT -66.930 228.060 -66.580 228.335 ;
        RECT -67.890 227.695 -66.580 228.060 ;
        RECT -67.890 227.690 -67.050 227.695 ;
        RECT -68.520 227.440 -68.125 227.445 ;
        RECT -67.755 227.440 -65.975 227.470 ;
        RECT -65.625 227.440 -65.165 227.465 ;
        RECT -68.520 227.270 -65.165 227.440 ;
        RECT -68.520 227.265 -68.125 227.270 ;
        RECT -68.520 226.465 -68.350 227.265 ;
        RECT -67.755 227.235 -65.975 227.270 ;
        RECT -65.625 227.245 -65.165 227.270 ;
        RECT -67.720 226.950 -67.290 226.955 ;
        RECT -68.180 226.780 -67.290 226.950 ;
        RECT -67.720 226.775 -67.290 226.780 ;
        RECT -68.520 226.460 -68.075 226.465 ;
        RECT -68.520 226.290 -67.640 226.460 ;
        RECT -68.520 226.255 -68.075 226.290 ;
        RECT -68.520 225.495 -68.350 226.255 ;
        RECT -68.180 225.965 -67.640 225.970 ;
        RECT -67.460 225.965 -67.290 226.775 ;
        RECT -67.020 226.610 -66.650 227.235 ;
        RECT -66.455 226.950 -66.080 226.970 ;
        RECT -66.455 226.780 -65.565 226.950 ;
        RECT -66.455 226.765 -66.080 226.780 ;
        RECT -68.180 225.800 -67.290 225.965 ;
        RECT -67.730 225.785 -67.290 225.800 ;
        RECT -68.520 225.480 -68.070 225.495 ;
        RECT -68.520 225.310 -67.640 225.480 ;
        RECT -68.520 225.285 -68.070 225.310 ;
        RECT -68.520 224.515 -68.350 225.285 ;
        RECT -67.460 224.995 -67.290 225.785 ;
        RECT -67.730 224.990 -67.290 224.995 ;
        RECT -68.180 224.820 -67.290 224.990 ;
        RECT -67.730 224.815 -67.290 224.820 ;
        RECT -67.460 224.690 -67.290 224.815 ;
        RECT -66.455 225.980 -66.285 226.765 ;
        RECT -65.335 226.485 -65.165 227.245 ;
        RECT -65.680 226.460 -65.165 226.485 ;
        RECT -66.105 226.290 -65.165 226.460 ;
        RECT -65.680 226.265 -65.165 226.290 ;
        RECT -66.455 225.970 -66.040 225.980 ;
        RECT -66.455 225.800 -65.565 225.970 ;
        RECT -66.455 225.775 -66.040 225.800 ;
        RECT -66.455 225.010 -66.285 225.775 ;
        RECT -65.335 225.505 -65.165 226.265 ;
        RECT -65.680 225.480 -65.165 225.505 ;
        RECT -66.105 225.310 -65.165 225.480 ;
        RECT -65.680 225.285 -65.165 225.310 ;
        RECT -66.455 224.990 -66.040 225.010 ;
        RECT -66.455 224.820 -65.565 224.990 ;
        RECT -66.455 224.805 -66.040 224.820 ;
        RECT -66.455 224.690 -66.285 224.805 ;
        RECT -68.520 224.500 -68.095 224.515 ;
        RECT -68.520 224.330 -67.640 224.500 ;
        RECT -68.520 224.305 -68.095 224.330 ;
        RECT -67.460 224.025 -66.285 224.690 ;
        RECT -65.335 224.520 -65.165 225.285 ;
        RECT -65.625 224.500 -65.165 224.520 ;
        RECT -66.105 224.330 -65.165 224.500 ;
        RECT -65.625 224.300 -65.165 224.330 ;
        RECT -67.680 224.010 -66.035 224.025 ;
        RECT -68.180 223.840 -65.565 224.010 ;
        RECT -67.680 223.820 -66.035 223.840 ;
        RECT -67.680 223.815 -66.250 223.820 ;
        RECT -66.745 223.440 -66.445 223.815 ;
        RECT -64.090 222.970 -63.895 244.925 ;
        RECT -62.280 244.505 -62.015 245.490 ;
        RECT -62.630 244.500 -61.200 244.505 ;
        RECT -62.845 244.480 -61.200 244.500 ;
        RECT -63.315 244.310 -60.700 244.480 ;
        RECT -62.845 244.295 -61.200 244.310 ;
        RECT -63.715 243.990 -63.255 244.020 ;
        RECT -63.715 243.820 -62.775 243.990 ;
        RECT -63.715 243.800 -63.255 243.820 ;
        RECT -63.715 243.035 -63.545 243.800 ;
        RECT -62.595 243.630 -61.420 244.295 ;
        RECT -60.785 243.990 -60.360 244.015 ;
        RECT -61.240 243.820 -60.360 243.990 ;
        RECT -60.785 243.805 -60.360 243.820 ;
        RECT -62.595 243.515 -62.425 243.630 ;
        RECT -62.840 243.500 -62.425 243.515 ;
        RECT -63.315 243.330 -62.425 243.500 ;
        RECT -62.840 243.310 -62.425 243.330 ;
        RECT -63.715 243.010 -63.200 243.035 ;
        RECT -63.715 242.840 -62.775 243.010 ;
        RECT -63.715 242.815 -63.200 242.840 ;
        RECT -63.715 242.055 -63.545 242.815 ;
        RECT -62.595 242.545 -62.425 243.310 ;
        RECT -62.840 242.520 -62.425 242.545 ;
        RECT -63.315 242.350 -62.425 242.520 ;
        RECT -62.840 242.340 -62.425 242.350 ;
        RECT -63.715 242.030 -63.200 242.055 ;
        RECT -63.715 241.860 -62.775 242.030 ;
        RECT -63.715 241.835 -63.200 241.860 ;
        RECT -63.715 241.075 -63.545 241.835 ;
        RECT -62.595 241.555 -62.425 242.340 ;
        RECT -61.590 243.505 -61.420 243.630 ;
        RECT -61.590 243.500 -61.150 243.505 ;
        RECT -61.590 243.330 -60.700 243.500 ;
        RECT -61.590 243.325 -61.150 243.330 ;
        RECT -61.590 242.535 -61.420 243.325 ;
        RECT -60.530 243.035 -60.360 243.805 ;
        RECT -60.810 243.010 -60.360 243.035 ;
        RECT -61.240 242.840 -60.360 243.010 ;
        RECT -60.810 242.825 -60.360 242.840 ;
        RECT -61.590 242.520 -61.150 242.535 ;
        RECT -61.590 242.355 -60.700 242.520 ;
        RECT -62.800 241.540 -62.425 241.555 ;
        RECT -63.315 241.370 -62.425 241.540 ;
        RECT -62.800 241.350 -62.425 241.370 ;
        RECT -62.230 241.085 -61.860 241.710 ;
        RECT -61.590 241.545 -61.420 242.355 ;
        RECT -61.240 242.350 -60.700 242.355 ;
        RECT -60.530 242.065 -60.360 242.825 ;
        RECT -60.805 242.030 -60.360 242.065 ;
        RECT -61.240 241.860 -60.360 242.030 ;
        RECT -60.805 241.855 -60.360 241.860 ;
        RECT -61.590 241.540 -61.160 241.545 ;
        RECT -61.590 241.370 -60.700 241.540 ;
        RECT -61.590 241.365 -61.160 241.370 ;
        RECT -63.715 241.050 -63.255 241.075 ;
        RECT -62.905 241.050 -61.125 241.085 ;
        RECT -60.530 241.055 -60.360 241.855 ;
        RECT -60.755 241.050 -60.360 241.055 ;
        RECT -63.715 240.880 -60.360 241.050 ;
        RECT -63.715 240.855 -63.255 240.880 ;
        RECT -62.905 240.850 -61.125 240.880 ;
        RECT -60.755 240.875 -60.360 240.880 ;
        RECT -61.830 240.625 -60.990 240.630 ;
        RECT -62.300 240.260 -60.990 240.625 ;
        RECT -62.300 239.985 -61.950 240.260 ;
        RECT -62.605 239.955 -61.585 239.985 ;
        RECT -63.065 239.785 -60.625 239.955 ;
        RECT -62.605 239.755 -61.585 239.785 ;
        RECT -62.140 239.005 -61.910 239.755 ;
        RECT -62.605 238.975 -61.585 239.005 ;
        RECT -63.065 238.805 -60.625 238.975 ;
        RECT -62.605 238.775 -61.585 238.805 ;
        RECT -62.140 238.025 -61.910 238.775 ;
        RECT -62.605 237.995 -60.645 238.025 ;
        RECT -63.065 237.825 -60.625 237.995 ;
        RECT -62.605 237.795 -60.645 237.825 ;
        RECT -55.060 237.785 -54.250 252.280 ;
        RECT -53.540 251.765 -53.360 253.455 ;
        RECT -56.430 237.230 -54.250 237.785 ;
        RECT -61.555 236.720 -60.735 237.005 ;
        RECT -61.350 235.925 -61.125 236.720 ;
        RECT -62.245 235.900 -61.125 235.925 ;
        RECT -62.820 235.700 -61.125 235.900 ;
        RECT -62.820 235.600 -62.020 235.700 ;
        RECT -62.245 235.350 -62.020 235.600 ;
        RECT -62.300 235.200 -61.950 235.350 ;
        RECT -62.605 235.170 -61.585 235.200 ;
        RECT -63.065 235.000 -60.625 235.170 ;
        RECT -62.605 234.970 -61.585 235.000 ;
        RECT -62.140 234.220 -61.910 234.970 ;
        RECT -62.605 234.190 -61.585 234.220 ;
        RECT -63.065 234.020 -60.625 234.190 ;
        RECT -62.605 233.990 -61.585 234.020 ;
        RECT -62.140 233.240 -61.910 233.990 ;
        RECT -62.605 233.210 -60.645 233.240 ;
        RECT -63.065 233.040 -60.625 233.210 ;
        RECT -62.605 233.010 -60.645 233.040 ;
        RECT -62.355 231.990 -61.985 232.830 ;
        RECT -62.315 231.005 -62.030 231.990 ;
        RECT -62.630 231.000 -61.200 231.005 ;
        RECT -62.845 230.995 -61.200 231.000 ;
        RECT -63.455 230.980 -61.200 230.995 ;
        RECT -63.455 230.810 -60.700 230.980 ;
        RECT -63.455 230.795 -61.200 230.810 ;
        RECT -63.455 230.765 -62.795 230.795 ;
        RECT -63.715 230.490 -63.255 230.520 ;
        RECT -63.715 230.320 -62.775 230.490 ;
        RECT -63.715 230.300 -63.255 230.320 ;
        RECT -63.715 229.535 -63.545 230.300 ;
        RECT -62.595 230.130 -61.420 230.795 ;
        RECT -60.785 230.490 -60.360 230.515 ;
        RECT -61.240 230.320 -60.360 230.490 ;
        RECT -60.785 230.305 -60.360 230.320 ;
        RECT -62.595 230.015 -62.425 230.130 ;
        RECT -62.840 230.000 -62.425 230.015 ;
        RECT -63.315 229.830 -62.425 230.000 ;
        RECT -62.840 229.810 -62.425 229.830 ;
        RECT -63.715 229.510 -63.200 229.535 ;
        RECT -63.715 229.340 -62.775 229.510 ;
        RECT -63.715 229.315 -63.200 229.340 ;
        RECT -63.715 228.555 -63.545 229.315 ;
        RECT -62.595 229.045 -62.425 229.810 ;
        RECT -62.840 229.020 -62.425 229.045 ;
        RECT -63.315 228.850 -62.425 229.020 ;
        RECT -62.840 228.840 -62.425 228.850 ;
        RECT -63.715 228.530 -63.200 228.555 ;
        RECT -63.715 228.360 -62.775 228.530 ;
        RECT -63.715 228.335 -63.200 228.360 ;
        RECT -63.715 227.575 -63.545 228.335 ;
        RECT -62.595 228.055 -62.425 228.840 ;
        RECT -61.590 230.005 -61.420 230.130 ;
        RECT -61.590 230.000 -61.150 230.005 ;
        RECT -61.590 229.830 -60.700 230.000 ;
        RECT -61.590 229.825 -61.150 229.830 ;
        RECT -61.590 229.035 -61.420 229.825 ;
        RECT -60.530 229.535 -60.360 230.305 ;
        RECT -60.810 229.510 -60.360 229.535 ;
        RECT -61.240 229.340 -60.360 229.510 ;
        RECT -60.810 229.325 -60.360 229.340 ;
        RECT -61.590 229.020 -61.150 229.035 ;
        RECT -61.590 228.855 -60.700 229.020 ;
        RECT -62.800 228.040 -62.425 228.055 ;
        RECT -63.315 227.870 -62.425 228.040 ;
        RECT -62.800 227.850 -62.425 227.870 ;
        RECT -62.230 227.585 -61.860 228.210 ;
        RECT -61.590 228.045 -61.420 228.855 ;
        RECT -61.240 228.850 -60.700 228.855 ;
        RECT -60.530 228.565 -60.360 229.325 ;
        RECT -60.805 228.530 -60.360 228.565 ;
        RECT -61.240 228.360 -60.360 228.530 ;
        RECT -60.805 228.355 -60.360 228.360 ;
        RECT -61.590 228.040 -61.160 228.045 ;
        RECT -61.590 227.870 -60.700 228.040 ;
        RECT -61.590 227.865 -61.160 227.870 ;
        RECT -63.715 227.550 -63.255 227.575 ;
        RECT -62.905 227.550 -61.125 227.585 ;
        RECT -60.530 227.555 -60.360 228.355 ;
        RECT -60.755 227.550 -60.360 227.555 ;
        RECT -63.715 227.380 -60.360 227.550 ;
        RECT -63.715 227.355 -63.255 227.380 ;
        RECT -62.905 227.350 -61.125 227.380 ;
        RECT -60.755 227.375 -60.360 227.380 ;
        RECT -61.830 227.125 -60.990 227.130 ;
        RECT -62.300 226.760 -60.990 227.125 ;
        RECT -62.300 226.485 -61.950 226.760 ;
        RECT -62.605 226.455 -61.585 226.485 ;
        RECT -63.065 226.285 -60.625 226.455 ;
        RECT -62.605 226.255 -61.585 226.285 ;
        RECT -62.140 225.505 -61.910 226.255 ;
        RECT -62.605 225.475 -61.585 225.505 ;
        RECT -63.065 225.305 -60.625 225.475 ;
        RECT -62.605 225.275 -61.585 225.305 ;
        RECT -62.140 224.525 -61.910 225.275 ;
        RECT -62.605 224.495 -60.645 224.525 ;
        RECT -63.065 224.325 -60.625 224.495 ;
        RECT -62.605 224.295 -60.645 224.325 ;
        RECT -62.355 223.275 -61.985 224.115 ;
        RECT -62.330 223.100 -62.040 223.275 ;
        RECT -61.555 223.220 -60.735 223.505 ;
        RECT -64.140 222.310 -63.840 222.970 ;
        RECT -62.270 222.815 -62.060 223.100 ;
        RECT -62.700 222.515 -62.040 222.815 ;
        RECT -62.270 222.225 -62.060 222.515 ;
        RECT -62.300 222.075 -61.950 222.225 ;
        RECT -62.605 222.045 -61.585 222.075 ;
        RECT -63.065 221.875 -60.625 222.045 ;
        RECT -62.605 221.845 -61.585 221.875 ;
        RECT -62.140 221.095 -61.910 221.845 ;
        RECT -62.605 221.065 -61.585 221.095 ;
        RECT -63.065 220.895 -60.625 221.065 ;
        RECT -62.605 220.865 -61.585 220.895 ;
        RECT -62.140 220.115 -61.910 220.865 ;
        RECT -62.605 220.085 -60.645 220.115 ;
        RECT -63.065 219.915 -60.625 220.085 ;
        RECT -62.605 219.885 -60.645 219.915 ;
        RECT -56.430 211.510 -55.875 237.230 ;
        RECT -55.060 231.875 -54.250 237.230 ;
        RECT -53.690 230.280 -53.220 251.765 ;
        RECT -41.300 245.600 -41.095 256.265 ;
        RECT -40.435 255.610 -40.225 257.655 ;
        RECT -40.435 255.590 -39.970 255.610 ;
        RECT -40.435 255.420 -39.015 255.590 ;
        RECT -40.435 255.400 -39.970 255.420 ;
        RECT -40.910 254.665 -40.630 255.390 ;
        RECT -40.855 246.885 -40.650 254.665 ;
        RECT -40.435 254.630 -40.225 255.400 ;
        RECT -40.435 254.610 -39.970 254.630 ;
        RECT -40.435 254.440 -39.015 254.610 ;
        RECT -40.435 254.420 -39.970 254.440 ;
        RECT -40.435 253.020 -40.155 253.745 ;
        RECT -40.395 247.880 -40.190 253.020 ;
        RECT -38.525 247.880 -37.770 247.920 ;
        RECT -22.020 247.880 -21.115 248.340 ;
        RECT -40.395 247.435 -21.115 247.880 ;
        RECT -22.020 247.355 -21.115 247.435 ;
        RECT -24.395 246.885 -23.350 247.040 ;
        RECT -40.855 246.225 -23.350 246.885 ;
        RECT -26.535 245.600 -25.180 245.645 ;
        RECT -24.395 245.635 -23.350 246.225 ;
        RECT -41.300 244.960 -25.180 245.600 ;
        RECT -49.475 243.115 -48.575 244.220 ;
        RECT -38.525 243.785 -37.770 244.550 ;
        RECT -49.365 239.245 -48.715 243.115 ;
        RECT -39.820 240.375 -39.000 240.865 ;
        RECT -50.755 238.830 -48.715 239.245 ;
        RECT -53.690 229.865 -51.860 230.280 ;
        RECT -53.690 228.390 -53.220 229.865 ;
        RECT -54.025 226.965 -52.930 228.390 ;
        RECT -56.480 211.165 -55.785 211.510 ;
        RECT -52.275 210.695 -51.860 229.865 ;
        RECT -50.755 212.325 -50.340 238.830 ;
        RECT -49.365 236.885 -48.715 238.830 ;
        RECT -50.025 234.315 -47.900 236.885 ;
        RECT -39.685 213.065 -39.070 240.375 ;
        RECT -39.705 212.815 -39.040 213.065 ;
        RECT -39.685 212.770 -39.070 212.815 ;
        RECT -50.815 212.005 -50.225 212.325 ;
        RECT -52.300 210.400 -51.825 210.695 ;
        RECT -38.340 208.995 -37.965 243.785 ;
        RECT -36.305 242.470 -34.815 243.805 ;
        RECT -30.595 242.635 -29.895 244.095 ;
        RECT -26.535 243.835 -25.180 244.960 ;
        RECT -36.170 215.745 -34.995 242.470 ;
        RECT -38.370 207.905 -37.925 208.995 ;
        RECT -30.595 207.765 -29.900 242.635 ;
        RECT -26.270 207.705 -25.410 243.835 ;
        RECT -27.095 206.705 -25.240 207.705 ;
        RECT -67.470 203.200 -67.200 203.895 ;
        RECT -56.215 203.250 -55.945 203.945 ;
        RECT -38.465 203.250 -38.195 203.945 ;
        RECT -27.210 203.200 -26.940 203.895 ;
        RECT -56.860 203.005 -54.690 203.030 ;
        RECT -39.720 203.005 -37.550 203.030 ;
        RECT -68.115 202.955 -65.945 202.980 ;
        RECT -69.070 202.785 -65.000 202.955 ;
        RECT -57.815 202.835 -53.745 203.005 ;
        RECT -40.665 202.835 -36.595 203.005 ;
        RECT -28.465 202.955 -26.295 202.980 ;
        RECT -56.860 202.815 -54.690 202.835 ;
        RECT -39.720 202.815 -37.550 202.835 ;
        RECT -68.115 202.765 -65.945 202.785 ;
        RECT -67.130 202.265 -66.900 202.765 ;
        RECT -55.875 202.315 -55.645 202.815 ;
        RECT -38.765 202.315 -38.535 202.815 ;
        RECT -29.410 202.785 -25.340 202.955 ;
        RECT -28.465 202.765 -26.295 202.785 ;
        RECT -27.510 202.265 -27.280 202.765 ;
        RECT -56.850 201.460 -54.700 201.480 ;
        RECT -39.710 201.460 -37.560 201.480 ;
        RECT -68.105 201.410 -65.955 201.430 ;
        RECT -69.070 201.240 -65.000 201.410 ;
        RECT -57.815 201.290 -53.745 201.460 ;
        RECT -40.665 201.290 -36.595 201.460 ;
        RECT -28.455 201.410 -26.305 201.430 ;
        RECT -56.850 201.265 -54.700 201.290 ;
        RECT -39.710 201.265 -37.560 201.290 ;
        RECT -68.105 201.215 -65.955 201.240 ;
        RECT -67.500 200.125 -67.230 200.820 ;
        RECT -66.410 200.735 -66.180 201.215 ;
        RECT -66.625 200.180 -65.000 200.350 ;
        RECT -69.070 199.690 -67.315 199.860 ;
        RECT -69.070 198.710 -67.685 198.880 ;
        RECT -67.855 197.980 -67.685 198.710 ;
        RECT -69.760 197.810 -67.685 197.980 ;
        RECT -69.760 195.490 -69.590 197.810 ;
        RECT -67.485 197.630 -67.315 199.690 ;
        RECT -66.625 198.880 -66.455 200.180 ;
        RECT -56.245 200.175 -55.975 200.870 ;
        RECT -55.155 200.785 -54.925 201.265 ;
        RECT -39.485 200.785 -39.255 201.265 ;
        RECT -29.410 201.240 -25.340 201.410 ;
        RECT -28.455 201.215 -26.305 201.240 ;
        RECT -55.370 200.230 -53.745 200.400 ;
        RECT -40.665 200.230 -39.040 200.400 ;
        RECT -65.085 199.860 -64.635 199.870 ;
        RECT -66.040 199.690 -64.635 199.860 ;
        RECT -57.815 199.740 -56.060 199.910 ;
        RECT -67.130 198.080 -66.860 198.775 ;
        RECT -66.625 198.710 -65.000 198.880 ;
        RECT -66.625 197.715 -66.455 198.710 ;
        RECT -69.415 197.460 -67.315 197.630 ;
        RECT -67.105 197.545 -66.455 197.715 ;
        RECT -66.190 198.220 -65.000 198.390 ;
        RECT -69.415 197.070 -69.245 197.460 ;
        RECT -67.105 197.155 -66.935 197.545 ;
        RECT -69.415 196.900 -68.030 197.070 ;
        RECT -67.850 196.985 -66.935 197.155 ;
        RECT -66.190 197.070 -65.995 198.220 ;
        RECT -69.415 196.090 -69.245 196.900 ;
        RECT -67.850 196.580 -67.680 196.985 ;
        RECT -66.190 196.900 -65.000 197.070 ;
        RECT -66.190 196.890 -65.995 196.900 ;
        RECT -69.070 196.410 -67.680 196.580 ;
        RECT -69.415 195.920 -68.030 196.090 ;
        RECT -69.760 195.320 -68.030 195.490 ;
        RECT -69.760 194.510 -69.590 195.320 ;
        RECT -67.850 195.000 -67.680 196.410 ;
        RECT -69.070 194.830 -67.680 195.000 ;
        RECT -69.760 194.340 -68.030 194.510 ;
        RECT -67.850 192.920 -67.680 194.830 ;
        RECT -67.280 194.335 -67.010 195.030 ;
        RECT -64.815 195.000 -64.635 199.690 ;
        RECT -57.815 198.760 -56.430 198.930 ;
        RECT -56.600 198.030 -56.430 198.760 ;
        RECT -66.040 194.830 -64.635 195.000 ;
        RECT -58.505 197.860 -56.430 198.030 ;
        RECT -58.505 195.540 -58.335 197.860 ;
        RECT -56.230 197.680 -56.060 199.740 ;
        RECT -55.370 198.930 -55.200 200.230 ;
        RECT -53.830 199.910 -53.380 199.920 ;
        RECT -54.785 199.740 -53.380 199.910 ;
        RECT -55.875 198.130 -55.605 198.825 ;
        RECT -55.370 198.760 -53.745 198.930 ;
        RECT -55.370 197.765 -55.200 198.760 ;
        RECT -58.160 197.510 -56.060 197.680 ;
        RECT -55.850 197.595 -55.200 197.765 ;
        RECT -54.935 198.270 -53.745 198.440 ;
        RECT -58.160 197.120 -57.990 197.510 ;
        RECT -55.850 197.205 -55.680 197.595 ;
        RECT -58.160 196.950 -56.775 197.120 ;
        RECT -56.595 197.035 -55.680 197.205 ;
        RECT -54.935 197.120 -54.740 198.270 ;
        RECT -58.160 196.140 -57.990 196.950 ;
        RECT -56.595 196.630 -56.425 197.035 ;
        RECT -54.935 196.950 -53.745 197.120 ;
        RECT -54.935 196.940 -54.740 196.950 ;
        RECT -57.815 196.460 -56.425 196.630 ;
        RECT -58.160 195.970 -56.775 196.140 ;
        RECT -58.505 195.370 -56.775 195.540 ;
        RECT -58.505 194.560 -58.335 195.370 ;
        RECT -56.595 195.050 -56.425 196.460 ;
        RECT -57.815 194.880 -56.425 195.050 ;
        RECT -58.505 194.390 -56.775 194.560 ;
        RECT -56.595 194.135 -56.425 194.880 ;
        RECT -56.025 194.385 -55.755 195.080 ;
        RECT -53.560 195.050 -53.380 199.740 ;
        RECT -54.785 194.880 -53.380 195.050 ;
        RECT -41.030 199.910 -40.580 199.920 ;
        RECT -41.030 199.740 -39.625 199.910 ;
        RECT -41.030 195.050 -40.850 199.740 ;
        RECT -39.210 198.930 -39.040 200.230 ;
        RECT -38.435 200.175 -38.165 200.870 ;
        RECT -28.230 200.735 -28.000 201.215 ;
        RECT -29.410 200.180 -27.785 200.350 ;
        RECT -40.665 198.760 -39.040 198.930 ;
        RECT -38.350 199.740 -36.595 199.910 ;
        RECT -29.775 199.860 -29.325 199.870 ;
        RECT -40.665 198.270 -39.475 198.440 ;
        RECT -39.670 197.120 -39.475 198.270 ;
        RECT -39.210 197.765 -39.040 198.760 ;
        RECT -38.805 198.130 -38.535 198.825 ;
        RECT -39.210 197.595 -38.560 197.765 ;
        RECT -40.665 196.950 -39.475 197.120 ;
        RECT -38.730 197.205 -38.560 197.595 ;
        RECT -38.350 197.680 -38.180 199.740 ;
        RECT -29.775 199.690 -28.370 199.860 ;
        RECT -37.980 198.760 -36.595 198.930 ;
        RECT -37.980 198.030 -37.810 198.760 ;
        RECT -37.980 197.860 -35.905 198.030 ;
        RECT -38.350 197.510 -36.250 197.680 ;
        RECT -38.730 197.035 -37.815 197.205 ;
        RECT -36.420 197.120 -36.250 197.510 ;
        RECT -39.670 196.940 -39.475 196.950 ;
        RECT -37.985 196.630 -37.815 197.035 ;
        RECT -37.635 196.950 -36.250 197.120 ;
        RECT -37.985 196.460 -36.595 196.630 ;
        RECT -41.030 194.880 -39.625 195.050 ;
        RECT -38.655 194.385 -38.385 195.080 ;
        RECT -37.985 195.050 -37.815 196.460 ;
        RECT -36.420 196.140 -36.250 196.950 ;
        RECT -37.635 195.970 -36.250 196.140 ;
        RECT -36.075 195.540 -35.905 197.860 ;
        RECT -37.635 195.370 -35.905 195.540 ;
        RECT -37.985 194.880 -36.595 195.050 ;
        RECT -37.985 194.135 -37.815 194.880 ;
        RECT -36.075 194.560 -35.905 195.370 ;
        RECT -29.775 195.000 -29.595 199.690 ;
        RECT -27.955 198.880 -27.785 200.180 ;
        RECT -27.180 200.125 -26.910 200.820 ;
        RECT -29.410 198.710 -27.785 198.880 ;
        RECT -27.095 199.690 -25.340 199.860 ;
        RECT -29.410 198.220 -28.220 198.390 ;
        RECT -28.415 197.070 -28.220 198.220 ;
        RECT -27.955 197.715 -27.785 198.710 ;
        RECT -27.550 198.080 -27.280 198.775 ;
        RECT -27.955 197.545 -27.305 197.715 ;
        RECT -29.410 196.900 -28.220 197.070 ;
        RECT -27.475 197.155 -27.305 197.545 ;
        RECT -27.095 197.630 -26.925 199.690 ;
        RECT -26.725 198.710 -25.340 198.880 ;
        RECT -26.725 197.980 -26.555 198.710 ;
        RECT -26.725 197.810 -24.650 197.980 ;
        RECT -27.095 197.460 -24.995 197.630 ;
        RECT -27.475 196.985 -26.560 197.155 ;
        RECT -25.165 197.070 -24.995 197.460 ;
        RECT -28.415 196.890 -28.220 196.900 ;
        RECT -26.730 196.580 -26.560 196.985 ;
        RECT -26.380 196.900 -24.995 197.070 ;
        RECT -26.730 196.410 -25.340 196.580 ;
        RECT -29.775 194.830 -28.370 195.000 ;
        RECT -37.635 194.390 -35.905 194.560 ;
        RECT -27.400 194.335 -27.130 195.030 ;
        RECT -26.730 195.000 -26.560 196.410 ;
        RECT -25.165 196.090 -24.995 196.900 ;
        RECT -26.380 195.920 -24.995 196.090 ;
        RECT -24.820 195.490 -24.650 197.810 ;
        RECT -26.380 195.320 -24.650 195.490 ;
        RECT -26.730 194.830 -25.340 195.000 ;
        RECT -63.655 193.650 -55.600 193.820 ;
        RECT -63.655 193.140 -63.485 193.650 ;
        RECT -63.195 193.300 -55.990 193.470 ;
        RECT -65.845 192.920 -65.165 192.950 ;
        RECT -67.850 192.750 -65.165 192.920 ;
        RECT -65.845 192.720 -65.165 192.750 ;
        RECT -63.685 192.460 -63.455 193.140 ;
        RECT -63.195 191.940 -63.025 193.300 ;
        RECT -56.595 193.020 -56.410 193.115 ;
        RECT -56.635 192.345 -56.365 193.020 ;
        RECT -56.595 192.340 -56.365 192.345 ;
        RECT -57.870 191.975 -56.465 192.145 ;
        RECT -63.560 191.770 -63.025 191.940 ;
        RECT -67.470 188.200 -67.200 188.895 ;
        RECT -68.115 187.955 -65.945 187.980 ;
        RECT -69.070 187.785 -65.000 187.955 ;
        RECT -68.115 187.765 -65.945 187.785 ;
        RECT -67.130 187.265 -66.900 187.765 ;
        RECT -68.105 186.410 -65.955 186.430 ;
        RECT -69.070 186.240 -65.000 186.410 ;
        RECT -68.105 186.215 -65.955 186.240 ;
        RECT -67.500 185.125 -67.230 185.820 ;
        RECT -66.410 185.735 -66.180 186.215 ;
        RECT -66.625 185.180 -65.000 185.350 ;
        RECT -69.070 184.690 -67.315 184.860 ;
        RECT -69.070 183.710 -67.685 183.880 ;
        RECT -67.855 182.980 -67.685 183.710 ;
        RECT -69.760 182.810 -67.685 182.980 ;
        RECT -69.760 180.490 -69.590 182.810 ;
        RECT -67.485 182.630 -67.315 184.690 ;
        RECT -66.625 183.880 -66.455 185.180 ;
        RECT -65.085 184.860 -64.635 184.870 ;
        RECT -66.040 184.690 -64.635 184.860 ;
        RECT -67.130 183.080 -66.860 183.775 ;
        RECT -66.625 183.710 -65.000 183.880 ;
        RECT -66.625 182.715 -66.455 183.710 ;
        RECT -69.415 182.460 -67.315 182.630 ;
        RECT -67.105 182.545 -66.455 182.715 ;
        RECT -66.190 183.220 -65.000 183.390 ;
        RECT -69.415 182.070 -69.245 182.460 ;
        RECT -67.105 182.155 -66.935 182.545 ;
        RECT -69.415 181.900 -68.030 182.070 ;
        RECT -67.850 181.985 -66.935 182.155 ;
        RECT -66.190 182.070 -65.995 183.220 ;
        RECT -69.415 181.090 -69.245 181.900 ;
        RECT -67.850 181.580 -67.680 181.985 ;
        RECT -66.190 181.900 -65.000 182.070 ;
        RECT -66.190 181.890 -65.995 181.900 ;
        RECT -69.070 181.410 -67.680 181.580 ;
        RECT -69.415 180.920 -68.030 181.090 ;
        RECT -69.760 180.320 -68.030 180.490 ;
        RECT -69.760 179.510 -69.590 180.320 ;
        RECT -67.850 180.000 -67.680 181.410 ;
        RECT -69.070 179.830 -67.680 180.000 ;
        RECT -69.760 179.340 -68.030 179.510 ;
        RECT -67.850 178.390 -67.680 179.830 ;
        RECT -67.280 179.335 -67.010 180.030 ;
        RECT -64.815 180.000 -64.635 184.690 ;
        RECT -66.040 179.830 -64.635 180.000 ;
        RECT -63.560 178.615 -63.390 191.770 ;
        RECT -56.650 191.165 -56.465 191.975 ;
        RECT -56.180 191.340 -55.990 193.300 ;
        RECT -57.870 190.995 -56.465 191.165 ;
        RECT -56.650 190.185 -56.465 190.995 ;
        RECT -56.225 190.665 -55.955 191.340 ;
        RECT -55.770 190.400 -55.600 193.650 ;
        RECT -38.810 193.650 -30.755 193.820 ;
        RECT -55.320 192.465 -53.295 192.635 ;
        RECT -41.115 192.465 -39.090 192.635 ;
        RECT -55.320 191.655 -55.150 192.465 ;
        RECT -39.260 191.655 -39.090 192.465 ;
        RECT -55.320 191.485 -53.295 191.655 ;
        RECT -41.115 191.485 -39.090 191.655 ;
        RECT -55.320 190.595 -55.145 191.485 ;
        RECT -54.830 190.915 -52.630 191.085 ;
        RECT -53.335 190.910 -52.630 190.915 ;
        RECT -55.320 190.425 -53.290 190.595 ;
        RECT -55.320 190.420 -54.830 190.425 ;
        RECT -57.870 190.015 -56.465 190.185 ;
        RECT -56.650 189.555 -56.465 190.015 ;
        RECT -55.835 189.725 -55.565 190.400 ;
        RECT -52.815 190.105 -52.630 190.910 ;
        RECT -54.830 189.935 -52.630 190.105 ;
        RECT -53.345 189.930 -52.630 189.935 ;
        RECT -56.650 189.540 -55.150 189.555 ;
        RECT -56.650 189.370 -53.290 189.540 ;
        RECT -55.775 187.345 -55.590 189.370 ;
        RECT -55.320 188.560 -55.150 189.370 ;
        RECT -52.800 189.050 -52.630 189.930 ;
        RECT -54.830 188.880 -52.630 189.050 ;
        RECT -41.780 190.915 -39.580 191.085 ;
        RECT -41.780 190.910 -41.075 190.915 ;
        RECT -41.780 190.105 -41.595 190.910 ;
        RECT -39.265 190.595 -39.090 191.485 ;
        RECT -41.120 190.425 -39.090 190.595 ;
        RECT -39.580 190.420 -39.090 190.425 ;
        RECT -38.810 190.400 -38.640 193.650 ;
        RECT -38.420 193.300 -31.215 193.470 ;
        RECT -38.420 191.340 -38.230 193.300 ;
        RECT -38.000 193.020 -37.815 193.115 ;
        RECT -38.045 192.345 -37.775 193.020 ;
        RECT -38.045 192.340 -37.815 192.345 ;
        RECT -37.945 191.975 -36.540 192.145 ;
        RECT -38.455 190.665 -38.185 191.340 ;
        RECT -37.945 191.165 -37.760 191.975 ;
        RECT -31.385 191.940 -31.215 193.300 ;
        RECT -30.925 193.140 -30.755 193.650 ;
        RECT -30.955 192.460 -30.725 193.140 ;
        RECT -29.245 192.920 -28.565 192.950 ;
        RECT -26.730 192.920 -26.560 194.830 ;
        RECT -24.820 194.510 -24.650 195.320 ;
        RECT -26.380 194.340 -24.650 194.510 ;
        RECT -29.245 192.750 -26.560 192.920 ;
        RECT -29.245 192.720 -28.565 192.750 ;
        RECT -31.385 191.770 -30.850 191.940 ;
        RECT -37.945 190.995 -36.540 191.165 ;
        RECT -41.780 189.935 -39.580 190.105 ;
        RECT -41.780 189.930 -41.065 189.935 ;
        RECT -41.780 189.050 -41.610 189.930 ;
        RECT -38.845 189.725 -38.575 190.400 ;
        RECT -37.945 190.185 -37.760 190.995 ;
        RECT -37.945 190.015 -36.540 190.185 ;
        RECT -37.945 189.555 -37.760 190.015 ;
        RECT -39.260 189.540 -37.760 189.555 ;
        RECT -41.120 189.370 -37.760 189.540 ;
        RECT -41.780 188.880 -39.580 189.050 ;
        RECT -39.260 188.560 -39.090 189.370 ;
        RECT -55.320 188.390 -53.290 188.560 ;
        RECT -41.120 188.390 -39.090 188.560 ;
        RECT -38.820 187.345 -38.635 189.370 ;
        RECT -55.825 186.670 -55.555 187.345 ;
        RECT -38.855 186.670 -38.585 187.345 ;
        RECT -57.870 186.325 -53.290 186.495 ;
        RECT -41.120 186.325 -36.540 186.495 ;
        RECT -54.870 185.570 -54.580 186.325 ;
        RECT -52.305 185.570 -52.075 185.575 ;
        RECT -54.870 185.245 -52.075 185.570 ;
        RECT -63.115 184.850 -55.280 185.050 ;
        RECT -52.305 184.895 -52.075 185.245 ;
        RECT -42.335 185.570 -42.105 185.575 ;
        RECT -39.830 185.570 -39.540 186.325 ;
        RECT -42.335 185.245 -39.540 185.570 ;
        RECT -42.335 184.895 -42.105 185.245 ;
        RECT -65.845 178.395 -65.165 178.425 ;
        RECT -65.850 178.390 -65.165 178.395 ;
        RECT -67.850 178.220 -65.165 178.390 ;
        RECT -65.845 178.195 -65.165 178.220 ;
        RECT -63.605 177.935 -63.375 178.615 ;
        RECT -63.115 177.710 -62.945 184.850 ;
        RECT -63.905 177.540 -62.945 177.710 ;
        RECT -62.775 184.555 -55.770 184.655 ;
        RECT -62.775 184.475 -55.760 184.555 ;
        RECT -67.470 175.700 -67.200 176.395 ;
        RECT -68.115 175.455 -65.945 175.480 ;
        RECT -69.070 175.285 -65.000 175.455 ;
        RECT -68.115 175.265 -65.945 175.285 ;
        RECT -67.130 174.765 -66.900 175.265 ;
        RECT -68.105 173.910 -65.955 173.930 ;
        RECT -69.070 173.740 -65.000 173.910 ;
        RECT -68.105 173.715 -65.955 173.740 ;
        RECT -67.500 172.625 -67.230 173.320 ;
        RECT -66.410 173.235 -66.180 173.715 ;
        RECT -66.625 172.680 -65.000 172.850 ;
        RECT -69.070 172.190 -67.315 172.360 ;
        RECT -69.070 171.210 -67.685 171.380 ;
        RECT -67.855 170.480 -67.685 171.210 ;
        RECT -69.760 170.310 -67.685 170.480 ;
        RECT -69.760 167.990 -69.590 170.310 ;
        RECT -67.485 170.130 -67.315 172.190 ;
        RECT -66.625 171.380 -66.455 172.680 ;
        RECT -65.085 172.360 -64.635 172.370 ;
        RECT -66.040 172.190 -64.635 172.360 ;
        RECT -67.130 170.580 -66.860 171.275 ;
        RECT -66.625 171.210 -65.000 171.380 ;
        RECT -66.625 170.215 -66.455 171.210 ;
        RECT -69.415 169.960 -67.315 170.130 ;
        RECT -67.105 170.045 -66.455 170.215 ;
        RECT -66.190 170.720 -65.000 170.890 ;
        RECT -69.415 169.570 -69.245 169.960 ;
        RECT -67.105 169.655 -66.935 170.045 ;
        RECT -69.415 169.400 -68.030 169.570 ;
        RECT -67.850 169.485 -66.935 169.655 ;
        RECT -66.190 169.570 -65.995 170.720 ;
        RECT -69.415 168.590 -69.245 169.400 ;
        RECT -67.850 169.080 -67.680 169.485 ;
        RECT -66.190 169.400 -65.000 169.570 ;
        RECT -66.190 169.390 -65.995 169.400 ;
        RECT -69.070 168.910 -67.680 169.080 ;
        RECT -69.415 168.420 -68.030 168.590 ;
        RECT -69.760 167.820 -68.030 167.990 ;
        RECT -69.760 167.010 -69.590 167.820 ;
        RECT -67.850 167.500 -67.680 168.910 ;
        RECT -69.070 167.330 -67.680 167.500 ;
        RECT -69.760 166.840 -68.030 167.010 ;
        RECT -67.850 166.310 -67.680 167.330 ;
        RECT -67.280 166.835 -67.010 167.530 ;
        RECT -64.815 167.500 -64.635 172.190 ;
        RECT -63.905 167.700 -63.735 177.540 ;
        RECT -62.775 177.230 -62.595 184.475 ;
        RECT -55.960 184.295 -55.760 184.475 ;
        RECT -55.990 183.620 -55.720 184.295 ;
        RECT -55.480 184.030 -55.280 184.850 ;
        RECT -39.130 184.850 -31.295 185.050 ;
        RECT -39.130 184.030 -38.930 184.850 ;
        RECT -38.640 184.555 -31.635 184.655 ;
        RECT -38.650 184.475 -31.635 184.555 ;
        RECT -38.650 184.295 -38.450 184.475 ;
        RECT -55.480 184.025 -55.270 184.030 ;
        RECT -55.470 183.675 -55.270 184.025 ;
        RECT -39.140 184.025 -38.930 184.030 ;
        RECT -55.060 183.700 -53.520 183.870 ;
        RECT -40.890 183.700 -39.350 183.870 ;
        RECT -39.140 183.675 -38.940 184.025 ;
        RECT -57.745 183.210 -55.835 183.380 ;
        RECT -56.025 182.400 -55.835 183.210 ;
        RECT -57.745 182.230 -55.835 182.400 ;
        RECT -56.025 181.535 -55.835 182.230 ;
        RECT -55.470 181.970 -55.275 183.675 ;
        RECT -55.060 182.720 -53.520 182.890 ;
        RECT -40.890 182.720 -39.350 182.890 ;
        RECT -55.060 182.230 -53.520 182.400 ;
        RECT -40.890 182.230 -39.350 182.400 ;
        RECT -39.135 181.970 -38.940 183.675 ;
        RECT -38.690 183.620 -38.420 184.295 ;
        RECT -38.575 183.210 -36.665 183.380 ;
        RECT -38.575 182.400 -38.385 183.210 ;
        RECT -38.575 182.230 -36.665 182.400 ;
        RECT -55.600 181.600 -55.245 181.970 ;
        RECT -55.060 181.740 -53.520 181.910 ;
        RECT -40.890 181.740 -39.350 181.910 ;
        RECT -39.165 181.600 -38.810 181.970 ;
        RECT -56.835 181.425 -55.835 181.535 ;
        RECT -56.975 181.285 -55.835 181.425 ;
        RECT -38.575 181.535 -38.385 182.230 ;
        RECT -38.575 181.425 -37.575 181.535 ;
        RECT -38.575 181.285 -37.435 181.425 ;
        RECT -56.975 181.230 -55.875 181.285 ;
        RECT -38.535 181.230 -37.435 181.285 ;
        RECT -56.975 180.925 -56.770 181.230 ;
        RECT -37.640 180.925 -37.435 181.230 ;
        RECT -57.040 180.560 -56.740 180.925 ;
        RECT -37.670 180.560 -37.370 180.925 ;
        RECT -57.750 180.165 -57.210 180.335 ;
        RECT -37.200 180.165 -36.660 180.335 ;
        RECT -56.595 179.675 -56.055 179.845 ;
        RECT -38.355 179.675 -37.815 179.845 ;
        RECT -57.750 179.185 -57.210 179.355 ;
        RECT -37.200 179.185 -36.660 179.355 ;
        RECT -56.595 178.695 -56.055 178.865 ;
        RECT -38.355 178.695 -37.815 178.865 ;
        RECT -57.750 178.205 -56.540 178.375 ;
        RECT -56.890 177.735 -56.540 178.205 ;
        RECT -37.870 178.205 -36.660 178.375 ;
        RECT -37.870 177.735 -37.520 178.205 ;
        RECT -56.890 177.385 -52.635 177.735 ;
        RECT -63.515 177.050 -62.595 177.230 ;
        RECT -52.865 177.055 -52.635 177.385 ;
        RECT -41.775 177.385 -37.520 177.735 ;
        RECT -41.775 177.055 -41.545 177.385 ;
        RECT -31.815 177.230 -31.635 184.475 ;
        RECT -31.465 177.710 -31.295 184.850 ;
        RECT -31.020 178.615 -30.850 191.770 ;
        RECT -27.210 188.200 -26.940 188.895 ;
        RECT -28.465 187.955 -26.295 187.980 ;
        RECT -29.410 187.785 -25.340 187.955 ;
        RECT -28.465 187.765 -26.295 187.785 ;
        RECT -27.510 187.265 -27.280 187.765 ;
        RECT -28.455 186.410 -26.305 186.430 ;
        RECT -29.410 186.240 -25.340 186.410 ;
        RECT -28.455 186.215 -26.305 186.240 ;
        RECT -28.230 185.735 -28.000 186.215 ;
        RECT -29.410 185.180 -27.785 185.350 ;
        RECT -29.775 184.860 -29.325 184.870 ;
        RECT -29.775 184.690 -28.370 184.860 ;
        RECT -29.775 180.000 -29.595 184.690 ;
        RECT -27.955 183.880 -27.785 185.180 ;
        RECT -27.180 185.125 -26.910 185.820 ;
        RECT -29.410 183.710 -27.785 183.880 ;
        RECT -27.095 184.690 -25.340 184.860 ;
        RECT -29.410 183.220 -28.220 183.390 ;
        RECT -28.415 182.070 -28.220 183.220 ;
        RECT -27.955 182.715 -27.785 183.710 ;
        RECT -27.550 183.080 -27.280 183.775 ;
        RECT -27.955 182.545 -27.305 182.715 ;
        RECT -29.410 181.900 -28.220 182.070 ;
        RECT -27.475 182.155 -27.305 182.545 ;
        RECT -27.095 182.630 -26.925 184.690 ;
        RECT -26.725 183.710 -25.340 183.880 ;
        RECT -26.725 182.980 -26.555 183.710 ;
        RECT -26.725 182.810 -24.650 182.980 ;
        RECT -27.095 182.460 -24.995 182.630 ;
        RECT -27.475 181.985 -26.560 182.155 ;
        RECT -25.165 182.070 -24.995 182.460 ;
        RECT -28.415 181.890 -28.220 181.900 ;
        RECT -26.730 181.580 -26.560 181.985 ;
        RECT -26.380 181.900 -24.995 182.070 ;
        RECT -26.730 181.410 -25.340 181.580 ;
        RECT -29.775 179.830 -28.370 180.000 ;
        RECT -27.400 179.335 -27.130 180.030 ;
        RECT -26.730 180.000 -26.560 181.410 ;
        RECT -25.165 181.090 -24.995 181.900 ;
        RECT -26.380 180.920 -24.995 181.090 ;
        RECT -24.820 180.490 -24.650 182.810 ;
        RECT -26.380 180.320 -24.650 180.490 ;
        RECT -26.730 179.830 -25.340 180.000 ;
        RECT -31.035 177.935 -30.805 178.615 ;
        RECT -29.245 178.395 -28.565 178.425 ;
        RECT -29.245 178.390 -28.560 178.395 ;
        RECT -26.730 178.390 -26.560 179.830 ;
        RECT -24.820 179.510 -24.650 180.320 ;
        RECT -26.380 179.340 -24.650 179.510 ;
        RECT -29.245 178.220 -26.560 178.390 ;
        RECT -29.245 178.195 -28.565 178.220 ;
        RECT -31.465 177.540 -30.505 177.710 ;
        RECT -31.815 177.050 -30.895 177.230 ;
        RECT -66.040 167.330 -64.635 167.500 ;
        RECT -63.920 167.020 -63.690 167.700 ;
        RECT -63.905 166.855 -63.735 167.020 ;
        RECT -65.845 166.310 -65.165 166.340 ;
        RECT -67.855 166.140 -65.165 166.310 ;
        RECT -65.845 166.110 -65.165 166.140 ;
        RECT -67.470 163.200 -67.200 163.895 ;
        RECT -68.115 162.955 -65.945 162.980 ;
        RECT -69.070 162.785 -65.000 162.955 ;
        RECT -68.115 162.765 -65.945 162.785 ;
        RECT -67.130 162.265 -66.900 162.765 ;
        RECT -68.105 161.410 -65.955 161.430 ;
        RECT -69.070 161.240 -65.000 161.410 ;
        RECT -68.105 161.215 -65.955 161.240 ;
        RECT -67.500 160.125 -67.230 160.820 ;
        RECT -66.410 160.735 -66.180 161.215 ;
        RECT -66.625 160.180 -65.000 160.350 ;
        RECT -69.070 159.690 -67.315 159.860 ;
        RECT -69.070 158.710 -67.685 158.880 ;
        RECT -67.855 157.980 -67.685 158.710 ;
        RECT -69.760 157.810 -67.685 157.980 ;
        RECT -69.760 155.490 -69.590 157.810 ;
        RECT -67.485 157.630 -67.315 159.690 ;
        RECT -66.625 158.880 -66.455 160.180 ;
        RECT -65.085 159.860 -64.635 159.870 ;
        RECT -66.040 159.690 -64.635 159.860 ;
        RECT -67.130 158.080 -66.860 158.775 ;
        RECT -66.625 158.710 -65.000 158.880 ;
        RECT -66.625 157.715 -66.455 158.710 ;
        RECT -69.415 157.460 -67.315 157.630 ;
        RECT -67.105 157.545 -66.455 157.715 ;
        RECT -66.190 158.220 -65.000 158.390 ;
        RECT -69.415 157.070 -69.245 157.460 ;
        RECT -67.105 157.155 -66.935 157.545 ;
        RECT -69.415 156.900 -68.030 157.070 ;
        RECT -67.850 156.985 -66.935 157.155 ;
        RECT -66.190 157.070 -65.995 158.220 ;
        RECT -69.415 156.090 -69.245 156.900 ;
        RECT -67.850 156.580 -67.680 156.985 ;
        RECT -66.190 156.900 -65.000 157.070 ;
        RECT -66.190 156.890 -65.995 156.900 ;
        RECT -69.070 156.410 -67.680 156.580 ;
        RECT -69.415 155.920 -68.030 156.090 ;
        RECT -69.760 155.320 -68.030 155.490 ;
        RECT -69.760 154.510 -69.590 155.320 ;
        RECT -67.850 155.000 -67.680 156.410 ;
        RECT -69.070 154.830 -67.680 155.000 ;
        RECT -69.760 154.340 -68.030 154.510 ;
        RECT -67.850 153.910 -67.680 154.830 ;
        RECT -67.280 154.335 -67.010 155.030 ;
        RECT -64.815 155.000 -64.635 159.690 ;
        RECT -63.515 155.215 -63.335 177.050 ;
        RECT -60.400 176.710 -55.290 176.910 ;
        RECT -60.400 176.230 -60.170 176.710 ;
        RECT -55.960 176.485 -55.780 176.530 ;
        RECT -59.980 176.420 -55.780 176.485 ;
        RECT -59.980 176.305 -55.760 176.420 ;
        RECT -59.980 175.710 -59.750 176.305 ;
        RECT -56.000 176.270 -55.760 176.305 ;
        RECT -56.000 175.595 -55.730 176.270 ;
        RECT -55.490 176.005 -55.290 176.710 ;
        RECT -39.120 176.710 -34.010 176.910 ;
        RECT -39.120 176.005 -38.920 176.710 ;
        RECT -38.630 176.485 -38.450 176.530 ;
        RECT -38.630 176.420 -34.430 176.485 ;
        RECT -38.650 176.305 -34.430 176.420 ;
        RECT -38.650 176.270 -38.410 176.305 ;
        RECT -55.490 176.000 -55.280 176.005 ;
        RECT -55.480 175.650 -55.280 176.000 ;
        RECT -39.130 176.000 -38.920 176.005 ;
        RECT -55.070 175.675 -53.530 175.845 ;
        RECT -40.880 175.675 -39.340 175.845 ;
        RECT -39.130 175.650 -38.930 176.000 ;
        RECT -57.755 175.185 -55.845 175.355 ;
        RECT -56.035 174.375 -55.845 175.185 ;
        RECT -57.755 174.205 -55.845 174.375 ;
        RECT -56.035 173.510 -55.845 174.205 ;
        RECT -55.480 173.945 -55.285 175.650 ;
        RECT -55.070 174.695 -53.530 174.865 ;
        RECT -40.880 174.695 -39.340 174.865 ;
        RECT -55.070 174.205 -53.530 174.375 ;
        RECT -40.880 174.205 -39.340 174.375 ;
        RECT -39.125 173.945 -38.930 175.650 ;
        RECT -38.680 175.595 -38.410 176.270 ;
        RECT -34.660 175.710 -34.430 176.305 ;
        RECT -34.240 176.230 -34.010 176.710 ;
        RECT -38.565 175.185 -36.655 175.355 ;
        RECT -38.565 174.375 -38.375 175.185 ;
        RECT -38.565 174.205 -36.655 174.375 ;
        RECT -55.610 173.575 -55.255 173.945 ;
        RECT -55.070 173.715 -53.530 173.885 ;
        RECT -40.880 173.715 -39.340 173.885 ;
        RECT -39.155 173.575 -38.800 173.945 ;
        RECT -56.845 173.400 -55.845 173.510 ;
        RECT -56.985 173.260 -55.845 173.400 ;
        RECT -38.565 173.510 -38.375 174.205 ;
        RECT -38.565 173.400 -37.565 173.510 ;
        RECT -38.565 173.260 -37.425 173.400 ;
        RECT -56.985 173.205 -55.885 173.260 ;
        RECT -38.525 173.205 -37.425 173.260 ;
        RECT -56.985 172.900 -56.780 173.205 ;
        RECT -37.630 172.900 -37.425 173.205 ;
        RECT -57.050 172.535 -56.750 172.900 ;
        RECT -37.660 172.535 -37.360 172.900 ;
        RECT -57.760 172.140 -57.220 172.310 ;
        RECT -37.190 172.140 -36.650 172.310 ;
        RECT -56.605 171.650 -56.065 171.820 ;
        RECT -38.345 171.650 -37.805 171.820 ;
        RECT -57.760 171.160 -57.220 171.330 ;
        RECT -37.190 171.160 -36.650 171.330 ;
        RECT -56.605 170.670 -56.065 170.840 ;
        RECT -38.345 170.670 -37.805 170.840 ;
        RECT -57.760 170.180 -56.550 170.350 ;
        RECT -56.900 169.695 -56.550 170.180 ;
        RECT -37.860 170.180 -36.650 170.350 ;
        RECT -37.860 169.695 -37.510 170.180 ;
        RECT -56.900 169.525 -55.555 169.695 ;
        RECT -56.900 169.495 -56.550 169.525 ;
        RECT -56.140 168.670 -55.910 169.350 ;
        RECT -57.010 168.265 -56.320 168.495 ;
        RECT -56.590 167.535 -56.320 168.265 ;
        RECT -57.825 167.165 -56.420 167.335 ;
        RECT -56.605 166.355 -56.420 167.165 ;
        RECT -56.135 166.530 -55.945 168.670 ;
        RECT -57.825 166.185 -56.420 166.355 ;
        RECT -56.605 165.375 -56.420 166.185 ;
        RECT -56.180 165.855 -55.910 166.530 ;
        RECT -55.725 165.590 -55.555 169.525 ;
        RECT -38.855 169.525 -37.510 169.695 ;
        RECT -55.275 167.655 -53.250 167.825 ;
        RECT -41.160 167.655 -39.135 167.825 ;
        RECT -55.275 166.845 -55.105 167.655 ;
        RECT -39.305 166.845 -39.135 167.655 ;
        RECT -55.275 166.675 -53.250 166.845 ;
        RECT -41.160 166.675 -39.135 166.845 ;
        RECT -55.275 165.785 -55.100 166.675 ;
        RECT -54.785 166.105 -52.585 166.275 ;
        RECT -53.290 166.100 -52.585 166.105 ;
        RECT -55.275 165.615 -53.245 165.785 ;
        RECT -55.275 165.610 -54.785 165.615 ;
        RECT -57.825 165.205 -56.420 165.375 ;
        RECT -56.605 164.745 -56.420 165.205 ;
        RECT -55.790 164.915 -55.520 165.590 ;
        RECT -52.770 165.295 -52.585 166.100 ;
        RECT -54.785 165.125 -52.585 165.295 ;
        RECT -53.300 165.120 -52.585 165.125 ;
        RECT -56.605 164.730 -55.105 164.745 ;
        RECT -56.605 164.560 -53.245 164.730 ;
        RECT -55.730 162.535 -55.545 164.560 ;
        RECT -55.275 163.750 -55.105 164.560 ;
        RECT -52.755 164.240 -52.585 165.120 ;
        RECT -54.785 164.070 -52.585 164.240 ;
        RECT -41.825 166.105 -39.625 166.275 ;
        RECT -41.825 166.100 -41.120 166.105 ;
        RECT -41.825 165.295 -41.640 166.100 ;
        RECT -39.310 165.785 -39.135 166.675 ;
        RECT -41.165 165.615 -39.135 165.785 ;
        RECT -39.625 165.610 -39.135 165.615 ;
        RECT -38.855 165.590 -38.685 169.525 ;
        RECT -37.860 169.495 -37.510 169.525 ;
        RECT -38.500 168.670 -38.270 169.350 ;
        RECT -38.465 166.530 -38.275 168.670 ;
        RECT -38.090 168.265 -37.400 168.495 ;
        RECT -38.090 167.535 -37.820 168.265 ;
        RECT -37.990 167.165 -36.585 167.335 ;
        RECT -38.500 165.855 -38.230 166.530 ;
        RECT -37.990 166.355 -37.805 167.165 ;
        RECT -37.990 166.185 -36.585 166.355 ;
        RECT -41.825 165.125 -39.625 165.295 ;
        RECT -41.825 165.120 -41.110 165.125 ;
        RECT -41.825 164.240 -41.655 165.120 ;
        RECT -38.890 164.915 -38.620 165.590 ;
        RECT -37.990 165.375 -37.805 166.185 ;
        RECT -37.990 165.205 -36.585 165.375 ;
        RECT -37.990 164.745 -37.805 165.205 ;
        RECT -39.305 164.730 -37.805 164.745 ;
        RECT -41.165 164.560 -37.805 164.730 ;
        RECT -41.825 164.070 -39.625 164.240 ;
        RECT -39.305 163.750 -39.135 164.560 ;
        RECT -55.275 163.580 -53.245 163.750 ;
        RECT -41.165 163.580 -39.135 163.750 ;
        RECT -38.865 162.535 -38.680 164.560 ;
        RECT -55.780 161.860 -55.510 162.535 ;
        RECT -38.900 161.860 -38.630 162.535 ;
        RECT -57.825 161.515 -53.245 161.685 ;
        RECT -41.165 161.515 -36.585 161.685 ;
        RECT -55.775 160.760 -55.510 161.515 ;
        RECT -38.900 160.760 -38.635 161.515 ;
        RECT -57.890 158.995 -55.930 159.025 ;
        RECT -38.480 158.995 -36.520 159.025 ;
        RECT -57.910 158.825 -55.470 158.995 ;
        RECT -38.940 158.825 -36.500 158.995 ;
        RECT -57.890 158.795 -55.930 158.825 ;
        RECT -38.480 158.795 -36.520 158.825 ;
        RECT -56.625 158.045 -56.395 158.795 ;
        RECT -38.015 158.045 -37.785 158.795 ;
        RECT -56.950 158.015 -55.930 158.045 ;
        RECT -38.480 158.015 -37.460 158.045 ;
        RECT -57.910 157.845 -55.470 158.015 ;
        RECT -38.940 157.845 -36.500 158.015 ;
        RECT -56.950 157.815 -55.930 157.845 ;
        RECT -38.480 157.815 -37.460 157.845 ;
        RECT -56.625 157.065 -56.395 157.815 ;
        RECT -56.950 157.035 -55.930 157.065 ;
        RECT -57.910 156.865 -55.470 157.035 ;
        RECT -40.450 156.990 -40.150 157.650 ;
        RECT -38.015 157.065 -37.785 157.815 ;
        RECT -38.480 157.035 -37.460 157.065 ;
        RECT -56.950 156.835 -55.930 156.865 ;
        RECT -56.585 156.685 -56.235 156.835 ;
        RECT -56.475 156.395 -56.265 156.685 ;
        RECT -56.495 156.095 -55.835 156.395 ;
        RECT -56.475 155.810 -56.265 156.095 ;
        RECT -54.695 155.940 -54.395 156.600 ;
        RECT -57.800 155.405 -56.980 155.690 ;
        RECT -56.495 155.635 -56.205 155.810 ;
        RECT -66.040 154.830 -64.635 155.000 ;
        RECT -63.985 154.970 -63.335 155.215 ;
        RECT -63.985 154.535 -63.755 154.970 ;
        RECT -56.550 154.795 -56.180 155.635 ;
        RECT -57.890 154.585 -55.930 154.615 ;
        RECT -57.910 154.415 -55.470 154.585 ;
        RECT -57.890 154.385 -55.930 154.415 ;
        RECT -65.845 153.910 -65.165 153.940 ;
        RECT -67.850 153.740 -65.165 153.910 ;
        RECT -65.845 153.710 -65.165 153.740 ;
        RECT -56.625 153.635 -56.395 154.385 ;
        RECT -56.950 153.605 -55.930 153.635 ;
        RECT -57.910 153.435 -55.470 153.605 ;
        RECT -56.950 153.405 -55.930 153.435 ;
        RECT -56.625 152.655 -56.395 153.405 ;
        RECT -56.950 152.625 -55.930 152.655 ;
        RECT -57.910 152.455 -55.470 152.625 ;
        RECT -56.950 152.425 -55.930 152.455 ;
        RECT -56.585 152.150 -56.235 152.425 ;
        RECT -57.545 151.785 -56.235 152.150 ;
        RECT -57.545 151.780 -56.705 151.785 ;
        RECT -58.175 151.530 -57.780 151.535 ;
        RECT -57.410 151.530 -55.630 151.560 ;
        RECT -55.280 151.530 -54.820 151.555 ;
        RECT -67.470 150.700 -67.200 151.395 ;
        RECT -58.175 151.360 -54.820 151.530 ;
        RECT -58.175 151.355 -57.780 151.360 ;
        RECT -58.175 150.555 -58.005 151.355 ;
        RECT -57.410 151.325 -55.630 151.360 ;
        RECT -55.280 151.335 -54.820 151.360 ;
        RECT -57.375 151.040 -56.945 151.045 ;
        RECT -57.835 150.870 -56.945 151.040 ;
        RECT -57.375 150.865 -56.945 150.870 ;
        RECT -58.175 150.550 -57.730 150.555 ;
        RECT -68.115 150.455 -65.945 150.480 ;
        RECT -69.070 150.285 -65.000 150.455 ;
        RECT -58.175 150.380 -57.295 150.550 ;
        RECT -58.175 150.345 -57.730 150.380 ;
        RECT -68.115 150.265 -65.945 150.285 ;
        RECT -67.130 149.765 -66.900 150.265 ;
        RECT -58.175 149.585 -58.005 150.345 ;
        RECT -57.835 150.055 -57.295 150.060 ;
        RECT -57.115 150.055 -56.945 150.865 ;
        RECT -56.675 150.700 -56.305 151.325 ;
        RECT -56.110 151.040 -55.735 151.060 ;
        RECT -56.110 150.870 -55.220 151.040 ;
        RECT -56.110 150.855 -55.735 150.870 ;
        RECT -57.835 149.890 -56.945 150.055 ;
        RECT -57.385 149.875 -56.945 149.890 ;
        RECT -58.175 149.570 -57.725 149.585 ;
        RECT -58.175 149.400 -57.295 149.570 ;
        RECT -58.175 149.375 -57.725 149.400 ;
        RECT -68.105 148.910 -65.955 148.930 ;
        RECT -69.070 148.740 -65.000 148.910 ;
        RECT -68.105 148.715 -65.955 148.740 ;
        RECT -67.500 147.625 -67.230 148.320 ;
        RECT -66.410 148.235 -66.180 148.715 ;
        RECT -58.175 148.605 -58.005 149.375 ;
        RECT -57.115 149.085 -56.945 149.875 ;
        RECT -57.385 149.080 -56.945 149.085 ;
        RECT -57.835 148.910 -56.945 149.080 ;
        RECT -57.385 148.905 -56.945 148.910 ;
        RECT -57.115 148.780 -56.945 148.905 ;
        RECT -56.110 150.070 -55.940 150.855 ;
        RECT -54.990 150.575 -54.820 151.335 ;
        RECT -55.335 150.550 -54.820 150.575 ;
        RECT -55.760 150.380 -54.820 150.550 ;
        RECT -55.335 150.355 -54.820 150.380 ;
        RECT -56.110 150.060 -55.695 150.070 ;
        RECT -56.110 149.890 -55.220 150.060 ;
        RECT -56.110 149.865 -55.695 149.890 ;
        RECT -56.110 149.100 -55.940 149.865 ;
        RECT -54.990 149.595 -54.820 150.355 ;
        RECT -55.335 149.570 -54.820 149.595 ;
        RECT -55.760 149.400 -54.820 149.570 ;
        RECT -55.335 149.375 -54.820 149.400 ;
        RECT -56.110 149.080 -55.695 149.100 ;
        RECT -56.110 148.910 -55.220 149.080 ;
        RECT -56.110 148.895 -55.695 148.910 ;
        RECT -56.110 148.780 -55.940 148.895 ;
        RECT -58.175 148.590 -57.750 148.605 ;
        RECT -58.175 148.420 -57.295 148.590 ;
        RECT -58.175 148.395 -57.750 148.420 ;
        RECT -57.115 148.115 -55.940 148.780 ;
        RECT -54.990 148.610 -54.820 149.375 ;
        RECT -55.280 148.590 -54.820 148.610 ;
        RECT -55.760 148.420 -54.820 148.590 ;
        RECT -55.280 148.390 -54.820 148.420 ;
        RECT -55.740 148.115 -55.080 148.145 ;
        RECT -57.335 148.100 -55.080 148.115 ;
        RECT -57.835 147.930 -55.080 148.100 ;
        RECT -57.335 147.915 -55.080 147.930 ;
        RECT -57.335 147.910 -55.690 147.915 ;
        RECT -57.335 147.905 -55.905 147.910 ;
        RECT -66.625 147.680 -65.000 147.850 ;
        RECT -69.070 147.190 -67.315 147.360 ;
        RECT -69.070 146.210 -67.685 146.380 ;
        RECT -67.855 145.480 -67.685 146.210 ;
        RECT -69.760 145.310 -67.685 145.480 ;
        RECT -69.760 142.990 -69.590 145.310 ;
        RECT -67.485 145.130 -67.315 147.190 ;
        RECT -66.625 146.380 -66.455 147.680 ;
        RECT -65.085 147.360 -64.635 147.370 ;
        RECT -66.040 147.190 -64.635 147.360 ;
        RECT -67.130 145.580 -66.860 146.275 ;
        RECT -66.625 146.210 -65.000 146.380 ;
        RECT -66.625 145.215 -66.455 146.210 ;
        RECT -69.415 144.960 -67.315 145.130 ;
        RECT -67.105 145.045 -66.455 145.215 ;
        RECT -66.190 145.720 -65.000 145.890 ;
        RECT -69.415 144.570 -69.245 144.960 ;
        RECT -67.105 144.655 -66.935 145.045 ;
        RECT -69.415 144.400 -68.030 144.570 ;
        RECT -67.850 144.485 -66.935 144.655 ;
        RECT -66.190 144.570 -65.995 145.720 ;
        RECT -69.415 143.590 -69.245 144.400 ;
        RECT -67.850 144.080 -67.680 144.485 ;
        RECT -66.190 144.400 -65.000 144.570 ;
        RECT -66.190 144.390 -65.995 144.400 ;
        RECT -69.070 143.910 -67.680 144.080 ;
        RECT -69.415 143.420 -68.030 143.590 ;
        RECT -69.760 142.820 -68.030 142.990 ;
        RECT -69.760 142.010 -69.590 142.820 ;
        RECT -67.850 142.500 -67.680 143.910 ;
        RECT -69.070 142.330 -67.680 142.500 ;
        RECT -69.760 141.840 -68.030 142.010 ;
        RECT -67.850 141.170 -67.680 142.330 ;
        RECT -67.280 141.835 -67.010 142.530 ;
        RECT -64.815 142.500 -64.635 147.190 ;
        RECT -56.505 146.920 -56.220 147.905 ;
        RECT -56.550 146.080 -56.180 146.920 ;
        RECT -57.890 145.870 -55.930 145.900 ;
        RECT -57.910 145.700 -55.470 145.870 ;
        RECT -57.890 145.670 -55.930 145.700 ;
        RECT -56.625 144.920 -56.395 145.670 ;
        RECT -56.950 144.890 -55.930 144.920 ;
        RECT -57.910 144.720 -55.470 144.890 ;
        RECT -56.950 144.690 -55.930 144.720 ;
        RECT -56.625 143.940 -56.395 144.690 ;
        RECT -56.950 143.910 -55.930 143.940 ;
        RECT -57.910 143.740 -55.470 143.910 ;
        RECT -56.950 143.710 -55.930 143.740 ;
        RECT -56.585 143.560 -56.235 143.710 ;
        RECT -56.515 143.310 -56.290 143.560 ;
        RECT -56.515 143.210 -55.715 143.310 ;
        RECT -66.040 142.330 -64.635 142.500 ;
        RECT -57.410 143.010 -55.715 143.210 ;
        RECT -57.410 142.985 -56.290 143.010 ;
        RECT -57.410 142.190 -57.185 142.985 ;
        RECT -57.800 141.905 -56.980 142.190 ;
        RECT -65.865 141.170 -65.185 141.200 ;
        RECT -67.850 141.000 -65.185 141.170 ;
        RECT -65.865 140.970 -65.185 141.000 ;
        RECT -62.335 141.185 -61.655 141.200 ;
        RECT -60.390 141.185 -60.160 141.665 ;
        RECT -62.335 140.985 -60.160 141.185 ;
        RECT -57.890 141.085 -55.930 141.115 ;
        RECT -62.335 140.970 -61.655 140.985 ;
        RECT -57.910 140.915 -55.470 141.085 ;
        RECT -57.890 140.885 -55.930 140.915 ;
        RECT -56.625 140.135 -56.395 140.885 ;
        RECT -56.950 140.105 -55.930 140.135 ;
        RECT -57.910 139.935 -55.470 140.105 ;
        RECT -56.950 139.905 -55.930 139.935 ;
        RECT -56.625 139.155 -56.395 139.905 ;
        RECT -56.950 139.125 -55.930 139.155 ;
        RECT -57.910 138.955 -55.470 139.125 ;
        RECT -56.950 138.925 -55.930 138.955 ;
        RECT -67.470 138.200 -67.200 138.895 ;
        RECT -56.585 138.650 -56.235 138.925 ;
        RECT -57.545 138.285 -56.235 138.650 ;
        RECT -57.545 138.280 -56.705 138.285 ;
        RECT -58.175 138.030 -57.780 138.035 ;
        RECT -57.410 138.030 -55.630 138.060 ;
        RECT -55.280 138.030 -54.820 138.055 ;
        RECT -68.115 137.955 -65.945 137.980 ;
        RECT -69.070 137.785 -65.000 137.955 ;
        RECT -58.175 137.860 -54.820 138.030 ;
        RECT -58.175 137.855 -57.780 137.860 ;
        RECT -68.115 137.765 -65.945 137.785 ;
        RECT -67.130 137.265 -66.900 137.765 ;
        RECT -58.175 137.055 -58.005 137.855 ;
        RECT -57.410 137.825 -55.630 137.860 ;
        RECT -55.280 137.835 -54.820 137.860 ;
        RECT -57.375 137.540 -56.945 137.545 ;
        RECT -57.835 137.370 -56.945 137.540 ;
        RECT -57.375 137.365 -56.945 137.370 ;
        RECT -58.175 137.050 -57.730 137.055 ;
        RECT -58.175 136.880 -57.295 137.050 ;
        RECT -58.175 136.845 -57.730 136.880 ;
        RECT -68.105 136.410 -65.955 136.430 ;
        RECT -69.070 136.240 -65.000 136.410 ;
        RECT -68.105 136.215 -65.955 136.240 ;
        RECT -67.500 135.125 -67.230 135.820 ;
        RECT -66.410 135.735 -66.180 136.215 ;
        RECT -58.175 136.085 -58.005 136.845 ;
        RECT -57.835 136.555 -57.295 136.560 ;
        RECT -57.115 136.555 -56.945 137.365 ;
        RECT -56.675 137.200 -56.305 137.825 ;
        RECT -56.110 137.540 -55.735 137.560 ;
        RECT -56.110 137.370 -55.220 137.540 ;
        RECT -56.110 137.355 -55.735 137.370 ;
        RECT -57.835 136.390 -56.945 136.555 ;
        RECT -57.385 136.375 -56.945 136.390 ;
        RECT -58.175 136.070 -57.725 136.085 ;
        RECT -58.175 135.900 -57.295 136.070 ;
        RECT -58.175 135.875 -57.725 135.900 ;
        RECT -66.625 135.180 -65.000 135.350 ;
        RECT -69.070 134.690 -67.315 134.860 ;
        RECT -69.070 133.710 -67.685 133.880 ;
        RECT -67.855 132.980 -67.685 133.710 ;
        RECT -69.760 132.810 -67.685 132.980 ;
        RECT -69.760 130.490 -69.590 132.810 ;
        RECT -67.485 132.630 -67.315 134.690 ;
        RECT -66.625 133.880 -66.455 135.180 ;
        RECT -58.175 135.105 -58.005 135.875 ;
        RECT -57.115 135.585 -56.945 136.375 ;
        RECT -57.385 135.580 -56.945 135.585 ;
        RECT -57.835 135.410 -56.945 135.580 ;
        RECT -57.385 135.405 -56.945 135.410 ;
        RECT -57.115 135.280 -56.945 135.405 ;
        RECT -56.110 136.570 -55.940 137.355 ;
        RECT -54.990 137.075 -54.820 137.835 ;
        RECT -55.335 137.050 -54.820 137.075 ;
        RECT -55.760 136.880 -54.820 137.050 ;
        RECT -55.335 136.855 -54.820 136.880 ;
        RECT -56.110 136.560 -55.695 136.570 ;
        RECT -56.110 136.390 -55.220 136.560 ;
        RECT -56.110 136.365 -55.695 136.390 ;
        RECT -56.110 135.600 -55.940 136.365 ;
        RECT -54.990 136.095 -54.820 136.855 ;
        RECT -55.335 136.070 -54.820 136.095 ;
        RECT -55.760 135.900 -54.820 136.070 ;
        RECT -55.335 135.875 -54.820 135.900 ;
        RECT -56.110 135.580 -55.695 135.600 ;
        RECT -56.110 135.410 -55.220 135.580 ;
        RECT -56.110 135.395 -55.695 135.410 ;
        RECT -56.110 135.280 -55.940 135.395 ;
        RECT -58.175 135.090 -57.750 135.105 ;
        RECT -58.175 134.920 -57.295 135.090 ;
        RECT -58.175 134.895 -57.750 134.920 ;
        RECT -65.085 134.860 -64.635 134.870 ;
        RECT -66.040 134.690 -64.635 134.860 ;
        RECT -67.130 133.080 -66.860 133.775 ;
        RECT -66.625 133.710 -65.000 133.880 ;
        RECT -66.625 132.715 -66.455 133.710 ;
        RECT -69.415 132.460 -67.315 132.630 ;
        RECT -67.105 132.545 -66.455 132.715 ;
        RECT -66.190 133.220 -65.000 133.390 ;
        RECT -69.415 132.070 -69.245 132.460 ;
        RECT -67.105 132.155 -66.935 132.545 ;
        RECT -69.415 131.900 -68.030 132.070 ;
        RECT -67.850 131.985 -66.935 132.155 ;
        RECT -66.190 132.070 -65.995 133.220 ;
        RECT -69.415 131.090 -69.245 131.900 ;
        RECT -67.850 131.580 -67.680 131.985 ;
        RECT -66.190 131.900 -65.000 132.070 ;
        RECT -66.190 131.890 -65.995 131.900 ;
        RECT -69.070 131.410 -67.680 131.580 ;
        RECT -69.415 130.920 -68.030 131.090 ;
        RECT -69.760 130.320 -68.030 130.490 ;
        RECT -69.760 129.510 -69.590 130.320 ;
        RECT -67.850 130.000 -67.680 131.410 ;
        RECT -69.070 129.830 -67.680 130.000 ;
        RECT -69.760 129.340 -68.030 129.510 ;
        RECT -67.850 128.955 -67.680 129.830 ;
        RECT -67.280 129.335 -67.010 130.030 ;
        RECT -64.815 130.000 -64.635 134.690 ;
        RECT -57.115 134.615 -55.940 135.280 ;
        RECT -54.990 135.110 -54.820 135.875 ;
        RECT -55.280 135.090 -54.820 135.110 ;
        RECT -55.760 134.920 -54.820 135.090 ;
        RECT -55.280 134.890 -54.820 134.920 ;
        RECT -57.335 134.600 -55.690 134.615 ;
        RECT -57.835 134.430 -55.220 134.600 ;
        RECT -57.335 134.410 -55.690 134.430 ;
        RECT -57.335 134.405 -55.905 134.410 ;
        RECT -56.520 133.420 -56.255 134.405 ;
        RECT -54.640 133.985 -54.445 155.940 ;
        RECT -52.090 155.095 -51.790 155.470 ;
        RECT -42.620 155.095 -42.320 155.470 ;
        RECT -52.285 155.090 -50.855 155.095 ;
        RECT -52.500 155.070 -50.855 155.090 ;
        RECT -43.555 155.090 -42.125 155.095 ;
        RECT -43.555 155.070 -41.910 155.090 ;
        RECT -52.970 154.900 -50.355 155.070 ;
        RECT -44.055 154.900 -41.440 155.070 ;
        RECT -52.500 154.885 -50.855 154.900 ;
        RECT -43.555 154.885 -41.910 154.900 ;
        RECT -53.370 154.580 -52.910 154.610 ;
        RECT -53.370 154.410 -52.430 154.580 ;
        RECT -53.370 154.390 -52.910 154.410 ;
        RECT -53.370 153.625 -53.200 154.390 ;
        RECT -52.250 154.220 -51.075 154.885 ;
        RECT -50.440 154.580 -50.015 154.605 ;
        RECT -50.895 154.410 -50.015 154.580 ;
        RECT -50.440 154.395 -50.015 154.410 ;
        RECT -52.250 154.105 -52.080 154.220 ;
        RECT -52.495 154.090 -52.080 154.105 ;
        RECT -52.970 153.920 -52.080 154.090 ;
        RECT -52.495 153.900 -52.080 153.920 ;
        RECT -53.370 153.600 -52.855 153.625 ;
        RECT -53.370 153.430 -52.430 153.600 ;
        RECT -53.370 153.405 -52.855 153.430 ;
        RECT -53.370 152.645 -53.200 153.405 ;
        RECT -52.250 153.135 -52.080 153.900 ;
        RECT -52.495 153.110 -52.080 153.135 ;
        RECT -52.970 152.940 -52.080 153.110 ;
        RECT -52.495 152.930 -52.080 152.940 ;
        RECT -53.370 152.620 -52.855 152.645 ;
        RECT -53.370 152.450 -52.430 152.620 ;
        RECT -53.370 152.425 -52.855 152.450 ;
        RECT -53.370 151.665 -53.200 152.425 ;
        RECT -52.250 152.145 -52.080 152.930 ;
        RECT -51.245 154.095 -51.075 154.220 ;
        RECT -51.245 154.090 -50.805 154.095 ;
        RECT -51.245 153.920 -50.355 154.090 ;
        RECT -51.245 153.915 -50.805 153.920 ;
        RECT -51.245 153.125 -51.075 153.915 ;
        RECT -50.185 153.625 -50.015 154.395 ;
        RECT -50.465 153.600 -50.015 153.625 ;
        RECT -50.895 153.430 -50.015 153.600 ;
        RECT -50.465 153.415 -50.015 153.430 ;
        RECT -51.245 153.110 -50.805 153.125 ;
        RECT -51.245 152.945 -50.355 153.110 ;
        RECT -52.455 152.130 -52.080 152.145 ;
        RECT -52.970 151.960 -52.080 152.130 ;
        RECT -52.455 151.940 -52.080 151.960 ;
        RECT -51.885 151.675 -51.515 152.300 ;
        RECT -51.245 152.135 -51.075 152.945 ;
        RECT -50.895 152.940 -50.355 152.945 ;
        RECT -50.185 152.655 -50.015 153.415 ;
        RECT -50.460 152.620 -50.015 152.655 ;
        RECT -50.895 152.450 -50.015 152.620 ;
        RECT -50.460 152.445 -50.015 152.450 ;
        RECT -51.245 152.130 -50.815 152.135 ;
        RECT -51.245 151.960 -50.355 152.130 ;
        RECT -51.245 151.955 -50.815 151.960 ;
        RECT -53.370 151.640 -52.910 151.665 ;
        RECT -52.560 151.640 -50.780 151.675 ;
        RECT -50.185 151.645 -50.015 152.445 ;
        RECT -50.410 151.640 -50.015 151.645 ;
        RECT -53.370 151.470 -50.015 151.640 ;
        RECT -53.370 151.445 -52.910 151.470 ;
        RECT -52.560 151.440 -50.780 151.470 ;
        RECT -50.410 151.465 -50.015 151.470 ;
        RECT -44.395 154.580 -43.970 154.605 ;
        RECT -44.395 154.410 -43.515 154.580 ;
        RECT -44.395 154.395 -43.970 154.410 ;
        RECT -44.395 153.625 -44.225 154.395 ;
        RECT -43.335 154.220 -42.160 154.885 ;
        RECT -41.500 154.580 -41.040 154.610 ;
        RECT -41.980 154.410 -41.040 154.580 ;
        RECT -41.500 154.390 -41.040 154.410 ;
        RECT -43.335 154.095 -43.165 154.220 ;
        RECT -43.605 154.090 -43.165 154.095 ;
        RECT -44.055 153.920 -43.165 154.090 ;
        RECT -43.605 153.915 -43.165 153.920 ;
        RECT -44.395 153.600 -43.945 153.625 ;
        RECT -44.395 153.430 -43.515 153.600 ;
        RECT -44.395 153.415 -43.945 153.430 ;
        RECT -44.395 152.655 -44.225 153.415 ;
        RECT -43.335 153.125 -43.165 153.915 ;
        RECT -43.605 153.110 -43.165 153.125 ;
        RECT -44.055 152.945 -43.165 153.110 ;
        RECT -44.055 152.940 -43.515 152.945 ;
        RECT -44.395 152.620 -43.950 152.655 ;
        RECT -44.395 152.450 -43.515 152.620 ;
        RECT -44.395 152.445 -43.950 152.450 ;
        RECT -44.395 151.645 -44.225 152.445 ;
        RECT -43.335 152.135 -43.165 152.945 ;
        RECT -42.330 154.105 -42.160 154.220 ;
        RECT -42.330 154.090 -41.915 154.105 ;
        RECT -42.330 153.920 -41.440 154.090 ;
        RECT -42.330 153.900 -41.915 153.920 ;
        RECT -42.330 153.135 -42.160 153.900 ;
        RECT -41.210 153.625 -41.040 154.390 ;
        RECT -41.555 153.600 -41.040 153.625 ;
        RECT -41.980 153.430 -41.040 153.600 ;
        RECT -41.555 153.405 -41.040 153.430 ;
        RECT -42.330 153.110 -41.915 153.135 ;
        RECT -42.330 152.940 -41.440 153.110 ;
        RECT -42.330 152.930 -41.915 152.940 ;
        RECT -43.595 152.130 -43.165 152.135 ;
        RECT -44.055 151.960 -43.165 152.130 ;
        RECT -43.595 151.955 -43.165 151.960 ;
        RECT -42.895 151.675 -42.525 152.300 ;
        RECT -42.330 152.145 -42.160 152.930 ;
        RECT -41.210 152.645 -41.040 153.405 ;
        RECT -41.555 152.620 -41.040 152.645 ;
        RECT -41.980 152.450 -41.040 152.620 ;
        RECT -41.555 152.425 -41.040 152.450 ;
        RECT -42.330 152.130 -41.955 152.145 ;
        RECT -42.330 151.960 -41.440 152.130 ;
        RECT -42.330 151.940 -41.955 151.960 ;
        RECT -44.395 151.640 -44.000 151.645 ;
        RECT -43.630 151.640 -41.850 151.675 ;
        RECT -41.210 151.665 -41.040 152.425 ;
        RECT -41.500 151.640 -41.040 151.665 ;
        RECT -44.395 151.470 -41.040 151.640 ;
        RECT -44.395 151.465 -44.000 151.470 ;
        RECT -43.630 151.440 -41.850 151.470 ;
        RECT -41.500 151.445 -41.040 151.470 ;
        RECT -51.485 151.215 -50.645 151.220 ;
        RECT -51.955 150.850 -50.645 151.215 ;
        RECT -43.765 151.215 -42.925 151.220 ;
        RECT -43.765 150.850 -42.455 151.215 ;
        RECT -51.955 150.575 -51.605 150.850 ;
        RECT -42.805 150.575 -42.455 150.850 ;
        RECT -52.260 150.545 -51.240 150.575 ;
        RECT -43.170 150.545 -42.150 150.575 ;
        RECT -52.720 150.375 -50.280 150.545 ;
        RECT -44.130 150.375 -41.690 150.545 ;
        RECT -52.260 150.345 -51.240 150.375 ;
        RECT -43.170 150.345 -42.150 150.375 ;
        RECT -51.795 149.595 -51.565 150.345 ;
        RECT -42.845 149.595 -42.615 150.345 ;
        RECT -52.260 149.565 -51.240 149.595 ;
        RECT -43.170 149.565 -42.150 149.595 ;
        RECT -52.720 149.395 -50.280 149.565 ;
        RECT -44.130 149.395 -41.690 149.565 ;
        RECT -52.260 149.365 -51.240 149.395 ;
        RECT -43.170 149.365 -42.150 149.395 ;
        RECT -51.795 148.615 -51.565 149.365 ;
        RECT -42.845 148.615 -42.615 149.365 ;
        RECT -52.260 148.585 -50.300 148.615 ;
        RECT -44.110 148.585 -42.150 148.615 ;
        RECT -52.720 148.415 -50.280 148.585 ;
        RECT -44.130 148.415 -41.690 148.585 ;
        RECT -52.260 148.385 -50.300 148.415 ;
        RECT -44.110 148.385 -42.150 148.415 ;
        RECT -51.210 147.310 -50.390 147.595 ;
        RECT -44.020 147.310 -43.200 147.595 ;
        RECT -42.770 147.365 -42.400 148.205 ;
        RECT -40.395 147.580 -40.200 156.990 ;
        RECT -38.940 156.865 -36.500 157.035 ;
        RECT -38.480 156.835 -37.460 156.865 ;
        RECT -38.175 156.685 -37.825 156.835 ;
        RECT -38.145 156.395 -37.935 156.685 ;
        RECT -38.575 156.095 -37.915 156.395 ;
        RECT -37.430 155.405 -36.610 155.690 ;
        RECT -31.075 155.215 -30.895 177.050 ;
        RECT -30.675 167.700 -30.505 177.540 ;
        RECT -27.210 175.700 -26.940 176.395 ;
        RECT -28.465 175.455 -26.295 175.480 ;
        RECT -29.410 175.285 -25.340 175.455 ;
        RECT -28.465 175.265 -26.295 175.285 ;
        RECT -27.510 174.765 -27.280 175.265 ;
        RECT -28.455 173.910 -26.305 173.930 ;
        RECT -29.410 173.740 -25.340 173.910 ;
        RECT -28.455 173.715 -26.305 173.740 ;
        RECT -28.230 173.235 -28.000 173.715 ;
        RECT -29.410 172.680 -27.785 172.850 ;
        RECT -29.775 172.360 -29.325 172.370 ;
        RECT -29.775 172.190 -28.370 172.360 ;
        RECT -30.720 167.020 -30.490 167.700 ;
        RECT -29.775 167.500 -29.595 172.190 ;
        RECT -27.955 171.380 -27.785 172.680 ;
        RECT -27.180 172.625 -26.910 173.320 ;
        RECT -29.410 171.210 -27.785 171.380 ;
        RECT -27.095 172.190 -25.340 172.360 ;
        RECT -29.410 170.720 -28.220 170.890 ;
        RECT -28.415 169.570 -28.220 170.720 ;
        RECT -27.955 170.215 -27.785 171.210 ;
        RECT -27.550 170.580 -27.280 171.275 ;
        RECT -27.955 170.045 -27.305 170.215 ;
        RECT -29.410 169.400 -28.220 169.570 ;
        RECT -27.475 169.655 -27.305 170.045 ;
        RECT -27.095 170.130 -26.925 172.190 ;
        RECT -26.725 171.210 -25.340 171.380 ;
        RECT -26.725 170.480 -26.555 171.210 ;
        RECT -26.725 170.310 -24.650 170.480 ;
        RECT -27.095 169.960 -24.995 170.130 ;
        RECT -27.475 169.485 -26.560 169.655 ;
        RECT -25.165 169.570 -24.995 169.960 ;
        RECT -28.415 169.390 -28.220 169.400 ;
        RECT -26.730 169.080 -26.560 169.485 ;
        RECT -26.380 169.400 -24.995 169.570 ;
        RECT -26.730 168.910 -25.340 169.080 ;
        RECT -29.775 167.330 -28.370 167.500 ;
        RECT -30.675 166.855 -30.505 167.020 ;
        RECT -27.400 166.835 -27.130 167.530 ;
        RECT -26.730 167.500 -26.560 168.910 ;
        RECT -25.165 168.590 -24.995 169.400 ;
        RECT -26.380 168.420 -24.995 168.590 ;
        RECT -24.820 167.990 -24.650 170.310 ;
        RECT -26.380 167.820 -24.650 167.990 ;
        RECT -26.730 167.330 -25.340 167.500 ;
        RECT -29.245 166.310 -28.565 166.340 ;
        RECT -26.730 166.310 -26.560 167.330 ;
        RECT -24.820 167.010 -24.650 167.820 ;
        RECT -26.380 166.840 -24.650 167.010 ;
        RECT -29.245 166.140 -26.555 166.310 ;
        RECT -29.245 166.110 -28.565 166.140 ;
        RECT -27.210 163.200 -26.940 163.895 ;
        RECT -28.465 162.955 -26.295 162.980 ;
        RECT -29.410 162.785 -25.340 162.955 ;
        RECT -28.465 162.765 -26.295 162.785 ;
        RECT -27.510 162.265 -27.280 162.765 ;
        RECT -28.455 161.410 -26.305 161.430 ;
        RECT -29.410 161.240 -25.340 161.410 ;
        RECT -28.455 161.215 -26.305 161.240 ;
        RECT -28.230 160.735 -28.000 161.215 ;
        RECT -29.410 160.180 -27.785 160.350 ;
        RECT -29.775 159.860 -29.325 159.870 ;
        RECT -29.775 159.690 -28.370 159.860 ;
        RECT -31.075 154.970 -30.425 155.215 ;
        RECT -38.480 154.585 -36.520 154.615 ;
        RECT -38.940 154.415 -36.500 154.585 ;
        RECT -30.655 154.535 -30.425 154.970 ;
        RECT -29.775 155.000 -29.595 159.690 ;
        RECT -27.955 158.880 -27.785 160.180 ;
        RECT -27.180 160.125 -26.910 160.820 ;
        RECT -29.410 158.710 -27.785 158.880 ;
        RECT -27.095 159.690 -25.340 159.860 ;
        RECT -29.410 158.220 -28.220 158.390 ;
        RECT -28.415 157.070 -28.220 158.220 ;
        RECT -27.955 157.715 -27.785 158.710 ;
        RECT -27.550 158.080 -27.280 158.775 ;
        RECT -27.955 157.545 -27.305 157.715 ;
        RECT -29.410 156.900 -28.220 157.070 ;
        RECT -27.475 157.155 -27.305 157.545 ;
        RECT -27.095 157.630 -26.925 159.690 ;
        RECT -26.725 158.710 -25.340 158.880 ;
        RECT -26.725 157.980 -26.555 158.710 ;
        RECT -26.725 157.810 -24.650 157.980 ;
        RECT -27.095 157.460 -24.995 157.630 ;
        RECT -27.475 156.985 -26.560 157.155 ;
        RECT -25.165 157.070 -24.995 157.460 ;
        RECT -28.415 156.890 -28.220 156.900 ;
        RECT -26.730 156.580 -26.560 156.985 ;
        RECT -26.380 156.900 -24.995 157.070 ;
        RECT -26.730 156.410 -25.340 156.580 ;
        RECT -29.775 154.830 -28.370 155.000 ;
        RECT -38.480 154.385 -36.520 154.415 ;
        RECT -38.015 153.635 -37.785 154.385 ;
        RECT -27.400 154.335 -27.130 155.030 ;
        RECT -26.730 155.000 -26.560 156.410 ;
        RECT -25.165 156.090 -24.995 156.900 ;
        RECT -26.380 155.920 -24.995 156.090 ;
        RECT -24.820 155.490 -24.650 157.810 ;
        RECT -26.380 155.320 -24.650 155.490 ;
        RECT -26.730 154.830 -25.340 155.000 ;
        RECT -29.245 153.910 -28.565 153.940 ;
        RECT -26.730 153.910 -26.560 154.830 ;
        RECT -24.820 154.510 -24.650 155.320 ;
        RECT -26.380 154.340 -24.650 154.510 ;
        RECT -29.245 153.740 -26.560 153.910 ;
        RECT -29.245 153.710 -28.565 153.740 ;
        RECT -38.480 153.605 -37.460 153.635 ;
        RECT -38.940 153.435 -36.500 153.605 ;
        RECT -38.480 153.405 -37.460 153.435 ;
        RECT -38.015 152.655 -37.785 153.405 ;
        RECT -38.480 152.625 -37.460 152.655 ;
        RECT -38.940 152.455 -36.500 152.625 ;
        RECT -38.480 152.425 -37.460 152.455 ;
        RECT -38.175 152.150 -37.825 152.425 ;
        RECT -38.175 151.785 -36.865 152.150 ;
        RECT -37.705 151.780 -36.865 151.785 ;
        RECT -39.590 151.530 -39.130 151.555 ;
        RECT -38.780 151.530 -37.000 151.560 ;
        RECT -36.630 151.530 -36.235 151.535 ;
        RECT -39.590 151.360 -36.235 151.530 ;
        RECT -39.590 151.335 -39.130 151.360 ;
        RECT -39.590 150.575 -39.420 151.335 ;
        RECT -38.780 151.325 -37.000 151.360 ;
        RECT -36.630 151.355 -36.235 151.360 ;
        RECT -38.675 151.040 -38.300 151.060 ;
        RECT -39.190 150.870 -38.300 151.040 ;
        RECT -38.675 150.855 -38.300 150.870 ;
        RECT -39.590 150.550 -39.075 150.575 ;
        RECT -39.590 150.380 -38.650 150.550 ;
        RECT -39.590 150.355 -39.075 150.380 ;
        RECT -39.590 149.595 -39.420 150.355 ;
        RECT -38.470 150.070 -38.300 150.855 ;
        RECT -38.105 150.700 -37.735 151.325 ;
        RECT -37.465 151.040 -37.035 151.045 ;
        RECT -37.465 150.870 -36.575 151.040 ;
        RECT -37.465 150.865 -37.035 150.870 ;
        RECT -38.715 150.060 -38.300 150.070 ;
        RECT -39.190 149.890 -38.300 150.060 ;
        RECT -38.715 149.865 -38.300 149.890 ;
        RECT -39.590 149.570 -39.075 149.595 ;
        RECT -39.590 149.400 -38.650 149.570 ;
        RECT -39.590 149.375 -39.075 149.400 ;
        RECT -39.590 148.610 -39.420 149.375 ;
        RECT -38.470 149.100 -38.300 149.865 ;
        RECT -38.715 149.080 -38.300 149.100 ;
        RECT -39.190 148.910 -38.300 149.080 ;
        RECT -38.715 148.895 -38.300 148.910 ;
        RECT -38.470 148.780 -38.300 148.895 ;
        RECT -37.465 150.055 -37.295 150.865 ;
        RECT -36.405 150.555 -36.235 151.355 ;
        RECT -27.210 150.700 -26.940 151.395 ;
        RECT -36.680 150.550 -36.235 150.555 ;
        RECT -37.115 150.380 -36.235 150.550 ;
        RECT -28.465 150.455 -26.295 150.480 ;
        RECT -36.680 150.345 -36.235 150.380 ;
        RECT -37.115 150.055 -36.575 150.060 ;
        RECT -37.465 149.890 -36.575 150.055 ;
        RECT -37.465 149.875 -37.025 149.890 ;
        RECT -37.465 149.085 -37.295 149.875 ;
        RECT -36.405 149.585 -36.235 150.345 ;
        RECT -29.410 150.285 -25.340 150.455 ;
        RECT -28.465 150.265 -26.295 150.285 ;
        RECT -27.510 149.765 -27.280 150.265 ;
        RECT -36.685 149.570 -36.235 149.585 ;
        RECT -37.115 149.400 -36.235 149.570 ;
        RECT -36.685 149.375 -36.235 149.400 ;
        RECT -37.465 149.080 -37.025 149.085 ;
        RECT -37.465 148.910 -36.575 149.080 ;
        RECT -37.465 148.905 -37.025 148.910 ;
        RECT -37.465 148.780 -37.295 148.905 ;
        RECT -39.590 148.590 -39.130 148.610 ;
        RECT -39.590 148.420 -38.650 148.590 ;
        RECT -39.590 148.390 -39.130 148.420 ;
        RECT -39.330 148.115 -38.670 148.145 ;
        RECT -38.470 148.115 -37.295 148.780 ;
        RECT -36.405 148.605 -36.235 149.375 ;
        RECT -28.455 148.910 -26.305 148.930 ;
        RECT -29.410 148.740 -25.340 148.910 ;
        RECT -28.455 148.715 -26.305 148.740 ;
        RECT -36.660 148.590 -36.235 148.605 ;
        RECT -37.115 148.420 -36.235 148.590 ;
        RECT -36.660 148.395 -36.235 148.420 ;
        RECT -28.230 148.235 -28.000 148.715 ;
        RECT -39.330 148.100 -37.075 148.115 ;
        RECT -39.330 147.930 -36.575 148.100 ;
        RECT -39.330 147.915 -37.075 147.930 ;
        RECT -38.720 147.910 -37.075 147.915 ;
        RECT -38.505 147.905 -37.075 147.910 ;
        RECT -50.960 146.880 -50.650 147.310 ;
        RECT -51.955 146.570 -50.650 146.880 ;
        RECT -43.760 146.880 -43.450 147.310 ;
        RECT -42.715 147.065 -41.605 147.365 ;
        RECT -40.445 146.920 -40.145 147.580 ;
        RECT -38.190 146.920 -37.905 147.905 ;
        RECT -29.410 147.680 -27.785 147.850 ;
        RECT -29.775 147.360 -29.325 147.370 ;
        RECT -29.775 147.190 -28.370 147.360 ;
        RECT -43.760 146.570 -42.455 146.880 ;
        RECT -51.955 146.390 -51.605 146.570 ;
        RECT -42.805 146.390 -42.455 146.570 ;
        RECT -52.260 146.360 -51.240 146.390 ;
        RECT -43.170 146.360 -42.150 146.390 ;
        RECT -52.720 146.190 -50.280 146.360 ;
        RECT -44.130 146.190 -41.690 146.360 ;
        RECT -52.260 146.160 -51.240 146.190 ;
        RECT -43.170 146.160 -42.150 146.190 ;
        RECT -51.795 145.410 -51.565 146.160 ;
        RECT -42.845 145.410 -42.615 146.160 ;
        RECT -52.260 145.380 -51.240 145.410 ;
        RECT -43.170 145.380 -42.150 145.410 ;
        RECT -52.720 145.210 -50.280 145.380 ;
        RECT -44.130 145.210 -41.690 145.380 ;
        RECT -52.260 145.180 -51.240 145.210 ;
        RECT -43.170 145.180 -42.150 145.210 ;
        RECT -51.795 144.430 -51.565 145.180 ;
        RECT -42.845 144.430 -42.615 145.180 ;
        RECT -52.260 144.400 -50.300 144.430 ;
        RECT -44.110 144.400 -42.150 144.430 ;
        RECT -52.720 144.230 -50.280 144.400 ;
        RECT -44.130 144.230 -41.690 144.400 ;
        RECT -52.260 144.200 -50.300 144.230 ;
        RECT -44.110 144.200 -42.150 144.230 ;
        RECT -52.010 143.180 -51.640 144.020 ;
        RECT -42.770 143.180 -42.400 144.020 ;
        RECT -51.975 143.070 -51.675 143.180 ;
        RECT -42.735 143.070 -42.435 143.180 ;
        RECT -40.395 142.875 -40.200 146.920 ;
        RECT -38.230 146.080 -37.860 146.920 ;
        RECT -38.480 145.870 -36.520 145.900 ;
        RECT -38.940 145.700 -36.500 145.870 ;
        RECT -38.480 145.670 -36.520 145.700 ;
        RECT -38.015 144.920 -37.785 145.670 ;
        RECT -38.480 144.890 -37.460 144.920 ;
        RECT -38.940 144.720 -36.500 144.890 ;
        RECT -38.480 144.690 -37.460 144.720 ;
        RECT -38.015 143.940 -37.785 144.690 ;
        RECT -38.480 143.910 -37.460 143.940 ;
        RECT -38.940 143.740 -36.500 143.910 ;
        RECT -38.480 143.710 -37.460 143.740 ;
        RECT -38.175 143.560 -37.825 143.710 ;
        RECT -38.120 143.310 -37.895 143.560 ;
        RECT -38.695 143.210 -37.895 143.310 ;
        RECT -38.695 143.010 -37.000 143.210 ;
        RECT -38.120 142.985 -37.000 143.010 ;
        RECT -40.450 142.190 -40.150 142.875 ;
        RECT -38.570 142.435 -37.910 142.735 ;
        RECT -52.080 141.595 -51.780 142.050 ;
        RECT -42.630 141.595 -42.330 142.050 ;
        RECT -52.285 141.590 -50.855 141.595 ;
        RECT -52.500 141.570 -50.855 141.590 ;
        RECT -43.555 141.590 -42.125 141.595 ;
        RECT -43.555 141.570 -41.910 141.590 ;
        RECT -52.970 141.400 -50.355 141.570 ;
        RECT -44.055 141.400 -41.440 141.570 ;
        RECT -52.500 141.385 -50.855 141.400 ;
        RECT -43.555 141.385 -41.910 141.400 ;
        RECT -53.370 141.080 -52.910 141.110 ;
        RECT -53.370 140.910 -52.430 141.080 ;
        RECT -53.370 140.890 -52.910 140.910 ;
        RECT -53.370 140.125 -53.200 140.890 ;
        RECT -52.250 140.720 -51.075 141.385 ;
        RECT -50.440 141.080 -50.015 141.105 ;
        RECT -50.895 140.910 -50.015 141.080 ;
        RECT -50.440 140.895 -50.015 140.910 ;
        RECT -52.250 140.605 -52.080 140.720 ;
        RECT -52.495 140.590 -52.080 140.605 ;
        RECT -52.970 140.420 -52.080 140.590 ;
        RECT -52.495 140.400 -52.080 140.420 ;
        RECT -53.370 140.100 -52.855 140.125 ;
        RECT -53.370 139.930 -52.430 140.100 ;
        RECT -53.370 139.905 -52.855 139.930 ;
        RECT -53.370 139.145 -53.200 139.905 ;
        RECT -52.250 139.635 -52.080 140.400 ;
        RECT -52.495 139.610 -52.080 139.635 ;
        RECT -52.970 139.440 -52.080 139.610 ;
        RECT -52.495 139.430 -52.080 139.440 ;
        RECT -53.370 139.120 -52.855 139.145 ;
        RECT -53.370 138.950 -52.430 139.120 ;
        RECT -53.370 138.925 -52.855 138.950 ;
        RECT -53.370 138.165 -53.200 138.925 ;
        RECT -52.250 138.645 -52.080 139.430 ;
        RECT -51.245 140.595 -51.075 140.720 ;
        RECT -51.245 140.590 -50.805 140.595 ;
        RECT -51.245 140.420 -50.355 140.590 ;
        RECT -51.245 140.415 -50.805 140.420 ;
        RECT -51.245 139.625 -51.075 140.415 ;
        RECT -50.185 140.125 -50.015 140.895 ;
        RECT -50.465 140.100 -50.015 140.125 ;
        RECT -50.895 139.930 -50.015 140.100 ;
        RECT -50.465 139.915 -50.015 139.930 ;
        RECT -51.245 139.610 -50.805 139.625 ;
        RECT -51.245 139.445 -50.355 139.610 ;
        RECT -52.455 138.630 -52.080 138.645 ;
        RECT -52.970 138.460 -52.080 138.630 ;
        RECT -52.455 138.440 -52.080 138.460 ;
        RECT -51.885 138.175 -51.515 138.800 ;
        RECT -51.245 138.635 -51.075 139.445 ;
        RECT -50.895 139.440 -50.355 139.445 ;
        RECT -50.185 139.155 -50.015 139.915 ;
        RECT -50.460 139.120 -50.015 139.155 ;
        RECT -50.895 138.950 -50.015 139.120 ;
        RECT -50.460 138.945 -50.015 138.950 ;
        RECT -51.245 138.630 -50.815 138.635 ;
        RECT -51.245 138.460 -50.355 138.630 ;
        RECT -51.245 138.455 -50.815 138.460 ;
        RECT -53.370 138.140 -52.910 138.165 ;
        RECT -52.560 138.140 -50.780 138.175 ;
        RECT -50.185 138.145 -50.015 138.945 ;
        RECT -50.410 138.140 -50.015 138.145 ;
        RECT -53.370 137.970 -50.015 138.140 ;
        RECT -53.370 137.945 -52.910 137.970 ;
        RECT -52.560 137.940 -50.780 137.970 ;
        RECT -50.410 137.965 -50.015 137.970 ;
        RECT -44.395 141.080 -43.970 141.105 ;
        RECT -44.395 140.910 -43.515 141.080 ;
        RECT -44.395 140.895 -43.970 140.910 ;
        RECT -44.395 140.125 -44.225 140.895 ;
        RECT -43.335 140.720 -42.160 141.385 ;
        RECT -41.500 141.080 -41.040 141.110 ;
        RECT -41.980 140.910 -41.040 141.080 ;
        RECT -41.500 140.890 -41.040 140.910 ;
        RECT -43.335 140.595 -43.165 140.720 ;
        RECT -43.605 140.590 -43.165 140.595 ;
        RECT -44.055 140.420 -43.165 140.590 ;
        RECT -43.605 140.415 -43.165 140.420 ;
        RECT -44.395 140.100 -43.945 140.125 ;
        RECT -44.395 139.930 -43.515 140.100 ;
        RECT -44.395 139.915 -43.945 139.930 ;
        RECT -44.395 139.155 -44.225 139.915 ;
        RECT -43.335 139.625 -43.165 140.415 ;
        RECT -43.605 139.610 -43.165 139.625 ;
        RECT -44.055 139.445 -43.165 139.610 ;
        RECT -44.055 139.440 -43.515 139.445 ;
        RECT -44.395 139.120 -43.950 139.155 ;
        RECT -44.395 138.950 -43.515 139.120 ;
        RECT -44.395 138.945 -43.950 138.950 ;
        RECT -44.395 138.145 -44.225 138.945 ;
        RECT -43.335 138.635 -43.165 139.445 ;
        RECT -42.330 140.605 -42.160 140.720 ;
        RECT -42.330 140.590 -41.915 140.605 ;
        RECT -42.330 140.420 -41.440 140.590 ;
        RECT -42.330 140.400 -41.915 140.420 ;
        RECT -42.330 139.635 -42.160 140.400 ;
        RECT -41.210 140.125 -41.040 140.890 ;
        RECT -41.555 140.100 -41.040 140.125 ;
        RECT -41.980 139.930 -41.040 140.100 ;
        RECT -41.555 139.905 -41.040 139.930 ;
        RECT -42.330 139.610 -41.915 139.635 ;
        RECT -42.330 139.440 -41.440 139.610 ;
        RECT -42.330 139.430 -41.915 139.440 ;
        RECT -43.595 138.630 -43.165 138.635 ;
        RECT -44.055 138.460 -43.165 138.630 ;
        RECT -43.595 138.455 -43.165 138.460 ;
        RECT -42.895 138.175 -42.525 138.800 ;
        RECT -42.330 138.645 -42.160 139.430 ;
        RECT -41.210 139.145 -41.040 139.905 ;
        RECT -41.555 139.120 -41.040 139.145 ;
        RECT -41.980 138.950 -41.040 139.120 ;
        RECT -41.555 138.925 -41.040 138.950 ;
        RECT -42.330 138.630 -41.955 138.645 ;
        RECT -42.330 138.460 -41.440 138.630 ;
        RECT -42.330 138.440 -41.955 138.460 ;
        RECT -44.395 138.140 -44.000 138.145 ;
        RECT -43.630 138.140 -41.850 138.175 ;
        RECT -41.210 138.165 -41.040 138.925 ;
        RECT -41.500 138.140 -41.040 138.165 ;
        RECT -44.395 137.970 -41.040 138.140 ;
        RECT -44.395 137.965 -44.000 137.970 ;
        RECT -43.630 137.940 -41.850 137.970 ;
        RECT -41.500 137.945 -41.040 137.970 ;
        RECT -51.485 137.715 -50.645 137.720 ;
        RECT -51.955 137.350 -50.645 137.715 ;
        RECT -43.765 137.715 -42.925 137.720 ;
        RECT -43.765 137.350 -42.455 137.715 ;
        RECT -51.955 137.075 -51.605 137.350 ;
        RECT -42.805 137.075 -42.455 137.350 ;
        RECT -52.260 137.045 -51.240 137.075 ;
        RECT -43.170 137.045 -42.150 137.075 ;
        RECT -52.720 136.875 -50.280 137.045 ;
        RECT -44.130 136.875 -41.690 137.045 ;
        RECT -52.260 136.845 -51.240 136.875 ;
        RECT -43.170 136.845 -42.150 136.875 ;
        RECT -51.795 136.095 -51.565 136.845 ;
        RECT -42.845 136.095 -42.615 136.845 ;
        RECT -52.260 136.065 -51.240 136.095 ;
        RECT -43.170 136.065 -42.150 136.095 ;
        RECT -52.720 135.895 -50.280 136.065 ;
        RECT -44.130 135.895 -41.690 136.065 ;
        RECT -52.260 135.865 -51.240 135.895 ;
        RECT -43.170 135.865 -42.150 135.895 ;
        RECT -51.795 135.115 -51.565 135.865 ;
        RECT -42.845 135.115 -42.615 135.865 ;
        RECT -52.260 135.085 -50.300 135.115 ;
        RECT -44.110 135.085 -42.150 135.115 ;
        RECT -52.720 134.915 -50.280 135.085 ;
        RECT -44.130 134.915 -41.690 135.085 ;
        RECT -52.260 134.885 -50.300 134.915 ;
        RECT -44.110 134.885 -42.150 134.915 ;
        RECT -56.550 132.580 -56.180 133.420 ;
        RECT -54.705 133.325 -54.405 133.985 ;
        RECT -52.010 133.865 -51.640 134.705 ;
        RECT -52.010 133.805 -51.695 133.865 ;
        RECT -51.210 133.810 -50.390 134.095 ;
        RECT -44.020 133.810 -43.200 134.095 ;
        RECT -52.730 133.690 -51.695 133.805 ;
        RECT -52.730 133.505 -51.700 133.690 ;
        RECT -50.955 133.325 -50.710 133.810 ;
        RECT -57.890 132.370 -55.930 132.400 ;
        RECT -57.910 132.200 -55.470 132.370 ;
        RECT -57.890 132.170 -55.930 132.200 ;
        RECT -56.625 131.420 -56.395 132.170 ;
        RECT -56.950 131.390 -55.930 131.420 ;
        RECT -57.910 131.220 -55.470 131.390 ;
        RECT -54.640 131.295 -54.445 133.325 ;
        RECT -51.955 133.095 -50.710 133.325 ;
        RECT -43.700 133.325 -43.455 133.810 ;
        RECT -43.700 133.095 -42.455 133.325 ;
        RECT -51.955 132.890 -51.605 133.095 ;
        RECT -42.805 132.890 -42.455 133.095 ;
        RECT -52.260 132.860 -51.240 132.890 ;
        RECT -43.170 132.860 -42.150 132.890 ;
        RECT -52.720 132.690 -50.280 132.860 ;
        RECT -44.130 132.690 -41.690 132.860 ;
        RECT -52.260 132.660 -51.240 132.690 ;
        RECT -43.170 132.660 -42.150 132.690 ;
        RECT -51.795 131.910 -51.565 132.660 ;
        RECT -42.845 131.910 -42.615 132.660 ;
        RECT -52.260 131.880 -51.240 131.910 ;
        RECT -43.170 131.880 -42.150 131.910 ;
        RECT -52.720 131.710 -50.280 131.880 ;
        RECT -44.130 131.710 -41.690 131.880 ;
        RECT -52.260 131.680 -51.240 131.710 ;
        RECT -43.170 131.680 -42.150 131.710 ;
        RECT -56.950 131.190 -55.930 131.220 ;
        RECT -56.625 130.440 -56.395 131.190 ;
        RECT -51.795 130.930 -51.565 131.680 ;
        RECT -42.845 130.930 -42.615 131.680 ;
        RECT -40.395 131.295 -40.200 142.190 ;
        RECT -38.205 142.135 -37.915 142.435 ;
        RECT -37.225 142.190 -37.000 142.985 ;
        RECT -29.775 142.500 -29.595 147.190 ;
        RECT -27.955 146.380 -27.785 147.680 ;
        RECT -27.180 147.625 -26.910 148.320 ;
        RECT -29.410 146.210 -27.785 146.380 ;
        RECT -27.095 147.190 -25.340 147.360 ;
        RECT -29.410 145.720 -28.220 145.890 ;
        RECT -28.415 144.570 -28.220 145.720 ;
        RECT -27.955 145.215 -27.785 146.210 ;
        RECT -27.550 145.580 -27.280 146.275 ;
        RECT -27.955 145.045 -27.305 145.215 ;
        RECT -29.410 144.400 -28.220 144.570 ;
        RECT -27.475 144.655 -27.305 145.045 ;
        RECT -27.095 145.130 -26.925 147.190 ;
        RECT -26.725 146.210 -25.340 146.380 ;
        RECT -26.725 145.480 -26.555 146.210 ;
        RECT -26.725 145.310 -24.650 145.480 ;
        RECT -27.095 144.960 -24.995 145.130 ;
        RECT -27.475 144.485 -26.560 144.655 ;
        RECT -25.165 144.570 -24.995 144.960 ;
        RECT -28.415 144.390 -28.220 144.400 ;
        RECT -26.730 144.080 -26.560 144.485 ;
        RECT -26.380 144.400 -24.995 144.570 ;
        RECT -26.730 143.910 -25.340 144.080 ;
        RECT -29.775 142.330 -28.370 142.500 ;
        RECT -38.230 141.295 -37.860 142.135 ;
        RECT -37.430 141.905 -36.610 142.190 ;
        RECT -27.400 141.835 -27.130 142.530 ;
        RECT -26.730 142.500 -26.560 143.910 ;
        RECT -25.165 143.590 -24.995 144.400 ;
        RECT -26.380 143.420 -24.995 143.590 ;
        RECT -24.820 142.990 -24.650 145.310 ;
        RECT -26.380 142.820 -24.650 142.990 ;
        RECT -26.730 142.330 -25.340 142.500 ;
        RECT -34.250 141.185 -34.020 141.665 ;
        RECT -32.755 141.185 -32.075 141.200 ;
        RECT -38.480 141.085 -36.520 141.115 ;
        RECT -38.940 140.915 -36.500 141.085 ;
        RECT -34.250 140.985 -32.075 141.185 ;
        RECT -32.755 140.970 -32.075 140.985 ;
        RECT -29.225 141.170 -28.545 141.200 ;
        RECT -26.730 141.170 -26.560 142.330 ;
        RECT -24.820 142.010 -24.650 142.820 ;
        RECT -26.380 141.840 -24.650 142.010 ;
        RECT -29.225 141.000 -26.560 141.170 ;
        RECT -29.225 140.970 -28.545 141.000 ;
        RECT -38.480 140.885 -36.520 140.915 ;
        RECT -38.015 140.135 -37.785 140.885 ;
        RECT -38.480 140.105 -37.460 140.135 ;
        RECT -38.940 139.935 -36.500 140.105 ;
        RECT -38.480 139.905 -37.460 139.935 ;
        RECT -38.015 139.155 -37.785 139.905 ;
        RECT -38.480 139.125 -37.460 139.155 ;
        RECT -38.940 138.955 -36.500 139.125 ;
        RECT -31.700 139.060 -31.020 139.290 ;
        RECT -38.480 138.925 -37.460 138.955 ;
        RECT -38.175 138.650 -37.825 138.925 ;
        RECT -38.175 138.285 -36.865 138.650 ;
        RECT -37.705 138.280 -36.865 138.285 ;
        RECT -39.590 138.030 -39.130 138.055 ;
        RECT -38.780 138.030 -37.000 138.060 ;
        RECT -36.630 138.030 -36.235 138.035 ;
        RECT -39.590 137.860 -36.235 138.030 ;
        RECT -39.590 137.835 -39.130 137.860 ;
        RECT -39.590 137.075 -39.420 137.835 ;
        RECT -38.780 137.825 -37.000 137.860 ;
        RECT -36.630 137.855 -36.235 137.860 ;
        RECT -38.675 137.540 -38.300 137.560 ;
        RECT -39.190 137.370 -38.300 137.540 ;
        RECT -38.675 137.355 -38.300 137.370 ;
        RECT -39.590 137.050 -39.075 137.075 ;
        RECT -39.590 136.880 -38.650 137.050 ;
        RECT -39.590 136.855 -39.075 136.880 ;
        RECT -39.590 136.095 -39.420 136.855 ;
        RECT -38.470 136.570 -38.300 137.355 ;
        RECT -38.105 137.200 -37.735 137.825 ;
        RECT -37.465 137.540 -37.035 137.545 ;
        RECT -37.465 137.370 -36.575 137.540 ;
        RECT -37.465 137.365 -37.035 137.370 ;
        RECT -38.715 136.560 -38.300 136.570 ;
        RECT -39.190 136.390 -38.300 136.560 ;
        RECT -38.715 136.365 -38.300 136.390 ;
        RECT -39.590 136.070 -39.075 136.095 ;
        RECT -39.590 135.900 -38.650 136.070 ;
        RECT -39.590 135.875 -39.075 135.900 ;
        RECT -39.590 135.110 -39.420 135.875 ;
        RECT -38.470 135.600 -38.300 136.365 ;
        RECT -38.715 135.580 -38.300 135.600 ;
        RECT -39.190 135.410 -38.300 135.580 ;
        RECT -38.715 135.395 -38.300 135.410 ;
        RECT -38.470 135.280 -38.300 135.395 ;
        RECT -37.465 136.555 -37.295 137.365 ;
        RECT -36.405 137.055 -36.235 137.855 ;
        RECT -36.680 137.050 -36.235 137.055 ;
        RECT -37.115 136.880 -36.235 137.050 ;
        RECT -36.680 136.845 -36.235 136.880 ;
        RECT -37.115 136.555 -36.575 136.560 ;
        RECT -37.465 136.390 -36.575 136.555 ;
        RECT -37.465 136.375 -37.025 136.390 ;
        RECT -37.465 135.585 -37.295 136.375 ;
        RECT -36.405 136.085 -36.235 136.845 ;
        RECT -36.685 136.070 -36.235 136.085 ;
        RECT -37.115 135.900 -36.235 136.070 ;
        RECT -36.685 135.875 -36.235 135.900 ;
        RECT -37.465 135.580 -37.025 135.585 ;
        RECT -37.465 135.410 -36.575 135.580 ;
        RECT -37.465 135.405 -37.025 135.410 ;
        RECT -37.465 135.280 -37.295 135.405 ;
        RECT -39.590 135.090 -39.130 135.110 ;
        RECT -39.590 134.920 -38.650 135.090 ;
        RECT -39.590 134.890 -39.130 134.920 ;
        RECT -38.470 134.615 -37.295 135.280 ;
        RECT -36.405 135.105 -36.235 135.875 ;
        RECT -36.660 135.090 -36.235 135.105 ;
        RECT -37.115 134.920 -36.235 135.090 ;
        RECT -36.660 134.895 -36.235 134.920 ;
        RECT -38.720 134.600 -37.075 134.615 ;
        RECT -39.190 134.430 -36.575 134.600 ;
        RECT -38.720 134.410 -37.075 134.430 ;
        RECT -38.505 134.405 -37.075 134.410 ;
        RECT -38.155 133.420 -37.890 134.405 ;
        RECT -31.700 134.175 -31.350 139.060 ;
        RECT -27.210 138.200 -26.940 138.895 ;
        RECT -28.465 137.955 -26.295 137.980 ;
        RECT -29.410 137.785 -25.340 137.955 ;
        RECT -28.465 137.765 -26.295 137.785 ;
        RECT -27.950 136.635 -27.680 137.330 ;
        RECT -27.510 137.265 -27.280 137.765 ;
        RECT -28.455 136.410 -26.305 136.430 ;
        RECT -29.410 136.240 -25.340 136.410 ;
        RECT -28.455 136.215 -26.305 136.240 ;
        RECT -28.230 135.735 -28.000 136.215 ;
        RECT -29.410 135.180 -27.785 135.350 ;
        RECT -29.775 134.860 -29.325 134.870 ;
        RECT -29.775 134.690 -28.370 134.860 ;
        RECT -32.065 134.145 -31.045 134.175 ;
        RECT -33.025 133.975 -30.585 134.145 ;
        RECT -32.065 133.945 -31.045 133.975 ;
        RECT -38.230 132.580 -37.860 133.420 ;
        RECT -31.740 133.195 -31.510 133.945 ;
        RECT -32.065 133.165 -31.045 133.195 ;
        RECT -33.025 132.995 -30.585 133.165 ;
        RECT -32.065 132.965 -31.045 132.995 ;
        RECT -38.480 132.370 -36.520 132.400 ;
        RECT -38.940 132.200 -36.500 132.370 ;
        RECT -31.740 132.215 -31.510 132.965 ;
        RECT -38.480 132.170 -36.520 132.200 ;
        RECT -33.005 132.185 -31.045 132.215 ;
        RECT -38.015 131.420 -37.785 132.170 ;
        RECT -33.025 132.015 -30.585 132.185 ;
        RECT -33.005 131.985 -31.045 132.015 ;
        RECT -38.480 131.390 -37.460 131.420 ;
        RECT -38.940 131.220 -36.500 131.390 ;
        RECT -38.480 131.190 -37.460 131.220 ;
        RECT -52.260 130.900 -50.300 130.930 ;
        RECT -44.110 130.900 -42.150 130.930 ;
        RECT -52.720 130.730 -50.280 130.900 ;
        RECT -44.130 130.730 -41.690 130.900 ;
        RECT -52.260 130.700 -50.300 130.730 ;
        RECT -44.110 130.700 -42.150 130.730 ;
        RECT -56.950 130.410 -55.930 130.440 ;
        RECT -57.910 130.240 -55.470 130.410 ;
        RECT -56.950 130.210 -55.930 130.240 ;
        RECT -56.585 130.060 -56.235 130.210 ;
        RECT -66.040 129.830 -64.635 130.000 ;
        RECT -56.540 129.885 -56.345 130.060 ;
        RECT -54.555 129.885 -53.870 129.940 ;
        RECT -52.010 129.885 -51.640 130.520 ;
        RECT -56.540 129.680 -51.640 129.885 ;
        RECT -42.770 129.885 -42.400 130.520 ;
        RECT -38.015 130.440 -37.785 131.190 ;
        RECT -38.480 130.410 -37.460 130.440 ;
        RECT -38.940 130.240 -36.500 130.410 ;
        RECT -38.480 130.210 -37.460 130.240 ;
        RECT -38.175 130.060 -37.825 130.210 ;
        RECT -40.540 129.885 -39.855 129.940 ;
        RECT -38.065 129.885 -37.870 130.060 ;
        RECT -42.770 129.680 -37.870 129.885 ;
        RECT -29.775 130.000 -29.595 134.690 ;
        RECT -27.955 133.880 -27.785 135.180 ;
        RECT -27.180 135.125 -26.910 135.820 ;
        RECT -29.410 133.710 -27.785 133.880 ;
        RECT -27.095 134.690 -25.340 134.860 ;
        RECT -29.410 133.220 -28.220 133.390 ;
        RECT -28.415 132.070 -28.220 133.220 ;
        RECT -27.955 132.715 -27.785 133.710 ;
        RECT -27.550 133.080 -27.280 133.775 ;
        RECT -27.955 132.545 -27.305 132.715 ;
        RECT -29.410 131.900 -28.220 132.070 ;
        RECT -27.475 132.155 -27.305 132.545 ;
        RECT -27.095 132.630 -26.925 134.690 ;
        RECT -26.725 133.710 -25.340 133.880 ;
        RECT -26.725 132.980 -26.555 133.710 ;
        RECT -26.725 132.810 -24.650 132.980 ;
        RECT -27.095 132.460 -24.995 132.630 ;
        RECT -27.475 131.985 -26.560 132.155 ;
        RECT -25.165 132.070 -24.995 132.460 ;
        RECT -28.415 131.890 -28.220 131.900 ;
        RECT -27.920 131.245 -27.650 131.940 ;
        RECT -26.730 131.580 -26.560 131.985 ;
        RECT -26.380 131.900 -24.995 132.070 ;
        RECT -26.730 131.410 -25.340 131.580 ;
        RECT -29.775 129.830 -28.370 130.000 ;
        RECT -56.540 129.650 -51.790 129.680 ;
        RECT -56.530 129.645 -51.790 129.650 ;
        RECT -42.620 129.650 -37.870 129.680 ;
        RECT -42.620 129.645 -37.880 129.650 ;
        RECT -54.555 129.640 -53.870 129.645 ;
        RECT -40.540 129.640 -39.855 129.645 ;
        RECT -27.400 129.335 -27.130 130.030 ;
        RECT -26.730 130.000 -26.560 131.410 ;
        RECT -25.165 131.090 -24.995 131.900 ;
        RECT -26.380 130.920 -24.995 131.090 ;
        RECT -24.820 130.490 -24.650 132.810 ;
        RECT -26.380 130.320 -24.650 130.490 ;
        RECT -26.730 129.830 -25.340 130.000 ;
        RECT -60.025 128.955 -59.795 129.265 ;
        RECT -67.850 128.785 -59.795 128.955 ;
        RECT -34.660 128.955 -34.430 129.265 ;
        RECT -26.730 128.955 -26.560 129.830 ;
        RECT -24.820 129.510 -24.650 130.320 ;
        RECT -26.380 129.340 -24.650 129.510 ;
        RECT -34.660 128.785 -26.560 128.955 ;
        RECT -60.025 128.585 -59.795 128.785 ;
        RECT -53.425 127.950 -53.105 128.660 ;
        RECT -40.305 128.035 -39.985 128.785 ;
        RECT -34.660 128.585 -34.430 128.785 ;
        RECT -40.305 127.970 -28.520 128.035 ;
        RECT -70.865 126.520 -69.990 127.335 ;
        RECT -70.770 68.735 -70.090 126.520 ;
        RECT -53.360 126.135 -53.190 127.950 ;
        RECT -40.300 127.865 -28.520 127.970 ;
        RECT -52.835 126.575 -52.395 127.235 ;
        RECT -53.420 125.360 -53.145 126.135 ;
        RECT -53.670 125.100 -53.120 125.130 ;
        RECT -55.130 124.930 -53.120 125.100 ;
        RECT -53.670 124.905 -53.120 124.930 ;
        RECT -53.320 123.575 -53.120 124.905 ;
        RECT -52.835 124.785 -52.655 126.575 ;
        RECT -28.690 126.000 -28.520 127.865 ;
        RECT -28.165 126.575 -27.630 127.235 ;
        RECT -52.425 125.590 -51.950 125.610 ;
        RECT -52.425 125.420 -49.030 125.590 ;
        RECT -52.425 125.400 -51.950 125.420 ;
        RECT -52.880 124.010 -52.605 124.785 ;
        RECT -52.425 124.550 -52.245 125.400 ;
        RECT -28.750 125.225 -28.475 126.000 ;
        RECT -29.000 124.965 -28.450 124.995 ;
        RECT -30.460 124.795 -28.450 124.965 ;
        RECT -29.000 124.770 -28.450 124.795 ;
        RECT -52.425 124.535 -51.980 124.550 ;
        RECT -49.070 124.535 -48.690 124.555 ;
        RECT -52.425 124.365 -48.690 124.535 ;
        RECT -52.425 124.340 -51.980 124.365 ;
        RECT -49.070 124.345 -48.690 124.365 ;
        RECT -52.435 124.045 -51.970 124.065 ;
        RECT -52.435 123.875 -49.030 124.045 ;
        RECT -52.435 123.855 -51.970 123.875 ;
        RECT -52.435 123.575 -52.240 123.855 ;
        RECT -53.320 123.360 -52.240 123.575 ;
        RECT -48.860 123.565 -48.690 124.345 ;
        RECT -49.080 123.555 -48.690 123.565 ;
        RECT -52.070 123.385 -48.690 123.555 ;
        RECT -53.420 122.930 -53.220 123.170 ;
        RECT -53.635 122.910 -53.220 122.930 ;
        RECT -55.130 122.740 -53.220 122.910 ;
        RECT -53.635 122.710 -53.220 122.740 ;
        RECT -53.435 122.500 -53.220 122.710 ;
        RECT -52.770 122.670 -52.495 123.360 ;
        RECT -49.080 123.355 -48.690 123.385 ;
        RECT -28.650 123.440 -28.450 124.770 ;
        RECT -28.165 124.650 -27.985 126.575 ;
        RECT -27.755 125.455 -27.280 125.475 ;
        RECT -27.755 125.285 -24.360 125.455 ;
        RECT -27.755 125.265 -27.280 125.285 ;
        RECT -28.210 123.875 -27.935 124.650 ;
        RECT -27.755 124.415 -27.575 125.265 ;
        RECT -27.755 124.400 -27.310 124.415 ;
        RECT -24.400 124.400 -24.020 124.420 ;
        RECT -27.755 124.230 -24.020 124.400 ;
        RECT -27.755 124.205 -27.310 124.230 ;
        RECT -24.400 124.210 -24.020 124.230 ;
        RECT -27.765 123.910 -27.300 123.930 ;
        RECT -27.765 123.740 -24.360 123.910 ;
        RECT -27.765 123.720 -27.300 123.740 ;
        RECT -27.765 123.440 -27.570 123.720 ;
        RECT -28.650 123.225 -27.570 123.440 ;
        RECT -24.190 123.430 -24.020 124.210 ;
        RECT -24.410 123.420 -24.020 123.430 ;
        RECT -27.400 123.250 -24.020 123.420 ;
        RECT -28.750 122.795 -28.550 123.035 ;
        RECT -28.965 122.775 -28.550 122.795 ;
        RECT -30.460 122.605 -28.550 122.775 ;
        RECT -28.965 122.575 -28.550 122.605 ;
        RECT -53.435 122.495 -52.000 122.500 ;
        RECT -53.435 122.325 -49.030 122.495 ;
        RECT -28.765 122.365 -28.550 122.575 ;
        RECT -28.100 122.535 -27.825 123.225 ;
        RECT -24.410 123.220 -24.020 123.250 ;
        RECT -28.765 122.360 -27.330 122.365 ;
        RECT -53.435 122.285 -52.000 122.325 ;
        RECT -69.555 120.835 -68.700 121.835 ;
        RECT -69.500 68.930 -68.820 120.835 ;
        RECT -55.215 120.575 -54.845 120.675 ;
        RECT -53.435 120.575 -53.220 122.285 ;
        RECT -28.765 122.190 -24.360 122.360 ;
        RECT -28.765 122.150 -27.330 122.190 ;
        RECT -36.735 120.900 -36.125 121.780 ;
        RECT -55.215 120.380 -52.680 120.575 ;
        RECT -55.215 119.835 -54.845 120.380 ;
        RECT -56.555 119.625 -54.595 119.655 ;
        RECT -56.575 119.455 -54.135 119.625 ;
        RECT -56.555 119.425 -54.595 119.455 ;
        RECT -55.290 118.675 -55.060 119.425 ;
        RECT -55.615 118.645 -54.595 118.675 ;
        RECT -56.575 118.475 -54.135 118.645 ;
        RECT -55.615 118.445 -54.595 118.475 ;
        RECT -55.290 117.695 -55.060 118.445 ;
        RECT -55.615 117.665 -54.595 117.695 ;
        RECT -56.575 117.495 -54.135 117.665 ;
        RECT -55.615 117.465 -54.595 117.495 ;
        RECT -55.250 117.315 -54.900 117.465 ;
        RECT -55.140 117.025 -54.930 117.315 ;
        RECT -55.160 116.725 -54.500 117.025 ;
        RECT -55.140 116.440 -54.930 116.725 ;
        RECT -53.360 116.570 -53.060 117.230 ;
        RECT -56.465 116.035 -55.645 116.320 ;
        RECT -55.160 116.265 -54.870 116.440 ;
        RECT -55.215 115.425 -54.845 116.265 ;
        RECT -56.555 115.215 -54.595 115.245 ;
        RECT -56.575 115.045 -54.135 115.215 ;
        RECT -56.555 115.015 -54.595 115.045 ;
        RECT -55.290 114.265 -55.060 115.015 ;
        RECT -55.615 114.235 -54.595 114.265 ;
        RECT -56.575 114.065 -54.135 114.235 ;
        RECT -55.615 114.035 -54.595 114.065 ;
        RECT -55.290 113.285 -55.060 114.035 ;
        RECT -55.615 113.255 -54.595 113.285 ;
        RECT -56.575 113.085 -54.135 113.255 ;
        RECT -55.615 113.055 -54.595 113.085 ;
        RECT -55.250 112.780 -54.900 113.055 ;
        RECT -56.210 112.415 -54.900 112.780 ;
        RECT -56.210 112.410 -55.370 112.415 ;
        RECT -56.840 112.160 -56.445 112.165 ;
        RECT -56.075 112.160 -54.295 112.190 ;
        RECT -53.945 112.160 -53.485 112.185 ;
        RECT -56.840 111.990 -53.485 112.160 ;
        RECT -56.840 111.985 -56.445 111.990 ;
        RECT -56.840 111.185 -56.670 111.985 ;
        RECT -56.075 111.955 -54.295 111.990 ;
        RECT -53.945 111.965 -53.485 111.990 ;
        RECT -56.040 111.670 -55.610 111.675 ;
        RECT -56.500 111.500 -55.610 111.670 ;
        RECT -56.040 111.495 -55.610 111.500 ;
        RECT -56.840 111.180 -56.395 111.185 ;
        RECT -56.840 111.010 -55.960 111.180 ;
        RECT -56.840 110.975 -56.395 111.010 ;
        RECT -56.840 110.215 -56.670 110.975 ;
        RECT -56.500 110.685 -55.960 110.690 ;
        RECT -55.780 110.685 -55.610 111.495 ;
        RECT -55.340 111.330 -54.970 111.955 ;
        RECT -54.775 111.670 -54.400 111.690 ;
        RECT -54.775 111.500 -53.885 111.670 ;
        RECT -54.775 111.485 -54.400 111.500 ;
        RECT -56.500 110.520 -55.610 110.685 ;
        RECT -56.050 110.505 -55.610 110.520 ;
        RECT -56.840 110.200 -56.390 110.215 ;
        RECT -56.840 110.030 -55.960 110.200 ;
        RECT -56.840 110.005 -56.390 110.030 ;
        RECT -56.840 109.235 -56.670 110.005 ;
        RECT -55.780 109.715 -55.610 110.505 ;
        RECT -56.050 109.710 -55.610 109.715 ;
        RECT -56.500 109.540 -55.610 109.710 ;
        RECT -56.050 109.535 -55.610 109.540 ;
        RECT -55.780 109.410 -55.610 109.535 ;
        RECT -54.775 110.700 -54.605 111.485 ;
        RECT -53.655 111.205 -53.485 111.965 ;
        RECT -54.000 111.180 -53.485 111.205 ;
        RECT -54.425 111.010 -53.485 111.180 ;
        RECT -54.000 110.985 -53.485 111.010 ;
        RECT -54.775 110.690 -54.360 110.700 ;
        RECT -54.775 110.520 -53.885 110.690 ;
        RECT -54.775 110.495 -54.360 110.520 ;
        RECT -54.775 109.730 -54.605 110.495 ;
        RECT -53.655 110.225 -53.485 110.985 ;
        RECT -54.000 110.200 -53.485 110.225 ;
        RECT -54.425 110.030 -53.485 110.200 ;
        RECT -54.000 110.005 -53.485 110.030 ;
        RECT -54.775 109.710 -54.360 109.730 ;
        RECT -54.775 109.540 -53.885 109.710 ;
        RECT -54.775 109.525 -54.360 109.540 ;
        RECT -54.775 109.410 -54.605 109.525 ;
        RECT -56.840 109.220 -56.415 109.235 ;
        RECT -56.840 109.050 -55.960 109.220 ;
        RECT -56.840 109.025 -56.415 109.050 ;
        RECT -55.780 108.745 -54.605 109.410 ;
        RECT -53.655 109.240 -53.485 110.005 ;
        RECT -53.945 109.220 -53.485 109.240 ;
        RECT -54.425 109.050 -53.485 109.220 ;
        RECT -53.945 109.020 -53.485 109.050 ;
        RECT -54.405 108.745 -53.745 108.775 ;
        RECT -56.000 108.730 -53.745 108.745 ;
        RECT -56.500 108.560 -53.745 108.730 ;
        RECT -56.000 108.545 -53.745 108.560 ;
        RECT -56.000 108.540 -54.355 108.545 ;
        RECT -56.000 108.535 -54.570 108.540 ;
        RECT -55.170 107.550 -54.885 108.535 ;
        RECT -55.215 106.710 -54.845 107.550 ;
        RECT -56.555 106.500 -54.595 106.530 ;
        RECT -56.575 106.330 -54.135 106.500 ;
        RECT -56.555 106.300 -54.595 106.330 ;
        RECT -55.290 105.550 -55.060 106.300 ;
        RECT -55.615 105.520 -54.595 105.550 ;
        RECT -56.575 105.350 -54.135 105.520 ;
        RECT -55.615 105.320 -54.595 105.350 ;
        RECT -55.290 104.570 -55.060 105.320 ;
        RECT -55.615 104.540 -54.595 104.570 ;
        RECT -56.575 104.370 -54.135 104.540 ;
        RECT -55.615 104.340 -54.595 104.370 ;
        RECT -55.250 104.190 -54.900 104.340 ;
        RECT -55.180 103.940 -54.955 104.190 ;
        RECT -55.180 103.840 -54.380 103.940 ;
        RECT -56.075 103.640 -54.380 103.840 ;
        RECT -56.075 103.615 -54.955 103.640 ;
        RECT -56.075 102.820 -55.850 103.615 ;
        RECT -55.165 103.065 -54.505 103.365 ;
        RECT -56.465 102.535 -55.645 102.820 ;
        RECT -55.160 102.765 -54.870 103.065 ;
        RECT -55.215 101.925 -54.845 102.765 ;
        RECT -56.555 101.715 -54.595 101.745 ;
        RECT -56.575 101.545 -54.135 101.715 ;
        RECT -56.555 101.515 -54.595 101.545 ;
        RECT -55.290 100.765 -55.060 101.515 ;
        RECT -55.615 100.735 -54.595 100.765 ;
        RECT -56.575 100.565 -54.135 100.735 ;
        RECT -55.615 100.535 -54.595 100.565 ;
        RECT -55.290 99.785 -55.060 100.535 ;
        RECT -55.615 99.755 -54.595 99.785 ;
        RECT -56.575 99.585 -54.135 99.755 ;
        RECT -55.615 99.555 -54.595 99.585 ;
        RECT -55.250 99.280 -54.900 99.555 ;
        RECT -56.210 98.915 -54.900 99.280 ;
        RECT -56.210 98.910 -55.370 98.915 ;
        RECT -56.840 98.660 -56.445 98.665 ;
        RECT -56.075 98.660 -54.295 98.690 ;
        RECT -53.945 98.660 -53.485 98.685 ;
        RECT -56.840 98.490 -53.485 98.660 ;
        RECT -56.840 98.485 -56.445 98.490 ;
        RECT -56.840 97.685 -56.670 98.485 ;
        RECT -56.075 98.455 -54.295 98.490 ;
        RECT -53.945 98.465 -53.485 98.490 ;
        RECT -56.040 98.170 -55.610 98.175 ;
        RECT -56.500 98.000 -55.610 98.170 ;
        RECT -56.040 97.995 -55.610 98.000 ;
        RECT -56.840 97.680 -56.395 97.685 ;
        RECT -56.840 97.510 -55.960 97.680 ;
        RECT -56.840 97.475 -56.395 97.510 ;
        RECT -56.840 96.715 -56.670 97.475 ;
        RECT -56.500 97.185 -55.960 97.190 ;
        RECT -55.780 97.185 -55.610 97.995 ;
        RECT -55.340 97.830 -54.970 98.455 ;
        RECT -54.775 98.170 -54.400 98.190 ;
        RECT -54.775 98.000 -53.885 98.170 ;
        RECT -54.775 97.985 -54.400 98.000 ;
        RECT -56.500 97.020 -55.610 97.185 ;
        RECT -56.050 97.005 -55.610 97.020 ;
        RECT -56.840 96.700 -56.390 96.715 ;
        RECT -56.840 96.530 -55.960 96.700 ;
        RECT -56.840 96.505 -56.390 96.530 ;
        RECT -56.840 95.735 -56.670 96.505 ;
        RECT -55.780 96.215 -55.610 97.005 ;
        RECT -56.050 96.210 -55.610 96.215 ;
        RECT -56.500 96.040 -55.610 96.210 ;
        RECT -56.050 96.035 -55.610 96.040 ;
        RECT -55.780 95.910 -55.610 96.035 ;
        RECT -54.775 97.200 -54.605 97.985 ;
        RECT -53.655 97.705 -53.485 98.465 ;
        RECT -54.000 97.680 -53.485 97.705 ;
        RECT -54.425 97.510 -53.485 97.680 ;
        RECT -54.000 97.485 -53.485 97.510 ;
        RECT -54.775 97.190 -54.360 97.200 ;
        RECT -54.775 97.020 -53.885 97.190 ;
        RECT -54.775 96.995 -54.360 97.020 ;
        RECT -54.775 96.230 -54.605 96.995 ;
        RECT -53.655 96.725 -53.485 97.485 ;
        RECT -54.000 96.700 -53.485 96.725 ;
        RECT -54.425 96.530 -53.485 96.700 ;
        RECT -54.000 96.505 -53.485 96.530 ;
        RECT -54.775 96.210 -54.360 96.230 ;
        RECT -54.775 96.040 -53.885 96.210 ;
        RECT -54.775 96.025 -54.360 96.040 ;
        RECT -54.775 95.910 -54.605 96.025 ;
        RECT -56.840 95.720 -56.415 95.735 ;
        RECT -56.840 95.550 -55.960 95.720 ;
        RECT -56.840 95.525 -56.415 95.550 ;
        RECT -55.780 95.245 -54.605 95.910 ;
        RECT -53.655 95.740 -53.485 96.505 ;
        RECT -53.945 95.720 -53.485 95.740 ;
        RECT -54.425 95.550 -53.485 95.720 ;
        RECT -53.945 95.520 -53.485 95.550 ;
        RECT -56.000 95.230 -54.355 95.245 ;
        RECT -56.500 95.060 -53.885 95.230 ;
        RECT -56.000 95.040 -54.355 95.060 ;
        RECT -56.000 95.035 -54.570 95.040 ;
        RECT -55.185 94.050 -54.920 95.035 ;
        RECT -53.305 94.615 -53.110 116.570 ;
        RECT -52.875 108.210 -52.680 120.380 ;
        RECT -50.755 115.725 -50.455 116.100 ;
        RECT -50.950 115.720 -49.520 115.725 ;
        RECT -51.165 115.700 -49.520 115.720 ;
        RECT -51.635 115.530 -49.020 115.700 ;
        RECT -51.165 115.515 -49.520 115.530 ;
        RECT -52.035 115.210 -51.575 115.240 ;
        RECT -52.035 115.040 -51.095 115.210 ;
        RECT -52.035 115.020 -51.575 115.040 ;
        RECT -52.035 114.255 -51.865 115.020 ;
        RECT -50.915 114.850 -49.740 115.515 ;
        RECT -49.105 115.210 -48.680 115.235 ;
        RECT -49.560 115.040 -48.680 115.210 ;
        RECT -49.105 115.025 -48.680 115.040 ;
        RECT -50.915 114.735 -50.745 114.850 ;
        RECT -51.160 114.720 -50.745 114.735 ;
        RECT -51.635 114.550 -50.745 114.720 ;
        RECT -51.160 114.530 -50.745 114.550 ;
        RECT -52.035 114.230 -51.520 114.255 ;
        RECT -52.035 114.060 -51.095 114.230 ;
        RECT -52.035 114.035 -51.520 114.060 ;
        RECT -52.035 113.275 -51.865 114.035 ;
        RECT -50.915 113.765 -50.745 114.530 ;
        RECT -51.160 113.740 -50.745 113.765 ;
        RECT -51.635 113.570 -50.745 113.740 ;
        RECT -51.160 113.560 -50.745 113.570 ;
        RECT -52.035 113.250 -51.520 113.275 ;
        RECT -52.035 113.080 -51.095 113.250 ;
        RECT -52.035 113.055 -51.520 113.080 ;
        RECT -52.035 112.295 -51.865 113.055 ;
        RECT -50.915 112.775 -50.745 113.560 ;
        RECT -49.910 114.725 -49.740 114.850 ;
        RECT -49.910 114.720 -49.470 114.725 ;
        RECT -49.910 114.550 -49.020 114.720 ;
        RECT -49.910 114.545 -49.470 114.550 ;
        RECT -49.910 113.755 -49.740 114.545 ;
        RECT -48.850 114.255 -48.680 115.025 ;
        RECT -49.130 114.230 -48.680 114.255 ;
        RECT -49.560 114.060 -48.680 114.230 ;
        RECT -49.130 114.045 -48.680 114.060 ;
        RECT -49.910 113.740 -49.470 113.755 ;
        RECT -49.910 113.575 -49.020 113.740 ;
        RECT -51.120 112.760 -50.745 112.775 ;
        RECT -51.635 112.590 -50.745 112.760 ;
        RECT -51.120 112.570 -50.745 112.590 ;
        RECT -50.550 112.305 -50.180 112.930 ;
        RECT -49.910 112.765 -49.740 113.575 ;
        RECT -49.560 113.570 -49.020 113.575 ;
        RECT -48.850 113.285 -48.680 114.045 ;
        RECT -49.125 113.250 -48.680 113.285 ;
        RECT -49.560 113.080 -48.680 113.250 ;
        RECT -49.125 113.075 -48.680 113.080 ;
        RECT -49.910 112.760 -49.480 112.765 ;
        RECT -49.910 112.590 -49.020 112.760 ;
        RECT -49.910 112.585 -49.480 112.590 ;
        RECT -52.035 112.270 -51.575 112.295 ;
        RECT -51.225 112.270 -49.445 112.305 ;
        RECT -48.850 112.275 -48.680 113.075 ;
        RECT -49.075 112.270 -48.680 112.275 ;
        RECT -52.035 112.100 -48.680 112.270 ;
        RECT -52.035 112.075 -51.575 112.100 ;
        RECT -51.225 112.070 -49.445 112.100 ;
        RECT -49.075 112.095 -48.680 112.100 ;
        RECT -50.150 111.845 -49.310 111.850 ;
        RECT -50.620 111.480 -49.310 111.845 ;
        RECT -50.620 111.205 -50.270 111.480 ;
        RECT -50.925 111.175 -49.905 111.205 ;
        RECT -51.385 111.005 -48.945 111.175 ;
        RECT -50.925 110.975 -49.905 111.005 ;
        RECT -50.460 110.225 -50.230 110.975 ;
        RECT -50.925 110.195 -49.905 110.225 ;
        RECT -51.385 110.025 -48.945 110.195 ;
        RECT -50.925 109.995 -49.905 110.025 ;
        RECT -50.460 109.245 -50.230 109.995 ;
        RECT -50.925 109.215 -48.965 109.245 ;
        RECT -51.385 109.045 -48.945 109.215 ;
        RECT -50.925 109.015 -48.965 109.045 ;
        RECT -52.930 107.550 -52.630 108.210 ;
        RECT -50.675 107.995 -50.305 108.835 ;
        RECT -37.215 108.345 -36.855 108.465 ;
        RECT -51.470 107.695 -50.360 107.995 ;
        RECT -49.875 107.940 -49.055 108.225 ;
        RECT -44.250 107.995 -36.855 108.345 ;
        RECT -52.875 103.505 -52.680 107.550 ;
        RECT -49.625 107.510 -49.315 107.940 ;
        RECT -50.620 107.200 -49.315 107.510 ;
        RECT -50.620 107.020 -50.270 107.200 ;
        RECT -50.925 106.990 -49.905 107.020 ;
        RECT -51.385 106.820 -48.945 106.990 ;
        RECT -50.925 106.790 -49.905 106.820 ;
        RECT -50.460 106.040 -50.230 106.790 ;
        RECT -44.250 106.655 -43.900 107.995 ;
        RECT -37.215 107.940 -36.855 107.995 ;
        RECT -36.340 107.025 -36.125 120.900 ;
        RECT -30.580 120.575 -30.210 120.675 ;
        RECT -28.765 120.575 -28.550 122.150 ;
        RECT -30.580 120.380 -28.045 120.575 ;
        RECT -30.580 119.835 -30.210 120.380 ;
        RECT -28.765 120.360 -28.550 120.380 ;
        RECT -31.920 119.625 -29.960 119.655 ;
        RECT -31.940 119.455 -29.500 119.625 ;
        RECT -31.920 119.425 -29.960 119.455 ;
        RECT -30.655 118.675 -30.425 119.425 ;
        RECT -30.980 118.645 -29.960 118.675 ;
        RECT -31.940 118.475 -29.500 118.645 ;
        RECT -30.980 118.445 -29.960 118.475 ;
        RECT -30.655 117.695 -30.425 118.445 ;
        RECT -30.980 117.665 -29.960 117.695 ;
        RECT -31.940 117.495 -29.500 117.665 ;
        RECT -30.980 117.465 -29.960 117.495 ;
        RECT -30.615 117.315 -30.265 117.465 ;
        RECT -30.505 117.025 -30.295 117.315 ;
        RECT -30.525 116.725 -29.865 117.025 ;
        RECT -30.505 116.440 -30.295 116.725 ;
        RECT -28.725 116.570 -28.425 117.230 ;
        RECT -31.830 116.035 -31.010 116.320 ;
        RECT -30.525 116.265 -30.235 116.440 ;
        RECT -30.580 115.425 -30.210 116.265 ;
        RECT -31.920 115.215 -29.960 115.245 ;
        RECT -31.940 115.045 -29.500 115.215 ;
        RECT -31.920 115.015 -29.960 115.045 ;
        RECT -30.655 114.265 -30.425 115.015 ;
        RECT -30.980 114.235 -29.960 114.265 ;
        RECT -31.940 114.065 -29.500 114.235 ;
        RECT -30.980 114.035 -29.960 114.065 ;
        RECT -30.655 113.285 -30.425 114.035 ;
        RECT -30.980 113.255 -29.960 113.285 ;
        RECT -31.940 113.085 -29.500 113.255 ;
        RECT -30.980 113.055 -29.960 113.085 ;
        RECT -30.615 112.780 -30.265 113.055 ;
        RECT -31.575 112.415 -30.265 112.780 ;
        RECT -31.575 112.410 -30.735 112.415 ;
        RECT -32.205 112.160 -31.810 112.165 ;
        RECT -31.440 112.160 -29.660 112.190 ;
        RECT -29.310 112.160 -28.850 112.185 ;
        RECT -32.205 111.990 -28.850 112.160 ;
        RECT -32.205 111.985 -31.810 111.990 ;
        RECT -32.205 111.185 -32.035 111.985 ;
        RECT -31.440 111.955 -29.660 111.990 ;
        RECT -29.310 111.965 -28.850 111.990 ;
        RECT -31.405 111.670 -30.975 111.675 ;
        RECT -31.865 111.500 -30.975 111.670 ;
        RECT -31.405 111.495 -30.975 111.500 ;
        RECT -32.205 111.180 -31.760 111.185 ;
        RECT -32.205 111.010 -31.325 111.180 ;
        RECT -32.205 110.975 -31.760 111.010 ;
        RECT -32.205 110.215 -32.035 110.975 ;
        RECT -31.865 110.685 -31.325 110.690 ;
        RECT -31.145 110.685 -30.975 111.495 ;
        RECT -30.705 111.330 -30.335 111.955 ;
        RECT -30.140 111.670 -29.765 111.690 ;
        RECT -30.140 111.500 -29.250 111.670 ;
        RECT -30.140 111.485 -29.765 111.500 ;
        RECT -31.865 110.520 -30.975 110.685 ;
        RECT -31.415 110.505 -30.975 110.520 ;
        RECT -32.205 110.200 -31.755 110.215 ;
        RECT -32.205 110.030 -31.325 110.200 ;
        RECT -32.205 110.005 -31.755 110.030 ;
        RECT -32.205 109.235 -32.035 110.005 ;
        RECT -31.145 109.715 -30.975 110.505 ;
        RECT -31.415 109.710 -30.975 109.715 ;
        RECT -31.865 109.540 -30.975 109.710 ;
        RECT -31.415 109.535 -30.975 109.540 ;
        RECT -31.145 109.410 -30.975 109.535 ;
        RECT -30.140 110.700 -29.970 111.485 ;
        RECT -29.020 111.205 -28.850 111.965 ;
        RECT -29.365 111.180 -28.850 111.205 ;
        RECT -29.790 111.010 -28.850 111.180 ;
        RECT -29.365 110.985 -28.850 111.010 ;
        RECT -30.140 110.690 -29.725 110.700 ;
        RECT -30.140 110.520 -29.250 110.690 ;
        RECT -30.140 110.495 -29.725 110.520 ;
        RECT -30.140 109.730 -29.970 110.495 ;
        RECT -29.020 110.225 -28.850 110.985 ;
        RECT -29.365 110.200 -28.850 110.225 ;
        RECT -29.790 110.030 -28.850 110.200 ;
        RECT -29.365 110.005 -28.850 110.030 ;
        RECT -30.140 109.710 -29.725 109.730 ;
        RECT -30.140 109.540 -29.250 109.710 ;
        RECT -30.140 109.525 -29.725 109.540 ;
        RECT -30.140 109.410 -29.970 109.525 ;
        RECT -32.205 109.220 -31.780 109.235 ;
        RECT -32.205 109.050 -31.325 109.220 ;
        RECT -32.205 109.025 -31.780 109.050 ;
        RECT -31.145 108.745 -29.970 109.410 ;
        RECT -29.020 109.240 -28.850 110.005 ;
        RECT -29.310 109.220 -28.850 109.240 ;
        RECT -29.790 109.050 -28.850 109.220 ;
        RECT -29.310 109.020 -28.850 109.050 ;
        RECT -29.770 108.745 -29.110 108.775 ;
        RECT -31.365 108.730 -29.110 108.745 ;
        RECT -31.865 108.560 -29.110 108.730 ;
        RECT -31.365 108.545 -29.110 108.560 ;
        RECT -31.365 108.540 -29.720 108.545 ;
        RECT -31.365 108.535 -29.935 108.540 ;
        RECT -30.535 107.550 -30.250 108.535 ;
        RECT -37.560 106.985 -36.125 107.025 ;
        RECT -40.530 106.815 -36.125 106.985 ;
        RECT -37.560 106.810 -36.125 106.815 ;
        RECT -44.250 106.485 -43.040 106.655 ;
        RECT -50.925 106.010 -49.905 106.040 ;
        RECT -51.385 105.840 -48.945 106.010 ;
        RECT -44.735 105.995 -44.195 106.165 ;
        RECT -40.870 105.925 -40.480 105.955 ;
        RECT -37.065 105.950 -36.790 106.640 ;
        RECT -36.340 106.600 -36.125 106.810 ;
        RECT -30.580 106.710 -30.210 107.550 ;
        RECT -36.340 106.570 -35.925 106.600 ;
        RECT -36.340 106.400 -34.430 106.570 ;
        RECT -31.920 106.500 -29.960 106.530 ;
        RECT -36.340 106.380 -35.925 106.400 ;
        RECT -36.340 106.140 -36.140 106.380 ;
        RECT -31.940 106.330 -29.500 106.500 ;
        RECT -31.920 106.300 -29.960 106.330 ;
        RECT -50.925 105.810 -49.905 105.840 ;
        RECT -50.460 105.060 -50.230 105.810 ;
        RECT -40.870 105.755 -37.490 105.925 ;
        RECT -40.870 105.745 -40.480 105.755 ;
        RECT -43.580 105.505 -43.040 105.675 ;
        RECT -50.925 105.030 -48.965 105.060 ;
        RECT -51.385 104.860 -48.945 105.030 ;
        RECT -44.735 105.015 -44.195 105.185 ;
        RECT -40.870 104.965 -40.700 105.745 ;
        RECT -37.320 105.735 -36.240 105.950 ;
        RECT -37.320 105.455 -37.125 105.735 ;
        RECT -37.590 105.435 -37.125 105.455 ;
        RECT -40.530 105.265 -37.125 105.435 ;
        RECT -37.590 105.245 -37.125 105.265 ;
        RECT -40.870 104.945 -40.490 104.965 ;
        RECT -37.580 104.945 -37.135 104.970 ;
        RECT -50.925 104.830 -48.965 104.860 ;
        RECT -40.870 104.775 -37.135 104.945 ;
        RECT -40.870 104.755 -40.490 104.775 ;
        RECT -37.580 104.760 -37.135 104.775 ;
        RECT -50.675 103.810 -50.305 104.650 ;
        RECT -43.580 104.525 -43.040 104.695 ;
        RECT -44.050 103.935 -43.750 104.300 ;
        RECT -50.640 103.700 -50.340 103.810 ;
        RECT -44.020 103.630 -43.815 103.935 ;
        RECT -37.315 103.910 -37.135 104.760 ;
        RECT -36.955 104.525 -36.680 105.300 ;
        RECT -37.610 103.890 -37.135 103.910 ;
        RECT -40.530 103.720 -37.135 103.890 ;
        RECT -37.610 103.700 -37.135 103.720 ;
        RECT -44.915 103.575 -43.815 103.630 ;
        RECT -52.925 102.820 -52.625 103.505 ;
        RECT -44.955 103.435 -43.815 103.575 ;
        RECT -44.955 103.325 -43.955 103.435 ;
        RECT -47.270 102.950 -45.730 103.120 ;
        RECT -45.545 102.890 -45.190 103.260 ;
        RECT -55.215 93.210 -54.845 94.050 ;
        RECT -53.370 93.955 -53.070 94.615 ;
        RECT -56.555 93.000 -54.595 93.030 ;
        RECT -56.575 92.830 -54.135 93.000 ;
        RECT -56.555 92.800 -54.595 92.830 ;
        RECT -55.290 92.050 -55.060 92.800 ;
        RECT -55.615 92.020 -54.595 92.050 ;
        RECT -56.575 91.850 -54.135 92.020 ;
        RECT -53.305 91.925 -53.110 93.955 ;
        RECT -52.875 91.925 -52.680 102.820 ;
        RECT -50.745 102.225 -50.445 102.680 ;
        RECT -47.270 102.460 -45.730 102.630 ;
        RECT -50.950 102.220 -49.520 102.225 ;
        RECT -51.165 102.200 -49.520 102.220 ;
        RECT -51.635 102.030 -49.020 102.200 ;
        RECT -51.165 102.015 -49.520 102.030 ;
        RECT -52.035 101.710 -51.575 101.740 ;
        RECT -52.035 101.540 -51.095 101.710 ;
        RECT -52.035 101.520 -51.575 101.540 ;
        RECT -52.035 100.755 -51.865 101.520 ;
        RECT -50.915 101.350 -49.740 102.015 ;
        RECT -47.270 101.970 -45.730 102.140 ;
        RECT -49.105 101.710 -48.680 101.735 ;
        RECT -49.560 101.540 -48.680 101.710 ;
        RECT -49.105 101.525 -48.680 101.540 ;
        RECT -50.915 101.235 -50.745 101.350 ;
        RECT -51.160 101.220 -50.745 101.235 ;
        RECT -51.635 101.050 -50.745 101.220 ;
        RECT -51.160 101.030 -50.745 101.050 ;
        RECT -52.035 100.730 -51.520 100.755 ;
        RECT -52.035 100.560 -51.095 100.730 ;
        RECT -52.035 100.535 -51.520 100.560 ;
        RECT -52.035 99.775 -51.865 100.535 ;
        RECT -50.915 100.265 -50.745 101.030 ;
        RECT -51.160 100.240 -50.745 100.265 ;
        RECT -51.635 100.070 -50.745 100.240 ;
        RECT -51.160 100.060 -50.745 100.070 ;
        RECT -52.035 99.750 -51.520 99.775 ;
        RECT -52.035 99.580 -51.095 99.750 ;
        RECT -52.035 99.555 -51.520 99.580 ;
        RECT -52.035 98.795 -51.865 99.555 ;
        RECT -50.915 99.275 -50.745 100.060 ;
        RECT -49.910 101.225 -49.740 101.350 ;
        RECT -49.910 101.220 -49.470 101.225 ;
        RECT -49.910 101.050 -49.020 101.220 ;
        RECT -49.910 101.045 -49.470 101.050 ;
        RECT -49.910 100.255 -49.740 101.045 ;
        RECT -48.850 100.755 -48.680 101.525 ;
        RECT -45.515 101.185 -45.320 102.890 ;
        RECT -44.955 102.630 -44.765 103.325 ;
        RECT -39.230 102.850 -38.880 102.880 ;
        RECT -36.905 102.850 -36.725 104.525 ;
        RECT -36.440 104.405 -36.240 105.735 ;
        RECT -30.655 105.550 -30.425 106.300 ;
        RECT -30.980 105.520 -29.960 105.550 ;
        RECT -31.940 105.350 -29.500 105.520 ;
        RECT -30.980 105.320 -29.960 105.350 ;
        RECT -30.655 104.570 -30.425 105.320 ;
        RECT -30.980 104.540 -29.960 104.570 ;
        RECT -36.440 104.380 -35.890 104.405 ;
        RECT -36.440 104.210 -34.430 104.380 ;
        RECT -31.940 104.370 -29.500 104.540 ;
        RECT -30.980 104.340 -29.960 104.370 ;
        RECT -36.440 104.180 -35.890 104.210 ;
        RECT -30.615 104.190 -30.265 104.340 ;
        RECT -36.415 103.175 -36.140 103.950 ;
        RECT -30.545 103.940 -30.320 104.190 ;
        RECT -30.545 103.840 -29.745 103.940 ;
        RECT -31.440 103.640 -29.745 103.840 ;
        RECT -31.440 103.615 -30.320 103.640 ;
        RECT -36.370 102.990 -36.200 103.175 ;
        RECT -44.955 102.460 -43.045 102.630 ;
        RECT -39.230 102.500 -36.715 102.850 ;
        RECT -31.440 102.820 -31.215 103.615 ;
        RECT -30.530 103.065 -29.870 103.365 ;
        RECT -31.830 102.535 -31.010 102.820 ;
        RECT -30.525 102.765 -30.235 103.065 ;
        RECT -44.955 101.650 -44.765 102.460 ;
        RECT -39.230 101.660 -38.880 102.500 ;
        RECT -30.580 101.925 -30.210 102.765 ;
        RECT -31.920 101.715 -29.960 101.745 ;
        RECT -44.955 101.480 -43.045 101.650 ;
        RECT -40.090 101.490 -38.880 101.660 ;
        RECT -31.940 101.545 -29.500 101.715 ;
        RECT -31.920 101.515 -29.960 101.545 ;
        RECT -47.270 100.990 -45.730 101.160 ;
        RECT -45.520 100.835 -45.320 101.185 ;
        RECT -45.520 100.830 -45.310 100.835 ;
        RECT -49.130 100.730 -48.680 100.755 ;
        RECT -49.560 100.560 -48.680 100.730 ;
        RECT -49.130 100.545 -48.680 100.560 ;
        RECT -49.910 100.240 -49.470 100.255 ;
        RECT -49.910 100.075 -49.020 100.240 ;
        RECT -51.120 99.260 -50.745 99.275 ;
        RECT -51.635 99.090 -50.745 99.260 ;
        RECT -51.120 99.070 -50.745 99.090 ;
        RECT -50.550 98.805 -50.180 99.430 ;
        RECT -49.910 99.265 -49.740 100.075 ;
        RECT -49.560 100.070 -49.020 100.075 ;
        RECT -48.850 99.785 -48.680 100.545 ;
        RECT -49.125 99.750 -48.680 99.785 ;
        RECT -49.560 99.580 -48.680 99.750 ;
        RECT -49.125 99.575 -48.680 99.580 ;
        RECT -49.910 99.260 -49.480 99.265 ;
        RECT -49.910 99.090 -49.020 99.260 ;
        RECT -49.910 99.085 -49.480 99.090 ;
        RECT -52.035 98.770 -51.575 98.795 ;
        RECT -51.225 98.770 -49.445 98.805 ;
        RECT -48.850 98.775 -48.680 99.575 ;
        RECT -49.075 98.770 -48.680 98.775 ;
        RECT -52.035 98.600 -48.680 98.770 ;
        RECT -52.035 98.575 -51.575 98.600 ;
        RECT -51.225 98.570 -49.445 98.600 ;
        RECT -49.075 98.595 -48.680 98.600 ;
        RECT -50.150 98.345 -49.310 98.350 ;
        RECT -50.620 97.980 -49.310 98.345 ;
        RECT -45.510 98.255 -45.310 100.830 ;
        RECT -45.070 100.565 -44.800 101.240 ;
        RECT -38.935 101.000 -38.395 101.170 ;
        RECT -30.655 100.765 -30.425 101.515 ;
        RECT -30.980 100.735 -29.960 100.765 ;
        RECT -45.030 100.465 -44.830 100.565 ;
        RECT -40.090 100.510 -39.550 100.680 ;
        RECT -31.940 100.565 -29.500 100.735 ;
        RECT -30.980 100.535 -29.960 100.565 ;
        RECT -45.020 99.430 -44.840 100.465 ;
        RECT -38.935 100.020 -38.395 100.190 ;
        RECT -30.655 99.785 -30.425 100.535 ;
        RECT -30.980 99.755 -29.960 99.785 ;
        RECT -40.090 99.530 -39.550 99.700 ;
        RECT -31.940 99.585 -29.500 99.755 ;
        RECT -30.980 99.555 -29.960 99.585 ;
        RECT -39.380 98.940 -39.080 99.305 ;
        RECT -30.615 99.280 -30.265 99.555 ;
        RECT -44.730 98.575 -43.690 98.745 ;
        RECT -39.315 98.635 -39.110 98.940 ;
        RECT -31.575 98.915 -30.265 99.280 ;
        RECT -31.575 98.910 -30.735 98.915 ;
        RECT -32.205 98.660 -31.810 98.665 ;
        RECT -31.440 98.660 -29.660 98.690 ;
        RECT -29.310 98.660 -28.850 98.685 ;
        RECT -39.315 98.580 -38.215 98.635 ;
        RECT -39.315 98.440 -38.175 98.580 ;
        RECT -39.175 98.330 -38.175 98.440 ;
        RECT -46.380 98.090 -45.310 98.255 ;
        RECT -46.380 98.085 -45.340 98.090 ;
        RECT -50.620 97.705 -50.270 97.980 ;
        RECT -50.925 97.675 -49.905 97.705 ;
        RECT -51.385 97.505 -48.945 97.675 ;
        RECT -44.730 97.595 -43.690 97.765 ;
        RECT -38.365 97.635 -38.175 98.330 ;
        RECT -32.205 98.490 -28.850 98.660 ;
        RECT -32.205 98.485 -31.810 98.490 ;
        RECT -37.400 97.955 -35.860 98.125 ;
        RECT -32.205 97.685 -32.035 98.485 ;
        RECT -31.440 98.455 -29.660 98.490 ;
        RECT -29.310 98.465 -28.850 98.490 ;
        RECT -31.405 98.170 -30.975 98.175 ;
        RECT -31.865 98.000 -30.975 98.170 ;
        RECT -31.405 97.995 -30.975 98.000 ;
        RECT -32.205 97.680 -31.760 97.685 ;
        RECT -50.925 97.475 -49.905 97.505 ;
        RECT -50.460 96.725 -50.230 97.475 ;
        RECT -40.085 97.465 -38.175 97.635 ;
        RECT -37.400 97.465 -35.860 97.635 ;
        RECT -32.205 97.510 -31.325 97.680 ;
        RECT -32.205 97.475 -31.760 97.510 ;
        RECT -46.380 97.105 -45.340 97.275 ;
        RECT -50.925 96.695 -49.905 96.725 ;
        RECT -51.385 96.525 -48.945 96.695 ;
        RECT -44.730 96.615 -43.690 96.785 ;
        RECT -38.365 96.655 -38.175 97.465 ;
        RECT -37.400 96.975 -35.860 97.145 ;
        RECT -50.925 96.495 -49.905 96.525 ;
        RECT -50.460 95.745 -50.230 96.495 ;
        RECT -40.085 96.485 -38.175 96.655 ;
        RECT -32.205 96.715 -32.035 97.475 ;
        RECT -31.865 97.185 -31.325 97.190 ;
        RECT -31.145 97.185 -30.975 97.995 ;
        RECT -30.705 97.830 -30.335 98.455 ;
        RECT -30.140 98.170 -29.765 98.190 ;
        RECT -30.140 98.000 -29.250 98.170 ;
        RECT -30.140 97.985 -29.765 98.000 ;
        RECT -31.865 97.020 -30.975 97.185 ;
        RECT -31.415 97.005 -30.975 97.020 ;
        RECT -32.205 96.700 -31.755 96.715 ;
        RECT -32.205 96.530 -31.325 96.700 ;
        RECT -32.205 96.505 -31.755 96.530 ;
        RECT -50.925 95.715 -48.965 95.745 ;
        RECT -51.385 95.545 -48.945 95.715 ;
        RECT -38.330 95.570 -38.060 96.245 ;
        RECT -37.400 95.995 -35.860 96.165 ;
        RECT -32.205 95.735 -32.035 96.505 ;
        RECT -31.145 96.215 -30.975 97.005 ;
        RECT -31.415 96.210 -30.975 96.215 ;
        RECT -31.865 96.040 -30.975 96.210 ;
        RECT -31.415 96.035 -30.975 96.040 ;
        RECT -31.145 95.910 -30.975 96.035 ;
        RECT -30.140 97.200 -29.970 97.985 ;
        RECT -29.020 97.705 -28.850 98.465 ;
        RECT -29.365 97.680 -28.850 97.705 ;
        RECT -29.790 97.510 -28.850 97.680 ;
        RECT -29.365 97.485 -28.850 97.510 ;
        RECT -30.140 97.190 -29.725 97.200 ;
        RECT -30.140 97.020 -29.250 97.190 ;
        RECT -30.140 96.995 -29.725 97.020 ;
        RECT -30.140 96.230 -29.970 96.995 ;
        RECT -29.020 96.725 -28.850 97.485 ;
        RECT -29.365 96.700 -28.850 96.725 ;
        RECT -29.790 96.530 -28.850 96.700 ;
        RECT -29.365 96.505 -28.850 96.530 ;
        RECT -30.140 96.210 -29.725 96.230 ;
        RECT -30.140 96.040 -29.250 96.210 ;
        RECT -30.140 96.025 -29.725 96.040 ;
        RECT -30.140 95.910 -29.970 96.025 ;
        RECT -32.205 95.720 -31.780 95.735 ;
        RECT -50.925 95.515 -48.965 95.545 ;
        RECT -38.300 95.470 -38.100 95.570 ;
        RECT -32.205 95.550 -31.325 95.720 ;
        RECT -32.205 95.525 -31.780 95.550 ;
        RECT -50.675 94.495 -50.305 95.335 ;
        RECT -50.675 94.435 -50.360 94.495 ;
        RECT -49.875 94.440 -49.055 94.725 ;
        RECT -51.395 94.320 -50.360 94.435 ;
        RECT -51.395 94.135 -50.365 94.320 ;
        RECT -49.620 93.955 -49.375 94.440 ;
        RECT -38.290 94.200 -38.110 95.470 ;
        RECT -31.145 95.245 -29.970 95.910 ;
        RECT -29.020 95.740 -28.850 96.505 ;
        RECT -29.310 95.720 -28.850 95.740 ;
        RECT -29.790 95.550 -28.850 95.720 ;
        RECT -29.310 95.520 -28.850 95.550 ;
        RECT -31.365 95.230 -29.720 95.245 ;
        RECT -31.865 95.060 -29.250 95.230 ;
        RECT -31.365 95.040 -29.720 95.060 ;
        RECT -31.365 95.035 -29.935 95.040 ;
        RECT -50.620 93.725 -49.375 93.955 ;
        RECT -50.620 93.520 -50.270 93.725 ;
        RECT -50.925 93.490 -49.905 93.520 ;
        RECT -51.385 93.320 -48.945 93.490 ;
        RECT -50.925 93.290 -49.905 93.320 ;
        RECT -50.460 92.540 -50.230 93.290 ;
        RECT -38.595 93.270 -37.825 94.200 ;
        RECT -30.550 94.050 -30.285 95.035 ;
        RECT -28.670 94.615 -28.475 116.570 ;
        RECT -28.240 108.210 -28.045 120.380 ;
        RECT -26.120 115.725 -25.820 116.100 ;
        RECT -26.315 115.720 -24.885 115.725 ;
        RECT -26.530 115.700 -24.885 115.720 ;
        RECT -27.000 115.530 -24.385 115.700 ;
        RECT -26.530 115.515 -24.885 115.530 ;
        RECT -27.400 115.210 -26.940 115.240 ;
        RECT -27.400 115.040 -26.460 115.210 ;
        RECT -27.400 115.020 -26.940 115.040 ;
        RECT -27.400 114.255 -27.230 115.020 ;
        RECT -26.280 114.850 -25.105 115.515 ;
        RECT -24.470 115.210 -24.045 115.235 ;
        RECT -24.925 115.040 -24.045 115.210 ;
        RECT -24.470 115.025 -24.045 115.040 ;
        RECT -26.280 114.735 -26.110 114.850 ;
        RECT -26.525 114.720 -26.110 114.735 ;
        RECT -27.000 114.550 -26.110 114.720 ;
        RECT -26.525 114.530 -26.110 114.550 ;
        RECT -27.400 114.230 -26.885 114.255 ;
        RECT -27.400 114.060 -26.460 114.230 ;
        RECT -27.400 114.035 -26.885 114.060 ;
        RECT -27.400 113.275 -27.230 114.035 ;
        RECT -26.280 113.765 -26.110 114.530 ;
        RECT -26.525 113.740 -26.110 113.765 ;
        RECT -27.000 113.570 -26.110 113.740 ;
        RECT -26.525 113.560 -26.110 113.570 ;
        RECT -27.400 113.250 -26.885 113.275 ;
        RECT -27.400 113.080 -26.460 113.250 ;
        RECT -27.400 113.055 -26.885 113.080 ;
        RECT -27.400 112.295 -27.230 113.055 ;
        RECT -26.280 112.775 -26.110 113.560 ;
        RECT -25.275 114.725 -25.105 114.850 ;
        RECT -25.275 114.720 -24.835 114.725 ;
        RECT -25.275 114.550 -24.385 114.720 ;
        RECT -25.275 114.545 -24.835 114.550 ;
        RECT -25.275 113.755 -25.105 114.545 ;
        RECT -24.215 114.255 -24.045 115.025 ;
        RECT -24.495 114.230 -24.045 114.255 ;
        RECT -24.925 114.060 -24.045 114.230 ;
        RECT -24.495 114.045 -24.045 114.060 ;
        RECT -25.275 113.740 -24.835 113.755 ;
        RECT -25.275 113.575 -24.385 113.740 ;
        RECT -26.485 112.760 -26.110 112.775 ;
        RECT -27.000 112.590 -26.110 112.760 ;
        RECT -26.485 112.570 -26.110 112.590 ;
        RECT -25.915 112.305 -25.545 112.930 ;
        RECT -25.275 112.765 -25.105 113.575 ;
        RECT -24.925 113.570 -24.385 113.575 ;
        RECT -24.215 113.285 -24.045 114.045 ;
        RECT -24.490 113.250 -24.045 113.285 ;
        RECT -24.925 113.080 -24.045 113.250 ;
        RECT -24.490 113.075 -24.045 113.080 ;
        RECT -25.275 112.760 -24.845 112.765 ;
        RECT -25.275 112.590 -24.385 112.760 ;
        RECT -25.275 112.585 -24.845 112.590 ;
        RECT -27.400 112.270 -26.940 112.295 ;
        RECT -26.590 112.270 -24.810 112.305 ;
        RECT -24.215 112.275 -24.045 113.075 ;
        RECT -24.440 112.270 -24.045 112.275 ;
        RECT -27.400 112.100 -24.045 112.270 ;
        RECT -27.400 112.075 -26.940 112.100 ;
        RECT -26.590 112.070 -24.810 112.100 ;
        RECT -24.440 112.095 -24.045 112.100 ;
        RECT -25.515 111.845 -24.675 111.850 ;
        RECT -25.985 111.480 -24.675 111.845 ;
        RECT -25.985 111.205 -25.635 111.480 ;
        RECT -26.290 111.175 -25.270 111.205 ;
        RECT -26.750 111.005 -24.310 111.175 ;
        RECT -26.290 110.975 -25.270 111.005 ;
        RECT -25.825 110.225 -25.595 110.975 ;
        RECT -26.290 110.195 -25.270 110.225 ;
        RECT -26.750 110.025 -24.310 110.195 ;
        RECT -26.290 109.995 -25.270 110.025 ;
        RECT -25.825 109.245 -25.595 109.995 ;
        RECT -26.290 109.215 -24.330 109.245 ;
        RECT -26.750 109.045 -24.310 109.215 ;
        RECT -26.290 109.015 -24.330 109.045 ;
        RECT -28.295 107.550 -27.995 108.210 ;
        RECT -26.040 107.995 -25.670 108.835 ;
        RECT -26.835 107.695 -25.725 107.995 ;
        RECT -25.240 107.940 -24.420 108.225 ;
        RECT -28.240 103.505 -28.045 107.550 ;
        RECT -24.990 107.510 -24.680 107.940 ;
        RECT -25.985 107.200 -24.680 107.510 ;
        RECT -25.985 107.020 -25.635 107.200 ;
        RECT -26.290 106.990 -25.270 107.020 ;
        RECT -26.750 106.820 -24.310 106.990 ;
        RECT -26.290 106.790 -25.270 106.820 ;
        RECT -25.825 106.040 -25.595 106.790 ;
        RECT -26.290 106.010 -25.270 106.040 ;
        RECT -26.750 105.840 -24.310 106.010 ;
        RECT -26.290 105.810 -25.270 105.840 ;
        RECT -25.825 105.060 -25.595 105.810 ;
        RECT -26.290 105.030 -24.330 105.060 ;
        RECT -26.750 104.860 -24.310 105.030 ;
        RECT -26.290 104.830 -24.330 104.860 ;
        RECT -26.040 103.810 -25.670 104.650 ;
        RECT -26.005 103.700 -25.705 103.810 ;
        RECT -28.290 102.820 -27.990 103.505 ;
        RECT -30.580 93.210 -30.210 94.050 ;
        RECT -28.735 93.955 -28.435 94.615 ;
        RECT -31.920 93.000 -29.960 93.030 ;
        RECT -31.940 92.830 -29.500 93.000 ;
        RECT -31.920 92.800 -29.960 92.830 ;
        RECT -50.925 92.510 -49.905 92.540 ;
        RECT -51.385 92.340 -48.945 92.510 ;
        RECT -50.925 92.310 -49.905 92.340 ;
        RECT -55.615 91.820 -54.595 91.850 ;
        RECT -55.290 91.070 -55.060 91.820 ;
        RECT -50.460 91.560 -50.230 92.310 ;
        RECT -30.655 92.050 -30.425 92.800 ;
        RECT -30.980 92.020 -29.960 92.050 ;
        RECT -31.940 91.850 -29.500 92.020 ;
        RECT -28.670 91.925 -28.475 93.955 ;
        RECT -28.240 91.925 -28.045 102.820 ;
        RECT -26.110 102.225 -25.810 102.680 ;
        RECT -26.315 102.220 -24.885 102.225 ;
        RECT -26.530 102.200 -24.885 102.220 ;
        RECT -27.000 102.030 -24.385 102.200 ;
        RECT -26.530 102.015 -24.885 102.030 ;
        RECT -27.400 101.710 -26.940 101.740 ;
        RECT -27.400 101.540 -26.460 101.710 ;
        RECT -27.400 101.520 -26.940 101.540 ;
        RECT -27.400 100.755 -27.230 101.520 ;
        RECT -26.280 101.350 -25.105 102.015 ;
        RECT -24.470 101.710 -24.045 101.735 ;
        RECT -24.925 101.540 -24.045 101.710 ;
        RECT -24.470 101.525 -24.045 101.540 ;
        RECT -26.280 101.235 -26.110 101.350 ;
        RECT -26.525 101.220 -26.110 101.235 ;
        RECT -27.000 101.050 -26.110 101.220 ;
        RECT -26.525 101.030 -26.110 101.050 ;
        RECT -27.400 100.730 -26.885 100.755 ;
        RECT -27.400 100.560 -26.460 100.730 ;
        RECT -27.400 100.535 -26.885 100.560 ;
        RECT -27.400 99.775 -27.230 100.535 ;
        RECT -26.280 100.265 -26.110 101.030 ;
        RECT -26.525 100.240 -26.110 100.265 ;
        RECT -27.000 100.070 -26.110 100.240 ;
        RECT -26.525 100.060 -26.110 100.070 ;
        RECT -27.400 99.750 -26.885 99.775 ;
        RECT -27.400 99.580 -26.460 99.750 ;
        RECT -27.400 99.555 -26.885 99.580 ;
        RECT -27.400 98.795 -27.230 99.555 ;
        RECT -26.280 99.275 -26.110 100.060 ;
        RECT -25.275 101.225 -25.105 101.350 ;
        RECT -25.275 101.220 -24.835 101.225 ;
        RECT -25.275 101.050 -24.385 101.220 ;
        RECT -25.275 101.045 -24.835 101.050 ;
        RECT -25.275 100.255 -25.105 101.045 ;
        RECT -24.215 100.755 -24.045 101.525 ;
        RECT -24.495 100.730 -24.045 100.755 ;
        RECT -24.925 100.560 -24.045 100.730 ;
        RECT -24.495 100.545 -24.045 100.560 ;
        RECT -25.275 100.240 -24.835 100.255 ;
        RECT -25.275 100.075 -24.385 100.240 ;
        RECT -26.485 99.260 -26.110 99.275 ;
        RECT -27.000 99.090 -26.110 99.260 ;
        RECT -26.485 99.070 -26.110 99.090 ;
        RECT -25.915 98.805 -25.545 99.430 ;
        RECT -25.275 99.265 -25.105 100.075 ;
        RECT -24.925 100.070 -24.385 100.075 ;
        RECT -24.215 99.785 -24.045 100.545 ;
        RECT -24.490 99.750 -24.045 99.785 ;
        RECT -24.925 99.580 -24.045 99.750 ;
        RECT -24.490 99.575 -24.045 99.580 ;
        RECT -25.275 99.260 -24.845 99.265 ;
        RECT -25.275 99.090 -24.385 99.260 ;
        RECT -25.275 99.085 -24.845 99.090 ;
        RECT -27.400 98.770 -26.940 98.795 ;
        RECT -26.590 98.770 -24.810 98.805 ;
        RECT -24.215 98.775 -24.045 99.575 ;
        RECT -24.440 98.770 -24.045 98.775 ;
        RECT -27.400 98.600 -24.045 98.770 ;
        RECT -27.400 98.575 -26.940 98.600 ;
        RECT -26.590 98.570 -24.810 98.600 ;
        RECT -24.440 98.595 -24.045 98.600 ;
        RECT -25.515 98.345 -24.675 98.350 ;
        RECT -25.985 97.980 -24.675 98.345 ;
        RECT -25.985 97.705 -25.635 97.980 ;
        RECT -26.290 97.675 -25.270 97.705 ;
        RECT -26.750 97.505 -24.310 97.675 ;
        RECT -26.290 97.475 -25.270 97.505 ;
        RECT -25.825 96.725 -25.595 97.475 ;
        RECT -26.290 96.695 -25.270 96.725 ;
        RECT -26.750 96.525 -24.310 96.695 ;
        RECT -26.290 96.495 -25.270 96.525 ;
        RECT -25.825 95.745 -25.595 96.495 ;
        RECT -26.290 95.715 -24.330 95.745 ;
        RECT -26.750 95.545 -24.310 95.715 ;
        RECT -26.290 95.515 -24.330 95.545 ;
        RECT -26.040 94.495 -25.670 95.335 ;
        RECT -26.040 94.435 -25.725 94.495 ;
        RECT -25.240 94.440 -24.420 94.725 ;
        RECT -26.760 94.320 -25.725 94.435 ;
        RECT -26.760 94.135 -25.730 94.320 ;
        RECT -24.985 93.955 -24.740 94.440 ;
        RECT -25.985 93.725 -24.740 93.955 ;
        RECT -25.985 93.520 -25.635 93.725 ;
        RECT -26.290 93.490 -25.270 93.520 ;
        RECT -26.750 93.320 -24.310 93.490 ;
        RECT -26.290 93.290 -25.270 93.320 ;
        RECT -25.825 92.540 -25.595 93.290 ;
        RECT -26.290 92.510 -25.270 92.540 ;
        RECT -26.750 92.340 -24.310 92.510 ;
        RECT -26.290 92.310 -25.270 92.340 ;
        RECT -30.980 91.820 -29.960 91.850 ;
        RECT -50.925 91.530 -48.965 91.560 ;
        RECT -51.385 91.360 -48.945 91.530 ;
        RECT -50.925 91.330 -48.965 91.360 ;
        RECT -55.615 91.040 -54.595 91.070 ;
        RECT -56.575 90.870 -54.135 91.040 ;
        RECT -55.615 90.840 -54.595 90.870 ;
        RECT -55.250 90.690 -54.900 90.840 ;
        RECT -55.205 90.515 -55.010 90.690 ;
        RECT -53.220 90.515 -52.535 90.570 ;
        RECT -50.675 90.515 -50.305 91.150 ;
        RECT -30.655 91.070 -30.425 91.820 ;
        RECT -25.825 91.560 -25.595 92.310 ;
        RECT -26.290 91.530 -24.330 91.560 ;
        RECT -26.750 91.360 -24.310 91.530 ;
        RECT -26.290 91.330 -24.330 91.360 ;
        RECT -30.980 91.040 -29.960 91.070 ;
        RECT -31.940 90.870 -29.500 91.040 ;
        RECT -30.980 90.840 -29.960 90.870 ;
        RECT -30.615 90.690 -30.265 90.840 ;
        RECT -55.205 90.310 -50.305 90.515 ;
        RECT -30.570 90.515 -30.375 90.690 ;
        RECT -28.585 90.515 -27.900 90.570 ;
        RECT -26.040 90.515 -25.670 91.150 ;
        RECT -30.570 90.310 -25.670 90.515 ;
        RECT -55.205 90.280 -50.455 90.310 ;
        RECT -30.570 90.280 -25.820 90.310 ;
        RECT -55.195 90.275 -50.455 90.280 ;
        RECT -30.560 90.275 -25.820 90.280 ;
        RECT -53.220 90.270 -52.535 90.275 ;
        RECT -28.585 90.270 -27.900 90.275 ;
        RECT -56.725 85.895 -55.895 86.580 ;
        RECT -57.335 83.400 -56.975 83.520 ;
        RECT -64.370 83.050 -56.975 83.400 ;
        RECT -64.370 81.710 -64.020 83.050 ;
        RECT -57.335 82.995 -56.975 83.050 ;
        RECT -56.460 82.080 -56.245 85.895 ;
        RECT -46.050 85.790 -45.010 86.830 ;
        RECT -57.680 82.040 -56.245 82.080 ;
        RECT -60.650 81.870 -56.245 82.040 ;
        RECT -57.680 81.865 -56.245 81.870 ;
        RECT -64.370 81.540 -63.160 81.710 ;
        RECT -64.855 81.050 -64.315 81.220 ;
        RECT -60.990 80.980 -60.600 81.010 ;
        RECT -57.185 81.005 -56.910 81.695 ;
        RECT -56.460 81.655 -56.245 81.865 ;
        RECT -56.460 81.625 -56.045 81.655 ;
        RECT -56.460 81.455 -54.550 81.625 ;
        RECT -56.460 81.435 -56.045 81.455 ;
        RECT -56.460 81.195 -56.260 81.435 ;
        RECT -48.430 81.095 -47.105 82.435 ;
        RECT -60.990 80.810 -57.610 80.980 ;
        RECT -60.990 80.800 -60.600 80.810 ;
        RECT -63.700 80.560 -63.160 80.730 ;
        RECT -64.855 80.070 -64.315 80.240 ;
        RECT -60.990 80.020 -60.820 80.800 ;
        RECT -57.440 80.790 -56.360 81.005 ;
        RECT -57.440 80.510 -57.245 80.790 ;
        RECT -57.710 80.490 -57.245 80.510 ;
        RECT -60.650 80.320 -57.245 80.490 ;
        RECT -57.710 80.300 -57.245 80.320 ;
        RECT -60.990 80.000 -60.610 80.020 ;
        RECT -57.700 80.000 -57.255 80.025 ;
        RECT -60.990 79.830 -57.255 80.000 ;
        RECT -60.990 79.810 -60.610 79.830 ;
        RECT -57.700 79.815 -57.255 79.830 ;
        RECT -63.700 79.580 -63.160 79.750 ;
        RECT -64.170 78.990 -63.870 79.355 ;
        RECT -64.140 78.685 -63.935 78.990 ;
        RECT -57.435 78.965 -57.255 79.815 ;
        RECT -57.075 79.580 -56.800 80.355 ;
        RECT -57.730 78.945 -57.255 78.965 ;
        RECT -60.650 78.775 -57.255 78.945 ;
        RECT -57.730 78.755 -57.255 78.775 ;
        RECT -65.035 78.630 -63.935 78.685 ;
        RECT -65.075 78.490 -63.935 78.630 ;
        RECT -65.075 78.380 -64.075 78.490 ;
        RECT -67.390 78.005 -65.850 78.175 ;
        RECT -65.665 77.945 -65.310 78.315 ;
        RECT -67.390 77.515 -65.850 77.685 ;
        RECT -67.390 77.025 -65.850 77.195 ;
        RECT -65.635 76.240 -65.440 77.945 ;
        RECT -65.075 77.685 -64.885 78.380 ;
        RECT -59.350 77.905 -59.000 77.935 ;
        RECT -57.025 77.905 -56.845 79.580 ;
        RECT -56.560 79.460 -56.360 80.790 ;
        RECT -56.560 79.435 -56.010 79.460 ;
        RECT -56.560 79.265 -54.550 79.435 ;
        RECT -56.560 79.235 -56.010 79.265 ;
        RECT -56.535 78.230 -56.260 79.005 ;
        RECT -56.490 78.045 -56.320 78.230 ;
        RECT -65.075 77.515 -63.165 77.685 ;
        RECT -59.350 77.555 -56.835 77.905 ;
        RECT -65.075 76.705 -64.885 77.515 ;
        RECT -59.350 76.715 -59.000 77.555 ;
        RECT -65.075 76.535 -63.165 76.705 ;
        RECT -60.210 76.545 -59.000 76.715 ;
        RECT -67.390 76.045 -65.850 76.215 ;
        RECT -65.640 75.890 -65.440 76.240 ;
        RECT -65.640 75.885 -65.430 75.890 ;
        RECT -65.630 73.310 -65.430 75.885 ;
        RECT -65.190 75.620 -64.920 76.295 ;
        RECT -59.055 76.055 -58.515 76.225 ;
        RECT -65.150 75.520 -64.950 75.620 ;
        RECT -60.210 75.565 -59.670 75.735 ;
        RECT -65.140 74.485 -64.960 75.520 ;
        RECT -59.055 75.075 -58.515 75.245 ;
        RECT -60.210 74.585 -59.670 74.755 ;
        RECT -59.500 73.995 -59.200 74.360 ;
        RECT -64.850 73.630 -63.810 73.800 ;
        RECT -59.435 73.690 -59.230 73.995 ;
        RECT -59.435 73.635 -58.335 73.690 ;
        RECT -59.435 73.495 -58.295 73.635 ;
        RECT -59.295 73.385 -58.295 73.495 ;
        RECT -66.500 73.145 -65.430 73.310 ;
        RECT -66.500 73.140 -65.460 73.145 ;
        RECT -64.850 72.650 -63.810 72.820 ;
        RECT -58.485 72.690 -58.295 73.385 ;
        RECT -58.060 72.950 -57.705 73.320 ;
        RECT -57.520 73.010 -55.980 73.180 ;
        RECT -60.205 72.520 -58.295 72.690 ;
        RECT -66.500 72.160 -65.460 72.330 ;
        RECT -64.850 71.670 -63.810 71.840 ;
        RECT -58.485 71.710 -58.295 72.520 ;
        RECT -60.205 71.540 -58.295 71.710 ;
        RECT -65.320 71.080 -65.020 71.445 ;
        RECT -65.290 70.860 -65.085 71.080 ;
        RECT -65.750 70.210 -65.000 70.860 ;
        RECT -58.450 70.625 -58.180 71.300 ;
        RECT -57.930 71.245 -57.735 72.950 ;
        RECT -57.520 72.520 -55.980 72.690 ;
        RECT -57.520 72.030 -55.980 72.200 ;
        RECT -57.930 70.895 -57.730 71.245 ;
        RECT -57.520 71.050 -55.980 71.220 ;
        RECT -57.940 70.890 -57.730 70.895 ;
        RECT -58.420 70.525 -58.220 70.625 ;
        RECT -70.775 68.045 -70.090 68.735 ;
        RECT -71.265 67.355 -70.975 68.040 ;
        RECT -65.455 67.825 -65.115 70.210 ;
        RECT -58.410 68.615 -58.230 70.525 ;
        RECT -57.940 69.760 -57.740 70.890 ;
        RECT -58.770 68.030 -58.155 68.615 ;
        RECT -65.795 67.535 -65.110 67.825 ;
        RECT -71.260 52.805 -71.000 67.355 ;
        RECT -68.240 67.110 -67.555 67.400 ;
        RECT -68.215 59.080 -68.040 67.110 ;
        RECT -57.280 66.800 -56.990 67.410 ;
        RECT -57.280 66.735 -55.830 66.800 ;
        RECT -54.160 66.735 -53.650 66.770 ;
        RECT -57.280 66.565 -53.650 66.735 ;
        RECT -57.280 66.550 -55.830 66.565 ;
        RECT -57.280 66.270 -57.055 66.550 ;
        RECT -54.160 66.540 -53.650 66.565 ;
        RECT -57.280 65.220 -57.100 66.270 ;
        RECT -57.525 65.190 -57.100 65.220 ;
        RECT -58.520 65.020 -57.100 65.190 ;
        RECT -57.525 64.995 -57.100 65.020 ;
        RECT -56.410 66.245 -56.010 66.265 ;
        RECT -56.410 66.075 -54.020 66.245 ;
        RECT -56.410 66.040 -56.010 66.075 ;
        RECT -56.410 64.705 -56.230 66.040 ;
        RECT -53.840 65.780 -53.650 66.540 ;
        RECT -54.160 65.755 -53.650 65.780 ;
        RECT -56.060 65.585 -53.650 65.755 ;
        RECT -54.160 65.550 -53.650 65.585 ;
        RECT -56.410 64.700 -56.035 64.705 ;
        RECT -56.410 64.530 -54.020 64.700 ;
        RECT -56.410 64.525 -56.035 64.530 ;
        RECT -68.225 58.985 -68.040 59.080 ;
        RECT -67.810 62.485 -67.125 62.775 ;
        RECT -68.265 58.310 -67.995 58.985 ;
        RECT -69.500 57.940 -68.095 58.110 ;
        RECT -68.280 57.130 -68.095 57.940 ;
        RECT -67.810 57.305 -67.620 62.485 ;
        RECT -57.275 62.275 -56.985 62.755 ;
        RECT -57.275 62.210 -55.825 62.275 ;
        RECT -54.155 62.210 -53.645 62.245 ;
        RECT -57.275 62.040 -53.645 62.210 ;
        RECT -57.275 62.025 -55.825 62.040 ;
        RECT -57.275 61.745 -57.050 62.025 ;
        RECT -54.155 62.015 -53.645 62.040 ;
        RECT -57.275 60.695 -57.095 61.745 ;
        RECT -57.520 60.665 -57.095 60.695 ;
        RECT -58.515 60.495 -57.095 60.665 ;
        RECT -57.520 60.470 -57.095 60.495 ;
        RECT -56.405 61.720 -56.005 61.740 ;
        RECT -56.405 61.550 -54.015 61.720 ;
        RECT -56.405 61.515 -56.005 61.550 ;
        RECT -56.405 60.180 -56.225 61.515 ;
        RECT -53.835 61.255 -53.645 62.015 ;
        RECT -54.155 61.230 -53.645 61.255 ;
        RECT -56.055 61.060 -53.645 61.230 ;
        RECT -54.155 61.025 -53.645 61.060 ;
        RECT -56.405 60.175 -56.030 60.180 ;
        RECT -56.405 60.005 -54.015 60.175 ;
        RECT -56.405 60.000 -56.030 60.005 ;
        RECT -67.400 58.835 -66.715 59.125 ;
        RECT -69.500 56.960 -68.095 57.130 ;
        RECT -68.280 56.150 -68.095 56.960 ;
        RECT -67.855 56.630 -67.585 57.305 ;
        RECT -67.400 56.365 -67.230 58.835 ;
        RECT -66.950 58.430 -64.925 58.600 ;
        RECT -66.950 57.620 -66.780 58.430 ;
        RECT -59.020 57.890 -58.730 58.320 ;
        RECT -59.020 57.680 -57.600 57.890 ;
        RECT -54.400 57.730 -54.020 57.790 ;
        RECT -59.020 57.635 -58.730 57.680 ;
        RECT -66.950 57.450 -64.925 57.620 ;
        RECT -66.950 56.560 -66.775 57.450 ;
        RECT -66.460 56.880 -64.260 57.050 ;
        RECT -64.965 56.875 -64.260 56.880 ;
        RECT -66.950 56.390 -64.920 56.560 ;
        RECT -66.950 56.385 -66.460 56.390 ;
        RECT -69.500 55.980 -68.095 56.150 ;
        RECT -68.280 55.520 -68.095 55.980 ;
        RECT -67.465 55.690 -67.195 56.365 ;
        RECT -64.445 56.070 -64.260 56.875 ;
        RECT -66.460 55.900 -64.260 56.070 ;
        RECT -64.975 55.895 -64.260 55.900 ;
        RECT -68.280 55.505 -66.780 55.520 ;
        RECT -68.280 55.335 -64.920 55.505 ;
        RECT -67.405 53.310 -67.220 55.335 ;
        RECT -66.950 54.525 -66.780 55.335 ;
        RECT -64.430 55.015 -64.260 55.895 ;
        RECT -59.020 55.635 -58.810 57.635 ;
        RECT -57.810 57.260 -57.600 57.680 ;
        RECT -57.410 57.560 -54.020 57.730 ;
        RECT -54.400 57.510 -54.020 57.560 ;
        RECT -57.810 57.240 -57.320 57.260 ;
        RECT -57.810 57.070 -54.370 57.240 ;
        RECT -57.810 57.050 -57.320 57.070 ;
        RECT -54.190 56.800 -54.020 57.510 ;
        RECT -54.400 56.750 -54.020 56.800 ;
        RECT -57.410 56.580 -54.020 56.750 ;
        RECT -54.400 56.520 -54.020 56.580 ;
        RECT -59.275 55.615 -58.810 55.635 ;
        RECT -60.230 55.445 -58.810 55.615 ;
        RECT -59.275 55.425 -58.810 55.445 ;
        RECT -66.460 54.845 -64.260 55.015 ;
        RECT -59.020 54.655 -58.810 55.425 ;
        RECT -59.275 54.635 -58.810 54.655 ;
        RECT -66.950 54.355 -64.920 54.525 ;
        RECT -60.230 54.465 -58.810 54.635 ;
        RECT -59.275 54.445 -58.810 54.465 ;
        RECT -57.765 56.185 -57.355 56.200 ;
        RECT -57.765 56.015 -54.370 56.185 ;
        RECT -57.765 55.990 -57.355 56.015 ;
        RECT -57.765 55.220 -57.580 55.990 ;
        RECT -54.190 55.740 -54.020 56.520 ;
        RECT -54.400 55.695 -54.020 55.740 ;
        RECT -57.410 55.525 -54.020 55.695 ;
        RECT -54.400 55.475 -54.020 55.525 ;
        RECT -57.765 55.205 -57.360 55.220 ;
        RECT -57.765 55.035 -54.370 55.205 ;
        RECT -57.765 55.010 -57.360 55.035 ;
        RECT -57.765 54.160 -57.580 55.010 ;
        RECT -57.765 54.145 -57.325 54.160 ;
        RECT -57.765 53.975 -54.370 54.145 ;
        RECT -57.765 53.955 -57.325 53.975 ;
        RECT -71.415 52.015 -70.835 52.805 ;
        RECT -67.455 52.635 -67.185 53.310 ;
        RECT -69.500 52.290 -64.920 52.460 ;
        RECT -48.270 38.690 -47.340 81.095 ;
        RECT -46.040 69.140 -45.010 85.790 ;
        RECT -44.170 86.220 -31.245 87.135 ;
        RECT -44.170 82.410 -43.255 86.220 ;
        RECT -32.335 83.400 -31.975 83.520 ;
        RECT -39.370 83.050 -31.975 83.400 ;
        RECT -44.330 81.070 -43.005 82.410 ;
        RECT -39.370 81.710 -39.020 83.050 ;
        RECT -32.335 82.995 -31.975 83.050 ;
        RECT -31.460 82.080 -31.245 86.220 ;
        RECT -32.680 82.040 -31.245 82.080 ;
        RECT -35.650 81.870 -31.245 82.040 ;
        RECT -32.680 81.865 -31.245 81.870 ;
        RECT -39.370 81.540 -38.160 81.710 ;
        RECT -39.855 81.050 -39.315 81.220 ;
        RECT -35.990 80.980 -35.600 81.010 ;
        RECT -32.185 81.005 -31.910 81.695 ;
        RECT -31.460 81.655 -31.245 81.865 ;
        RECT -31.460 81.625 -31.045 81.655 ;
        RECT -31.460 81.455 -29.550 81.625 ;
        RECT -31.460 81.435 -31.045 81.455 ;
        RECT -31.460 81.195 -31.260 81.435 ;
        RECT -35.990 80.810 -32.610 80.980 ;
        RECT -35.990 80.800 -35.600 80.810 ;
        RECT -38.700 80.560 -38.160 80.730 ;
        RECT -39.855 80.070 -39.315 80.240 ;
        RECT -35.990 80.020 -35.820 80.800 ;
        RECT -32.440 80.790 -31.360 81.005 ;
        RECT -32.440 80.510 -32.245 80.790 ;
        RECT -32.710 80.490 -32.245 80.510 ;
        RECT -35.650 80.320 -32.245 80.490 ;
        RECT -32.710 80.300 -32.245 80.320 ;
        RECT -35.990 80.000 -35.610 80.020 ;
        RECT -32.700 80.000 -32.255 80.025 ;
        RECT -35.990 79.830 -32.255 80.000 ;
        RECT -35.990 79.810 -35.610 79.830 ;
        RECT -32.700 79.815 -32.255 79.830 ;
        RECT -38.700 79.580 -38.160 79.750 ;
        RECT -39.170 78.990 -38.870 79.355 ;
        RECT -39.140 78.685 -38.935 78.990 ;
        RECT -32.435 78.965 -32.255 79.815 ;
        RECT -32.075 79.580 -31.800 80.355 ;
        RECT -32.730 78.945 -32.255 78.965 ;
        RECT -35.650 78.775 -32.255 78.945 ;
        RECT -32.730 78.755 -32.255 78.775 ;
        RECT -40.035 78.630 -38.935 78.685 ;
        RECT -40.075 78.490 -38.935 78.630 ;
        RECT -40.075 78.380 -39.075 78.490 ;
        RECT -42.390 78.005 -40.850 78.175 ;
        RECT -40.665 77.945 -40.310 78.315 ;
        RECT -42.390 77.515 -40.850 77.685 ;
        RECT -42.390 77.025 -40.850 77.195 ;
        RECT -40.635 76.240 -40.440 77.945 ;
        RECT -40.075 77.685 -39.885 78.380 ;
        RECT -34.350 77.905 -34.000 77.935 ;
        RECT -32.025 77.905 -31.845 79.580 ;
        RECT -31.560 79.460 -31.360 80.790 ;
        RECT -31.560 79.435 -31.010 79.460 ;
        RECT -31.560 79.265 -29.550 79.435 ;
        RECT -31.560 79.235 -31.010 79.265 ;
        RECT -31.535 78.230 -31.260 79.005 ;
        RECT -31.490 78.045 -31.320 78.230 ;
        RECT -40.075 77.515 -38.165 77.685 ;
        RECT -34.350 77.555 -31.835 77.905 ;
        RECT -40.075 76.705 -39.885 77.515 ;
        RECT -34.350 76.715 -34.000 77.555 ;
        RECT -40.075 76.535 -38.165 76.705 ;
        RECT -35.210 76.545 -34.000 76.715 ;
        RECT -42.390 76.045 -40.850 76.215 ;
        RECT -40.640 75.890 -40.440 76.240 ;
        RECT -40.640 75.885 -40.430 75.890 ;
        RECT -40.630 73.310 -40.430 75.885 ;
        RECT -40.190 75.620 -39.920 76.295 ;
        RECT -34.055 76.055 -33.515 76.225 ;
        RECT -40.150 75.520 -39.950 75.620 ;
        RECT -35.210 75.565 -34.670 75.735 ;
        RECT -40.140 74.485 -39.960 75.520 ;
        RECT -34.055 75.075 -33.515 75.245 ;
        RECT -35.210 74.585 -34.670 74.755 ;
        RECT -34.500 73.995 -34.200 74.360 ;
        RECT -39.850 73.630 -38.810 73.800 ;
        RECT -34.435 73.690 -34.230 73.995 ;
        RECT -34.435 73.635 -33.335 73.690 ;
        RECT -34.435 73.495 -33.295 73.635 ;
        RECT -34.295 73.385 -33.295 73.495 ;
        RECT -41.500 73.145 -40.430 73.310 ;
        RECT -41.500 73.140 -40.460 73.145 ;
        RECT -39.850 72.650 -38.810 72.820 ;
        RECT -33.485 72.690 -33.295 73.385 ;
        RECT -33.060 72.950 -32.705 73.320 ;
        RECT -32.520 73.010 -30.980 73.180 ;
        RECT -35.205 72.520 -33.295 72.690 ;
        RECT -41.500 72.160 -40.460 72.330 ;
        RECT -39.850 71.670 -38.810 71.840 ;
        RECT -33.485 71.710 -33.295 72.520 ;
        RECT -35.205 71.540 -33.295 71.710 ;
        RECT -40.320 71.080 -40.020 71.445 ;
        RECT -32.930 71.245 -32.735 72.950 ;
        RECT -32.520 72.520 -30.980 72.690 ;
        RECT -32.520 72.030 -30.980 72.200 ;
        RECT -40.290 70.860 -40.085 71.080 ;
        RECT -32.930 70.895 -32.730 71.245 ;
        RECT -32.520 71.050 -30.980 71.220 ;
        RECT -32.940 70.890 -32.730 70.895 ;
        RECT -40.750 70.210 -40.000 70.860 ;
        RECT -40.500 68.335 -40.330 70.210 ;
        RECT -32.940 69.760 -32.740 70.890 ;
        RECT -30.005 70.385 -29.715 70.705 ;
        RECT -30.060 68.535 -29.710 70.385 ;
        RECT -30.060 68.365 -28.850 68.535 ;
        RECT -42.505 68.165 -37.925 68.335 ;
        RECT -40.240 67.315 -39.970 67.990 ;
        RECT -30.545 67.875 -30.005 68.045 ;
        RECT -29.390 67.385 -28.850 67.555 ;
        RECT -42.505 66.100 -40.475 66.270 ;
        RECT -43.165 65.610 -40.965 65.780 ;
        RECT -43.165 64.730 -42.995 65.610 ;
        RECT -40.645 65.290 -40.475 66.100 ;
        RECT -40.205 65.290 -40.020 67.315 ;
        RECT -30.545 66.895 -30.005 67.065 ;
        RECT -29.390 66.405 -28.850 66.575 ;
        RECT -29.860 65.815 -29.560 66.180 ;
        RECT -29.830 65.510 -29.625 65.815 ;
        RECT -30.725 65.455 -29.625 65.510 ;
        RECT -30.765 65.315 -29.625 65.455 ;
        RECT -42.505 65.120 -39.145 65.290 ;
        RECT -40.645 65.105 -39.145 65.120 ;
        RECT -43.165 64.725 -42.450 64.730 ;
        RECT -43.165 64.555 -40.965 64.725 ;
        RECT -43.165 63.750 -42.980 64.555 ;
        RECT -40.230 64.260 -39.960 64.935 ;
        RECT -39.330 64.645 -39.145 65.105 ;
        RECT -30.765 65.205 -29.765 65.315 ;
        RECT -33.080 64.830 -31.540 65.000 ;
        RECT -39.330 64.475 -37.925 64.645 ;
        RECT -30.765 64.510 -30.575 65.205 ;
        RECT -40.965 64.235 -40.475 64.240 ;
        RECT -42.505 64.065 -40.475 64.235 ;
        RECT -43.165 63.745 -42.460 63.750 ;
        RECT -43.165 63.575 -40.965 63.745 ;
        RECT -40.650 63.175 -40.475 64.065 ;
        RECT -42.500 63.005 -40.475 63.175 ;
        RECT -40.645 62.195 -40.475 63.005 ;
        RECT -42.500 62.025 -40.475 62.195 ;
        RECT -40.195 61.725 -40.025 64.260 ;
        RECT -39.840 63.320 -39.570 63.995 ;
        RECT -39.330 63.665 -39.145 64.475 ;
        RECT -33.080 64.340 -31.540 64.510 ;
        RECT -30.765 64.340 -28.855 64.510 ;
        RECT -33.080 63.850 -31.540 64.020 ;
        RECT -39.330 63.495 -37.925 63.665 ;
        RECT -30.765 63.530 -30.575 64.340 ;
        RECT -40.900 61.555 -40.025 61.725 ;
        RECT -40.900 60.870 -40.730 61.555 ;
        RECT -39.805 61.355 -39.615 63.320 ;
        RECT -39.330 62.685 -39.145 63.495 ;
        RECT -30.765 63.360 -28.855 63.530 ;
        RECT -33.080 62.870 -31.540 63.040 ;
        RECT -39.330 62.515 -37.925 62.685 ;
        RECT -39.430 61.640 -39.160 62.315 ;
        RECT 469.655 62.300 475.760 192.475 ;
        RECT -39.385 61.545 -39.200 61.640 ;
        RECT -40.260 61.065 -39.575 61.355 ;
        RECT -39.805 60.935 -39.615 61.065 ;
        RECT -40.915 60.580 -40.230 60.870 ;
        RECT -39.375 60.045 -39.200 61.545 ;
        RECT -39.605 59.840 -39.200 60.045 ;
        RECT -41.400 59.510 -40.715 59.800 ;
        RECT -39.605 58.825 -39.255 59.840 ;
        RECT -32.825 59.015 -28.245 59.185 ;
        RECT -39.605 58.655 -38.395 58.825 ;
        RECT -40.090 58.165 -39.550 58.335 ;
        RECT -30.560 58.165 -30.290 58.840 ;
        RECT -38.935 57.675 -38.395 57.845 ;
        RECT -40.090 57.185 -39.550 57.355 ;
        RECT -32.825 56.950 -30.795 57.120 ;
        RECT -38.935 56.695 -38.395 56.865 ;
        RECT -39.405 56.105 -39.105 56.470 ;
        RECT -33.485 56.460 -31.285 56.630 ;
        RECT -39.375 55.800 -39.170 56.105 ;
        RECT -40.270 55.745 -39.170 55.800 ;
        RECT -40.310 55.605 -39.170 55.745 ;
        RECT -40.310 55.495 -39.310 55.605 ;
        RECT -33.485 55.580 -33.315 56.460 ;
        RECT -30.965 56.140 -30.795 56.950 ;
        RECT -30.525 56.140 -30.340 58.165 ;
        RECT -32.825 55.970 -29.465 56.140 ;
        RECT -30.965 55.955 -29.465 55.970 ;
        RECT -33.485 55.575 -32.770 55.580 ;
        RECT -42.625 55.120 -41.085 55.290 ;
        RECT -40.310 54.800 -40.120 55.495 ;
        RECT -33.485 55.405 -31.285 55.575 ;
        RECT -29.650 55.495 -29.465 55.955 ;
        RECT -42.625 54.630 -41.085 54.800 ;
        RECT -40.310 54.630 -38.400 54.800 ;
        RECT -42.625 54.140 -41.085 54.310 ;
        RECT -40.310 53.820 -40.120 54.630 ;
        RECT -33.485 54.600 -33.300 55.405 ;
        RECT -29.650 55.325 -28.245 55.495 ;
        RECT -31.285 55.085 -30.795 55.090 ;
        RECT -32.825 54.915 -30.795 55.085 ;
        RECT -33.485 54.595 -32.780 54.600 ;
        RECT -33.485 54.425 -31.285 54.595 ;
        RECT -30.970 54.025 -30.795 54.915 ;
        RECT -32.820 53.855 -30.795 54.025 ;
        RECT -40.310 53.650 -38.400 53.820 ;
        RECT -42.625 53.160 -41.085 53.330 ;
        RECT -30.965 53.045 -30.795 53.855 ;
        RECT -29.650 54.515 -29.465 55.325 ;
        RECT -29.650 54.345 -28.245 54.515 ;
        RECT -29.650 53.535 -29.465 54.345 ;
        RECT -0.585 54.035 0.365 61.985 ;
        RECT -29.650 53.365 -28.245 53.535 ;
        RECT -32.820 52.875 -30.795 53.045 ;
        RECT 73.905 50.665 75.465 50.835 ;
        RECT 75.920 50.665 76.960 50.835 ;
        RECT 82.070 50.690 83.110 50.860 ;
        RECT 75.295 50.440 75.465 50.665 ;
        RECT 75.220 50.035 75.595 50.440 ;
        RECT 81.410 49.990 81.800 50.355 ;
        RECT 75.920 49.375 78.960 49.545 ;
        RECT 79.580 49.400 81.110 49.570 ;
        RECT 75.200 48.255 75.575 48.370 ;
        RECT 73.905 48.085 75.575 48.255 ;
        RECT 75.920 48.085 76.960 48.255 ;
        RECT 75.200 47.965 75.575 48.085 ;
        RECT 77.185 46.965 77.710 49.375 ;
        RECT 79.580 46.990 79.750 49.400 ;
        RECT 81.535 48.950 81.705 49.990 ;
        RECT 82.070 49.400 85.110 49.570 ;
        RECT 81.415 48.585 81.805 48.950 ;
        RECT 81.535 47.545 81.705 48.585 ;
        RECT 82.070 48.110 83.110 48.280 ;
        RECT 81.440 47.180 81.830 47.545 ;
        RECT 81.535 46.990 81.705 47.180 ;
        RECT 83.345 46.990 83.515 49.400 ;
        RECT 346.870 48.890 349.030 49.580 ;
        RECT 458.870 48.890 461.030 49.580 ;
        RECT 75.920 46.795 78.960 46.965 ;
        RECT 79.580 46.820 81.705 46.990 ;
        RECT 82.070 46.820 85.110 46.990 ;
        RECT 75.090 45.735 75.440 46.090 ;
        RECT 77.470 46.030 77.805 46.365 ;
        RECT 75.090 45.675 75.355 45.735 ;
        RECT 73.905 45.505 75.355 45.675 ;
        RECT 75.920 45.505 76.960 45.675 ;
        RECT 74.940 45.500 75.355 45.505 ;
        RECT 72.930 44.085 73.865 44.495 ;
        RECT 75.090 44.085 75.355 45.500 ;
        RECT 77.520 44.440 77.690 46.030 ;
        RECT 77.520 44.270 79.450 44.440 ;
        RECT 79.635 44.165 79.975 44.485 ;
        RECT 80.145 44.270 80.605 44.440 ;
        RECT 72.930 43.820 75.355 44.085 ;
        RECT 34.830 43.455 36.560 43.780 ;
        RECT 72.930 43.730 73.865 43.820 ;
        RECT 75.090 43.695 75.355 43.820 ;
        RECT 79.710 43.455 79.890 44.165 ;
        RECT 81.520 43.715 81.690 46.820 ;
        RECT 83.580 46.040 83.920 46.370 ;
        RECT 82.070 45.530 83.110 45.700 ;
        RECT 34.830 42.650 80.025 43.455 ;
        RECT 81.130 43.025 81.980 43.715 ;
        RECT 34.830 42.330 36.560 42.650 ;
        RECT 36.445 41.305 38.175 41.535 ;
        RECT 83.610 41.305 83.875 46.040 ;
        RECT 36.445 40.395 83.995 41.305 ;
        RECT 36.445 40.085 38.175 40.395 ;
        RECT -68.545 37.760 -47.340 38.690 ;
        RECT -68.545 13.425 -67.615 37.760 ;
        RECT 45.010 32.790 45.180 37.500 ;
        RECT 46.170 32.790 46.750 33.070 ;
        RECT 47.670 32.790 48.250 33.070 ;
        RECT 49.170 32.790 49.750 33.070 ;
        RECT 50.670 32.790 51.250 33.070 ;
        RECT 52.170 32.790 52.750 33.070 ;
        RECT 53.590 32.790 53.760 37.500 ;
        RECT 60.820 32.810 60.990 37.500 ;
        RECT 74.985 34.655 76.055 34.850 ;
        RECT 96.005 34.655 98.215 35.425 ;
        RECT 114.695 34.655 116.515 35.580 ;
        RECT 74.985 34.035 116.515 34.655 ;
        RECT 74.985 33.780 76.055 34.035 ;
        RECT 81.135 32.810 82.030 33.115 ;
        RECT 96.005 33.100 98.215 34.035 ;
        RECT 114.695 33.330 116.515 34.035 ;
        RECT 45.010 32.620 53.940 32.790 ;
        RECT 45.190 28.195 45.360 32.620 ;
        RECT 53.770 28.195 53.940 32.620 ;
        RECT 60.820 32.400 82.030 32.810 ;
        RECT 81.135 32.220 82.030 32.400 ;
        RECT 69.330 29.490 70.650 29.820 ;
        RECT 62.325 28.205 70.650 29.490 ;
        RECT 62.350 23.195 62.520 28.205 ;
        RECT 93.955 26.080 95.840 27.865 ;
        RECT 106.680 17.255 107.520 17.455 ;
        RECT 106.050 17.085 107.520 17.255 ;
        RECT 99.460 16.890 99.630 16.910 ;
        RECT 99.430 15.625 99.660 16.890 ;
        RECT 100.440 15.950 100.610 16.910 ;
        RECT 101.420 15.950 101.590 16.910 ;
        RECT 103.710 16.890 103.880 16.910 ;
        RECT 100.410 15.625 100.640 15.950 ;
        RECT 101.390 15.625 101.620 15.950 ;
        RECT 99.430 15.585 101.620 15.625 ;
        RECT 103.680 15.625 103.910 16.890 ;
        RECT 104.690 15.950 104.860 16.910 ;
        RECT 105.670 15.950 105.840 16.910 ;
        RECT 104.660 15.625 104.890 15.950 ;
        RECT 105.640 15.625 105.870 15.950 ;
        RECT 103.680 15.585 105.870 15.625 ;
        RECT 106.050 15.585 106.220 17.085 ;
        RECT 99.430 15.510 102.450 15.585 ;
        RECT 102.660 15.510 103.500 15.550 ;
        RECT 99.430 15.395 103.500 15.510 ;
        RECT 99.430 14.930 99.660 15.395 ;
        RECT 100.410 14.930 100.640 15.395 ;
        RECT 101.390 15.250 103.500 15.395 ;
        RECT 101.390 15.235 102.450 15.250 ;
        RECT 101.390 14.930 101.620 15.235 ;
        RECT 102.660 15.180 103.500 15.250 ;
        RECT 103.680 15.395 106.220 15.585 ;
        RECT 103.680 14.930 103.910 15.395 ;
        RECT 104.660 14.930 104.890 15.395 ;
        RECT 105.640 15.235 106.220 15.395 ;
        RECT 106.450 15.625 106.620 16.910 ;
        RECT 106.940 15.870 107.110 16.910 ;
        RECT 107.430 15.625 107.600 16.910 ;
        RECT 107.920 15.870 108.090 16.910 ;
        RECT 108.410 15.625 108.580 16.910 ;
        RECT 108.900 15.870 109.070 16.910 ;
        RECT 109.390 15.625 109.560 16.910 ;
        RECT 109.880 15.870 110.050 16.910 ;
        RECT 110.370 15.625 110.540 16.910 ;
        RECT 106.450 15.455 110.540 15.625 ;
        RECT 105.640 14.930 105.870 15.235 ;
        RECT 99.460 14.470 99.630 14.930 ;
        RECT 100.440 14.470 100.610 14.930 ;
        RECT 101.420 14.470 101.590 14.930 ;
        RECT 103.710 14.470 103.880 14.930 ;
        RECT 104.690 14.470 104.860 14.930 ;
        RECT 105.670 14.470 105.840 14.930 ;
        RECT 106.450 14.140 106.620 15.455 ;
        RECT 106.940 14.140 107.110 15.180 ;
        RECT 107.430 14.140 107.600 15.455 ;
        RECT 107.920 14.140 108.090 15.180 ;
        RECT 108.410 14.140 108.580 15.455 ;
        RECT 108.900 14.140 109.070 15.180 ;
        RECT 109.390 14.140 109.560 15.455 ;
        RECT 109.880 14.140 110.050 15.180 ;
        RECT 110.370 14.140 110.540 15.455 ;
        RECT 203.880 14.790 207.020 14.960 ;
        RECT 196.420 14.675 196.590 14.695 ;
        RECT -29.225 13.425 -27.695 13.820 ;
        RECT 111.580 13.555 112.770 14.500 ;
        RECT -68.545 12.740 -27.695 13.425 ;
        RECT -29.225 12.415 -27.695 12.740 ;
        RECT 1.310 12.710 5.555 12.975 ;
        RECT -10.210 10.550 -9.370 10.750 ;
        RECT -10.840 10.380 -9.370 10.550 ;
        RECT -17.430 10.185 -17.260 10.205 ;
        RECT -48.655 6.855 -48.295 7.125 ;
        RECT -46.925 6.855 -46.755 9.895 ;
        RECT -45.745 7.855 -45.575 9.895 ;
        RECT -44.565 7.855 -44.395 9.895 ;
        RECT -43.385 7.855 -43.215 9.895 ;
        RECT -42.205 7.855 -42.035 9.895 ;
        RECT -41.025 7.855 -40.855 9.895 ;
        RECT -39.845 7.855 -39.675 9.895 ;
        RECT -38.665 7.855 -38.495 9.895 ;
        RECT -48.655 6.685 -46.755 6.855 ;
        RECT -39.215 6.925 -38.855 7.295 ;
        RECT -36.835 6.925 -36.665 9.895 ;
        RECT -35.655 7.855 -35.485 9.895 ;
        RECT -34.475 7.855 -34.305 9.895 ;
        RECT -33.295 7.855 -33.125 9.895 ;
        RECT -31.465 7.525 -31.295 9.895 ;
        RECT -30.285 7.855 -30.115 9.895 ;
        RECT -17.460 8.920 -17.230 10.185 ;
        RECT -16.450 9.245 -16.280 10.205 ;
        RECT -15.470 9.245 -15.300 10.205 ;
        RECT -13.180 10.185 -13.010 10.205 ;
        RECT -16.480 8.920 -16.250 9.245 ;
        RECT -15.500 8.920 -15.270 9.245 ;
        RECT -17.460 8.880 -15.270 8.920 ;
        RECT -13.210 8.920 -12.980 10.185 ;
        RECT -12.200 9.245 -12.030 10.205 ;
        RECT -11.220 9.245 -11.050 10.205 ;
        RECT -12.230 8.920 -12.000 9.245 ;
        RECT -11.250 8.920 -11.020 9.245 ;
        RECT -13.210 8.880 -11.020 8.920 ;
        RECT -10.840 8.880 -10.670 10.380 ;
        RECT -17.460 8.805 -14.440 8.880 ;
        RECT -14.230 8.805 -13.390 8.845 ;
        RECT -17.460 8.690 -13.390 8.805 ;
        RECT -28.210 7.570 -27.870 7.605 ;
        RECT -32.335 7.355 -31.295 7.525 ;
        RECT -39.215 6.755 -36.665 6.925 ;
        RECT -34.560 6.910 -34.050 7.150 ;
        RECT -32.335 6.910 -32.165 7.355 ;
        RECT -48.655 6.345 -48.295 6.685 ;
        RECT -39.215 6.515 -38.855 6.755 ;
        RECT -34.560 6.740 -32.165 6.910 ;
        RECT -31.550 6.760 -31.170 7.060 ;
        RECT -28.895 6.760 -27.870 7.570 ;
        RECT -21.060 7.305 -20.495 7.675 ;
        RECT -17.920 7.510 -17.750 8.305 ;
        RECT -17.460 8.225 -17.230 8.690 ;
        RECT -17.430 7.765 -17.260 8.225 ;
        RECT -16.940 7.510 -16.770 8.305 ;
        RECT -16.480 8.225 -16.250 8.690 ;
        RECT -15.500 8.545 -13.390 8.690 ;
        RECT -15.500 8.530 -14.440 8.545 ;
        RECT -16.450 7.765 -16.280 8.225 ;
        RECT -15.960 7.510 -15.790 8.305 ;
        RECT -15.500 8.225 -15.270 8.530 ;
        RECT -14.230 8.475 -13.390 8.545 ;
        RECT -13.210 8.690 -10.670 8.880 ;
        RECT -15.470 7.765 -15.300 8.225 ;
        RECT -13.670 7.510 -13.500 8.305 ;
        RECT -13.210 8.225 -12.980 8.690 ;
        RECT -13.180 7.765 -13.010 8.225 ;
        RECT -12.690 7.510 -12.520 8.305 ;
        RECT -12.230 8.225 -12.000 8.690 ;
        RECT -11.250 8.530 -10.670 8.690 ;
        RECT -10.440 8.920 -10.270 10.205 ;
        RECT -9.950 9.165 -9.780 10.205 ;
        RECT -9.460 8.920 -9.290 10.205 ;
        RECT -8.970 9.165 -8.800 10.205 ;
        RECT -8.480 8.920 -8.310 10.205 ;
        RECT -7.990 9.165 -7.820 10.205 ;
        RECT -7.500 8.920 -7.330 10.205 ;
        RECT -7.010 9.165 -6.840 10.205 ;
        RECT -6.520 8.920 -6.350 10.205 ;
        RECT -10.440 8.750 -6.350 8.920 ;
        RECT -12.200 7.765 -12.030 8.225 ;
        RECT -11.710 7.510 -11.540 8.305 ;
        RECT -11.250 8.225 -11.020 8.530 ;
        RECT -11.220 7.765 -11.050 8.225 ;
        RECT -34.560 6.450 -34.050 6.740 ;
        RECT -31.550 6.495 -28.210 6.760 ;
        RECT -31.550 6.455 -28.505 6.495 ;
        RECT -66.685 6.175 -49.275 6.315 ;
        RECT -31.550 6.175 -31.170 6.455 ;
        RECT -66.685 5.855 -48.535 6.175 ;
        RECT -66.555 3.815 -66.385 5.855 ;
        RECT -65.965 3.815 -65.795 5.855 ;
        RECT -65.375 3.815 -65.205 5.855 ;
        RECT -64.785 3.815 -64.615 5.855 ;
        RECT -64.195 3.815 -64.025 5.855 ;
        RECT -63.605 3.815 -63.435 5.855 ;
        RECT -63.015 3.815 -62.845 5.855 ;
        RECT -62.425 3.815 -62.255 5.855 ;
        RECT -61.835 3.815 -61.665 5.855 ;
        RECT -61.245 3.815 -61.075 5.855 ;
        RECT -60.655 3.815 -60.485 5.855 ;
        RECT -60.065 3.815 -59.895 5.855 ;
        RECT -59.475 3.815 -59.305 5.855 ;
        RECT -58.885 3.815 -58.715 5.855 ;
        RECT -58.295 3.815 -58.125 5.855 ;
        RECT -57.705 3.815 -57.535 5.855 ;
        RECT -57.115 3.815 -56.945 5.855 ;
        RECT -56.525 3.815 -56.355 5.855 ;
        RECT -55.935 3.815 -55.765 5.855 ;
        RECT -55.345 3.815 -55.175 5.855 ;
        RECT -54.755 3.815 -54.585 5.855 ;
        RECT -54.165 3.815 -53.995 5.855 ;
        RECT -53.575 3.815 -53.405 5.855 ;
        RECT -52.985 3.815 -52.815 5.855 ;
        RECT -52.395 3.815 -52.225 5.855 ;
        RECT -51.805 3.815 -51.635 5.855 ;
        RECT -51.215 3.815 -51.045 5.855 ;
        RECT -50.625 3.815 -50.455 5.855 ;
        RECT -50.035 3.815 -49.865 5.855 ;
        RECT -49.445 3.815 -49.275 5.855 ;
        RECT -48.855 3.460 -48.685 5.855 ;
        RECT -47.675 3.460 -47.505 5.855 ;
        RECT -46.495 3.460 -46.325 5.855 ;
        RECT -45.315 3.460 -45.145 5.855 ;
        RECT -44.135 3.460 -43.965 5.855 ;
        RECT -42.955 3.460 -42.785 5.855 ;
        RECT -41.775 3.460 -41.605 5.855 ;
        RECT -40.595 3.460 -40.425 5.855 ;
        RECT -39.415 3.460 -39.245 5.855 ;
        RECT -38.825 3.815 -38.655 5.855 ;
        RECT -38.235 3.460 -38.065 5.855 ;
        RECT -37.645 3.815 -37.475 5.855 ;
        RECT -37.055 3.460 -36.885 5.855 ;
        RECT -36.465 3.815 -36.295 5.855 ;
        RECT -35.875 3.460 -35.705 5.855 ;
        RECT -35.285 3.815 -35.115 5.855 ;
        RECT -34.695 3.460 -34.525 5.855 ;
        RECT -34.105 3.815 -33.935 5.855 ;
        RECT -33.515 3.460 -33.345 5.855 ;
        RECT -32.925 3.815 -32.755 5.855 ;
        RECT -32.335 3.460 -32.165 5.855 ;
        RECT -31.745 3.815 -31.575 5.855 ;
        RECT -31.155 3.460 -30.985 5.855 ;
        RECT -66.605 3.400 -30.875 3.460 ;
        RECT -20.935 3.400 -20.510 7.305 ;
        RECT -17.965 7.170 -11.045 7.510 ;
        RECT -10.440 7.435 -10.270 8.750 ;
        RECT -9.950 7.435 -9.780 8.475 ;
        RECT -9.460 7.435 -9.290 8.750 ;
        RECT -8.970 7.435 -8.800 8.475 ;
        RECT -8.480 7.435 -8.310 8.750 ;
        RECT -7.990 7.435 -7.820 8.475 ;
        RECT -7.500 7.435 -7.330 8.750 ;
        RECT -7.010 7.435 -6.840 8.475 ;
        RECT -6.520 7.435 -6.350 8.750 ;
        RECT -13.715 6.485 -11.045 7.170 ;
        RECT -13.670 5.690 -13.500 6.485 ;
        RECT -13.180 5.770 -13.010 6.230 ;
        RECT -13.210 5.305 -12.980 5.770 ;
        RECT -12.690 5.690 -12.520 6.485 ;
        RECT -12.200 5.770 -12.030 6.230 ;
        RECT -12.230 5.305 -12.000 5.770 ;
        RECT -11.710 5.690 -11.540 6.485 ;
        RECT -11.220 5.770 -11.050 6.230 ;
        RECT -11.250 5.465 -11.020 5.770 ;
        RECT -9.950 5.520 -9.780 6.560 ;
        RECT -8.970 5.520 -8.800 6.560 ;
        RECT -7.990 5.520 -7.820 6.560 ;
        RECT -7.010 5.520 -6.840 6.560 ;
        RECT -11.250 5.305 -10.670 5.465 ;
        RECT -13.210 5.115 -10.670 5.305 ;
        RECT -13.210 5.075 -11.020 5.115 ;
        RECT -13.210 3.810 -12.980 5.075 ;
        RECT -12.230 4.750 -12.000 5.075 ;
        RECT -11.250 4.750 -11.020 5.075 ;
        RECT -13.180 3.790 -13.010 3.810 ;
        RECT -12.200 3.790 -12.030 4.750 ;
        RECT -11.220 3.790 -11.050 4.750 ;
        RECT -10.840 3.615 -10.670 5.115 ;
        RECT 1.310 4.890 1.575 12.710 ;
        RECT 5.170 12.505 5.555 12.710 ;
        RECT 3.690 12.335 4.875 12.485 ;
        RECT 2.345 12.140 4.875 12.335 ;
        RECT 2.345 9.615 2.540 12.140 ;
        RECT 3.690 12.005 4.875 12.140 ;
        RECT 5.170 12.025 10.060 12.505 ;
        RECT 103.710 12.475 103.880 12.935 ;
        RECT 104.690 12.475 104.860 12.935 ;
        RECT 105.670 12.475 105.840 12.935 ;
        RECT 103.680 12.010 103.910 12.475 ;
        RECT 104.660 12.010 104.890 12.475 ;
        RECT 105.640 12.170 105.870 12.475 ;
        RECT 106.940 12.225 107.110 13.265 ;
        RECT 107.920 12.225 108.090 13.265 ;
        RECT 108.900 12.225 109.070 13.265 ;
        RECT 109.880 12.225 110.050 13.265 ;
        RECT 105.640 12.010 106.220 12.170 ;
        RECT 103.680 11.820 106.220 12.010 ;
        RECT 103.680 11.780 105.870 11.820 ;
        RECT 30.285 11.430 31.125 11.630 ;
        RECT 29.655 11.260 31.125 11.430 ;
        RECT 4.475 10.740 4.875 11.110 ;
        RECT 5.130 10.740 5.520 11.105 ;
        RECT 6.830 10.740 7.220 11.110 ;
        RECT 8.000 11.075 8.395 11.170 ;
        RECT 8.000 10.865 8.970 11.075 ;
        RECT 8.000 10.770 8.395 10.865 ;
        RECT 3.125 9.615 3.295 10.445 ;
        RECT 4.355 9.930 4.525 10.570 ;
        RECT 4.945 9.930 5.115 10.570 ;
        RECT 5.535 9.930 5.705 10.570 ;
        RECT 6.565 9.930 6.735 10.570 ;
        RECT 2.325 9.420 3.295 9.615 ;
        RECT 3.125 8.245 3.295 9.420 ;
        RECT 3.465 9.660 3.865 9.750 ;
        RECT 7.005 9.660 7.175 10.570 ;
        RECT 8.015 9.955 8.185 10.595 ;
        RECT 8.455 9.955 8.625 10.595 ;
        RECT 3.465 9.420 7.955 9.660 ;
        RECT 8.795 9.620 8.970 10.865 ;
        RECT 9.260 10.800 11.425 11.190 ;
        RECT 23.065 11.065 23.235 11.085 ;
        RECT 9.145 9.990 9.315 10.630 ;
        RECT 9.290 9.620 10.095 9.785 ;
        RECT 3.465 9.295 4.300 9.420 ;
        RECT 3.885 9.270 4.300 9.295 ;
        RECT 4.805 8.475 4.975 9.115 ;
        RECT 5.685 8.475 5.855 9.420 ;
        RECT 6.565 8.475 6.735 9.420 ;
        RECT 7.155 9.285 7.955 9.420 ;
        RECT 8.175 9.285 8.585 9.615 ;
        RECT 8.795 9.445 10.095 9.620 ;
        RECT 9.290 9.285 10.095 9.445 ;
        RECT 10.325 9.625 10.495 10.630 ;
        RECT 11.505 9.625 11.675 10.630 ;
        RECT 12.370 9.660 12.770 9.750 ;
        RECT 11.935 9.625 12.770 9.660 ;
        RECT 10.325 9.455 12.770 9.625 ;
        RECT 5.585 7.870 5.945 8.275 ;
        RECT 6.470 7.865 6.830 8.270 ;
        RECT 7.570 8.175 7.740 9.285 ;
        RECT 8.010 8.175 8.180 9.115 ;
        RECT 9.770 9.110 9.940 9.115 ;
        RECT 10.325 9.110 10.495 9.455 ;
        RECT 11.935 9.295 12.770 9.455 ;
        RECT 12.940 9.660 13.110 10.445 ;
        RECT 13.915 9.660 14.315 9.750 ;
        RECT 12.940 9.420 14.315 9.660 ;
        RECT 11.935 9.270 12.350 9.295 ;
        RECT 9.770 8.925 10.495 9.110 ;
        RECT 9.770 8.310 9.940 8.925 ;
        RECT 10.325 8.310 10.495 8.925 ;
        RECT 9.770 8.125 10.495 8.310 ;
        RECT 12.940 8.245 13.110 9.420 ;
        RECT 13.480 9.295 14.315 9.420 ;
        RECT 14.485 9.615 14.655 10.445 ;
        RECT 23.035 9.800 23.265 11.065 ;
        RECT 24.045 10.125 24.215 11.085 ;
        RECT 25.025 10.125 25.195 11.085 ;
        RECT 27.315 11.065 27.485 11.085 ;
        RECT 24.015 9.800 24.245 10.125 ;
        RECT 24.995 9.800 25.225 10.125 ;
        RECT 23.035 9.760 25.225 9.800 ;
        RECT 27.285 9.800 27.515 11.065 ;
        RECT 28.295 10.125 28.465 11.085 ;
        RECT 29.275 10.125 29.445 11.085 ;
        RECT 28.265 9.800 28.495 10.125 ;
        RECT 29.245 9.800 29.475 10.125 ;
        RECT 27.285 9.760 29.475 9.800 ;
        RECT 29.655 9.760 29.825 11.260 ;
        RECT 23.035 9.685 26.055 9.760 ;
        RECT 26.265 9.685 27.105 9.725 ;
        RECT 14.485 9.420 20.365 9.615 ;
        RECT 13.480 9.270 13.895 9.295 ;
        RECT 14.485 8.245 14.655 9.420 ;
        RECT 20.170 8.190 20.365 9.420 ;
        RECT 23.035 9.570 27.105 9.685 ;
        RECT 23.035 9.105 23.265 9.570 ;
        RECT 24.015 9.105 24.245 9.570 ;
        RECT 24.995 9.425 27.105 9.570 ;
        RECT 24.995 9.410 26.055 9.425 ;
        RECT 24.995 9.105 25.225 9.410 ;
        RECT 26.265 9.355 27.105 9.425 ;
        RECT 27.285 9.570 29.825 9.760 ;
        RECT 27.285 9.105 27.515 9.570 ;
        RECT 28.265 9.105 28.495 9.570 ;
        RECT 29.245 9.410 29.825 9.570 ;
        RECT 30.055 9.800 30.225 11.085 ;
        RECT 30.545 10.045 30.715 11.085 ;
        RECT 31.035 9.800 31.205 11.085 ;
        RECT 31.525 10.045 31.695 11.085 ;
        RECT 32.015 9.800 32.185 11.085 ;
        RECT 32.505 10.045 32.675 11.085 ;
        RECT 32.995 9.800 33.165 11.085 ;
        RECT 33.485 10.045 33.655 11.085 ;
        RECT 33.975 9.800 34.145 11.085 ;
        RECT 30.055 9.630 34.145 9.800 ;
        RECT 29.245 9.105 29.475 9.410 ;
        RECT 23.065 8.645 23.235 9.105 ;
        RECT 24.045 8.645 24.215 9.105 ;
        RECT 25.025 8.645 25.195 9.105 ;
        RECT 27.315 8.645 27.485 9.105 ;
        RECT 28.295 8.645 28.465 9.105 ;
        RECT 29.275 8.645 29.445 9.105 ;
        RECT 30.055 8.315 30.225 9.630 ;
        RECT 30.545 8.315 30.715 9.355 ;
        RECT 31.035 8.315 31.205 9.630 ;
        RECT 31.525 8.315 31.695 9.355 ;
        RECT 32.015 8.315 32.185 9.630 ;
        RECT 32.505 8.315 32.675 9.355 ;
        RECT 32.995 8.315 33.165 9.630 ;
        RECT 33.485 8.315 33.655 9.355 ;
        RECT 33.975 8.315 34.145 9.630 ;
        RECT 35.270 9.225 36.515 10.395 ;
        RECT 38.680 9.265 38.850 11.305 ;
        RECT 19.950 7.495 20.530 8.190 ;
        RECT 35.480 7.840 36.170 9.225 ;
        RECT 39.860 8.935 40.030 11.305 ;
        RECT 41.690 9.265 41.860 11.305 ;
        RECT 42.870 9.265 43.040 11.305 ;
        RECT 44.050 9.265 44.220 11.305 ;
        RECT 39.860 8.765 40.900 8.935 ;
        RECT 36.685 8.170 37.350 8.400 ;
        RECT 39.735 8.170 40.115 8.470 ;
        RECT 36.685 7.865 40.115 8.170 ;
        RECT 40.730 8.320 40.900 8.765 ;
        RECT 42.615 8.320 43.125 8.560 ;
        RECT 40.730 8.150 43.125 8.320 ;
        RECT 45.230 8.335 45.400 11.305 ;
        RECT 47.060 9.265 47.230 11.305 ;
        RECT 48.240 9.265 48.410 11.305 ;
        RECT 49.420 9.265 49.590 11.305 ;
        RECT 50.600 9.265 50.770 11.305 ;
        RECT 51.780 9.265 51.950 11.305 ;
        RECT 52.960 9.265 53.130 11.305 ;
        RECT 54.140 9.265 54.310 11.305 ;
        RECT 47.420 8.335 47.780 8.705 ;
        RECT 45.230 8.165 47.780 8.335 ;
        RECT 27.315 6.650 27.485 7.110 ;
        RECT 28.295 6.650 28.465 7.110 ;
        RECT 29.275 6.650 29.445 7.110 ;
        RECT 3.125 4.890 3.295 6.065 ;
        RECT 5.585 6.035 5.945 6.440 ;
        RECT 6.470 6.040 6.830 6.445 ;
        RECT 27.285 6.185 27.515 6.650 ;
        RECT 28.265 6.185 28.495 6.650 ;
        RECT 29.245 6.345 29.475 6.650 ;
        RECT 30.545 6.400 30.715 7.440 ;
        RECT 31.525 6.400 31.695 7.440 ;
        RECT 32.505 6.400 32.675 7.440 ;
        RECT 33.485 6.400 33.655 7.440 ;
        RECT 35.145 6.670 36.390 7.840 ;
        RECT 36.685 7.810 37.350 7.865 ;
        RECT 39.735 7.585 40.115 7.865 ;
        RECT 42.615 7.860 43.125 8.150 ;
        RECT 47.420 7.925 47.780 8.165 ;
        RECT 55.320 8.265 55.490 11.305 ;
        RECT 103.680 10.515 103.910 11.780 ;
        RECT 104.660 11.455 104.890 11.780 ;
        RECT 105.640 11.455 105.870 11.780 ;
        RECT 103.710 10.495 103.880 10.515 ;
        RECT 104.690 10.495 104.860 11.455 ;
        RECT 105.670 10.495 105.840 11.455 ;
        RECT 106.050 10.320 106.220 11.820 ;
        RECT 106.940 10.495 107.110 11.535 ;
        RECT 107.920 10.495 108.090 11.535 ;
        RECT 108.900 10.495 109.070 11.535 ;
        RECT 109.880 10.495 110.050 11.535 ;
        RECT 111.880 11.485 112.660 13.555 ;
        RECT 196.390 13.410 196.620 14.675 ;
        RECT 197.400 13.735 197.570 14.695 ;
        RECT 198.380 13.735 198.550 14.695 ;
        RECT 200.830 14.675 201.000 14.695 ;
        RECT 199.725 13.765 200.010 14.585 ;
        RECT 197.370 13.410 197.600 13.735 ;
        RECT 198.350 13.410 198.580 13.735 ;
        RECT 196.390 13.370 198.580 13.410 ;
        RECT 200.800 13.410 201.030 14.675 ;
        RECT 201.810 13.735 201.980 14.695 ;
        RECT 202.790 13.735 202.960 14.695 ;
        RECT 203.880 14.565 204.060 14.790 ;
        RECT 201.780 13.410 202.010 13.735 ;
        RECT 202.760 13.410 202.990 13.735 ;
        RECT 200.800 13.370 202.990 13.410 ;
        RECT 203.265 13.490 203.635 14.330 ;
        RECT 203.885 14.195 204.055 14.565 ;
        RECT 203.265 13.370 203.630 13.490 ;
        RECT 195.370 12.965 196.210 13.335 ;
        RECT 196.390 13.260 198.730 13.370 ;
        RECT 199.780 13.280 200.620 13.335 ;
        RECT 199.020 13.260 199.320 13.280 ;
        RECT 199.605 13.260 200.620 13.280 ;
        RECT 196.390 13.180 200.620 13.260 ;
        RECT 125.305 11.485 126.665 11.860 ;
        RECT 111.880 10.705 126.665 11.485 ;
        RECT 125.305 10.425 126.665 10.705 ;
        RECT 129.775 11.365 130.555 11.665 ;
        RECT 129.775 10.725 137.940 11.365 ;
        RECT 138.955 11.045 139.760 11.200 ;
        RECT 138.955 10.895 140.030 11.045 ;
        RECT 140.315 10.895 141.095 11.010 ;
        RECT 138.955 10.805 141.095 10.895 ;
        RECT 129.775 10.580 130.555 10.725 ;
        RECT 139.565 10.700 141.095 10.805 ;
        RECT 140.315 10.625 141.095 10.700 ;
        RECT 145.505 10.545 146.345 10.975 ;
        RECT 106.050 10.150 107.520 10.320 ;
        RECT 106.680 9.950 107.520 10.150 ;
        RECT 140.545 9.095 140.715 10.305 ;
        RECT 142.125 9.265 142.295 10.305 ;
        RECT 143.705 9.095 143.875 10.305 ;
        RECT 144.355 9.290 144.525 10.330 ;
        RECT 145.935 9.095 146.105 10.330 ;
        RECT 152.440 10.080 152.610 12.500 ;
        RECT 154.020 10.080 154.190 12.500 ;
        RECT 163.235 10.860 164.060 11.165 ;
        RECT 164.590 10.860 165.370 10.975 ;
        RECT 163.235 10.765 165.370 10.860 ;
        RECT 163.710 10.665 165.370 10.765 ;
        RECT 164.590 10.590 165.370 10.665 ;
        RECT 169.780 10.510 170.620 10.940 ;
        RECT 148.210 9.610 152.185 10.020 ;
        RECT 152.440 9.910 154.190 10.080 ;
        RECT 148.210 9.095 148.620 9.610 ;
        RECT 140.000 8.890 149.015 9.095 ;
        RECT 56.860 8.265 57.220 8.535 ;
        RECT 55.320 8.095 57.220 8.265 ;
        RECT 56.860 7.755 57.220 8.095 ;
        RECT 29.245 6.185 29.825 6.345 ;
        RECT 4.805 5.195 4.975 5.835 ;
        RECT 3.885 5.015 4.300 5.040 ;
        RECT -9.950 3.790 -9.780 4.830 ;
        RECT -8.970 3.790 -8.800 4.830 ;
        RECT -7.990 3.790 -7.820 4.830 ;
        RECT -7.010 3.790 -6.840 4.830 ;
        RECT 1.310 4.695 3.295 4.890 ;
        RECT 1.310 4.625 2.540 4.695 ;
        RECT -10.840 3.445 -9.370 3.615 ;
        RECT -66.605 3.390 -20.510 3.400 ;
        RECT -66.710 2.975 -20.510 3.390 ;
        RECT -10.210 3.245 -9.370 3.445 ;
        RECT -66.710 2.790 -30.775 2.975 ;
        RECT 2.345 2.170 2.540 4.625 ;
        RECT 3.125 3.865 3.295 4.695 ;
        RECT 3.465 4.890 4.300 5.015 ;
        RECT 5.685 4.890 5.855 5.835 ;
        RECT 6.565 4.890 6.735 5.835 ;
        RECT 7.570 5.025 7.740 6.135 ;
        RECT 8.010 5.195 8.180 6.135 ;
        RECT 9.770 6.000 10.495 6.185 ;
        RECT 9.770 5.385 9.940 6.000 ;
        RECT 10.325 5.385 10.495 6.000 ;
        RECT 9.770 5.200 10.495 5.385 ;
        RECT 9.770 5.195 9.940 5.200 ;
        RECT 7.155 4.890 7.955 5.025 ;
        RECT 3.465 4.650 7.955 4.890 ;
        RECT 8.175 4.695 8.585 5.025 ;
        RECT 9.290 4.865 10.095 5.025 ;
        RECT 8.795 4.690 10.095 4.865 ;
        RECT 3.465 4.560 3.865 4.650 ;
        RECT 4.355 3.740 4.525 4.380 ;
        RECT 4.945 3.740 5.115 4.380 ;
        RECT 5.535 3.740 5.705 4.380 ;
        RECT 6.565 3.740 6.735 4.380 ;
        RECT 7.005 3.740 7.175 4.650 ;
        RECT 8.015 3.715 8.185 4.355 ;
        RECT 8.455 3.715 8.625 4.355 ;
        RECT 4.475 3.200 4.875 3.570 ;
        RECT 5.130 3.205 5.520 3.570 ;
        RECT 6.830 3.200 7.220 3.570 ;
        RECT 8.000 3.445 8.395 3.540 ;
        RECT 8.795 3.445 8.970 4.690 ;
        RECT 9.290 4.525 10.095 4.690 ;
        RECT 10.325 4.855 10.495 5.200 ;
        RECT 11.935 5.015 12.350 5.040 ;
        RECT 11.935 4.855 12.770 5.015 ;
        RECT 10.325 4.685 12.770 4.855 ;
        RECT 9.145 3.680 9.315 4.320 ;
        RECT 10.325 3.680 10.495 4.685 ;
        RECT 11.505 3.680 11.675 4.685 ;
        RECT 11.935 4.650 12.770 4.685 ;
        RECT 12.370 4.560 12.770 4.650 ;
        RECT 12.940 4.890 13.110 6.065 ;
        RECT 13.480 5.015 13.895 5.040 ;
        RECT 13.480 4.890 14.315 5.015 ;
        RECT 12.940 4.650 14.315 4.890 ;
        RECT 12.940 3.865 13.110 4.650 ;
        RECT 13.915 4.560 14.315 4.650 ;
        RECT 14.485 4.890 14.655 6.065 ;
        RECT 27.285 5.995 29.825 6.185 ;
        RECT 27.285 5.955 29.475 5.995 ;
        RECT 17.815 4.890 18.625 5.195 ;
        RECT 14.485 4.695 18.625 4.890 ;
        RECT 14.485 3.865 14.655 4.695 ;
        RECT 17.815 4.425 18.625 4.695 ;
        RECT 27.285 4.690 27.515 5.955 ;
        RECT 28.265 5.630 28.495 5.955 ;
        RECT 29.245 5.630 29.475 5.955 ;
        RECT 27.315 4.670 27.485 4.690 ;
        RECT 28.295 4.670 28.465 5.630 ;
        RECT 29.275 4.670 29.445 5.630 ;
        RECT 29.655 4.495 29.825 5.995 ;
        RECT 30.545 4.670 30.715 5.710 ;
        RECT 31.525 4.670 31.695 5.710 ;
        RECT 32.505 4.670 32.675 5.710 ;
        RECT 33.485 4.670 33.655 5.710 ;
        RECT 40.140 5.225 40.310 7.265 ;
        RECT 41.320 5.225 41.490 7.265 ;
        RECT 42.500 5.225 42.670 7.265 ;
        RECT 43.680 5.225 43.850 7.265 ;
        RECT 44.860 5.225 45.030 7.265 ;
        RECT 46.040 5.225 46.210 7.265 ;
        RECT 47.220 5.225 47.390 7.265 ;
        RECT 140.000 6.450 140.205 8.890 ;
        RECT 140.545 7.320 140.715 8.360 ;
        RECT 142.125 7.320 142.295 8.890 ;
        RECT 143.705 7.320 143.875 8.360 ;
        RECT 144.355 7.320 144.525 8.890 ;
        RECT 145.375 8.610 149.015 8.890 ;
        RECT 145.935 7.320 146.105 8.360 ;
        RECT 149.030 7.110 149.235 7.225 ;
        RECT 152.440 7.180 152.610 9.910 ;
        RECT 154.020 9.640 154.190 9.910 ;
        RECT 154.020 9.470 159.955 9.640 ;
        RECT 154.020 7.180 154.190 9.470 ;
        RECT 155.600 7.180 155.770 9.470 ;
        RECT 157.180 7.180 157.350 9.470 ;
        RECT 146.300 6.780 149.235 7.110 ;
        RECT 140.000 6.420 145.350 6.450 ;
        RECT 137.535 6.230 145.350 6.420 ;
        RECT 131.390 4.940 132.350 5.470 ;
        RECT 135.660 4.940 137.250 5.030 ;
        RECT 131.390 4.615 137.250 4.940 ;
        RECT 29.655 4.325 31.125 4.495 ;
        RECT 30.285 4.125 31.125 4.325 ;
        RECT 131.390 4.180 132.350 4.615 ;
        RECT 135.660 4.530 137.250 4.615 ;
        RECT 137.535 3.860 137.725 6.230 ;
        RECT 140.000 6.075 145.350 6.230 ;
        RECT 140.000 5.995 140.650 6.075 ;
        RECT 138.275 4.425 138.635 5.175 ;
        RECT 140.480 4.675 140.650 5.995 ;
        RECT 141.270 4.675 141.440 5.715 ;
        RECT 142.060 4.675 142.230 5.715 ;
        RECT 142.850 4.675 143.020 5.715 ;
        RECT 143.640 4.675 143.810 6.075 ;
        RECT 144.230 4.675 144.400 5.715 ;
        RECT 145.020 4.675 145.190 5.715 ;
        RECT 159.650 4.995 159.955 9.470 ;
        RECT 164.820 9.060 164.990 10.270 ;
        RECT 166.400 9.230 166.570 10.270 ;
        RECT 167.980 9.060 168.150 10.270 ;
        RECT 168.630 9.255 168.800 10.295 ;
        RECT 170.210 9.060 170.380 10.295 ;
        RECT 176.115 10.190 176.285 12.610 ;
        RECT 177.695 10.190 177.865 12.610 ;
        RECT 172.670 9.720 175.860 10.130 ;
        RECT 176.115 10.020 177.865 10.190 ;
        RECT 172.670 9.060 173.080 9.720 ;
        RECT 164.275 8.855 173.290 9.060 ;
        RECT 164.275 6.415 164.480 8.855 ;
        RECT 164.820 7.285 164.990 8.325 ;
        RECT 166.400 7.285 166.570 8.855 ;
        RECT 167.980 7.285 168.150 8.325 ;
        RECT 168.630 7.285 168.800 8.855 ;
        RECT 169.650 8.575 173.290 8.855 ;
        RECT 170.210 7.285 170.380 8.325 ;
        RECT 176.115 7.290 176.285 10.020 ;
        RECT 177.695 9.750 177.865 10.020 ;
        RECT 184.720 9.975 184.890 12.395 ;
        RECT 186.300 9.975 186.470 12.395 ;
        RECT 195.470 10.995 195.665 12.965 ;
        RECT 196.390 12.715 196.620 13.180 ;
        RECT 197.370 12.715 197.600 13.180 ;
        RECT 198.350 13.050 200.620 13.180 ;
        RECT 198.350 13.020 198.730 13.050 ;
        RECT 198.350 12.715 198.580 13.020 ;
        RECT 196.420 12.255 196.590 12.715 ;
        RECT 197.400 12.255 197.570 12.715 ;
        RECT 198.380 12.255 198.550 12.715 ;
        RECT 199.020 12.620 199.320 13.050 ;
        RECT 199.605 12.990 200.620 13.050 ;
        RECT 199.780 12.965 200.620 12.990 ;
        RECT 200.800 13.180 203.630 13.370 ;
        RECT 200.800 12.715 201.030 13.180 ;
        RECT 201.780 12.715 202.010 13.180 ;
        RECT 202.760 13.020 203.630 13.180 ;
        RECT 203.855 13.460 204.090 14.195 ;
        RECT 204.375 14.160 204.545 14.620 ;
        RECT 204.860 14.515 205.070 14.790 ;
        RECT 204.370 13.900 204.550 14.160 ;
        RECT 204.865 14.080 205.035 14.515 ;
        RECT 205.355 14.170 205.525 14.620 ;
        RECT 205.830 14.510 206.040 14.790 ;
        RECT 205.355 14.080 205.540 14.170 ;
        RECT 205.845 14.080 206.015 14.510 ;
        RECT 206.335 14.170 206.505 14.620 ;
        RECT 206.810 14.535 207.020 14.790 ;
        RECT 217.380 14.790 220.520 14.960 ;
        RECT 209.545 14.675 209.715 14.695 ;
        RECT 205.360 13.900 205.540 14.080 ;
        RECT 206.330 13.900 206.510 14.170 ;
        RECT 206.825 14.080 206.995 14.535 ;
        RECT 207.315 14.120 207.485 14.620 ;
        RECT 207.300 13.900 207.510 14.120 ;
        RECT 204.370 13.730 207.510 13.900 ;
        RECT 203.855 13.090 204.715 13.460 ;
        RECT 206.635 13.290 207.510 13.730 ;
        RECT 209.515 13.410 209.745 14.675 ;
        RECT 210.525 13.735 210.695 14.695 ;
        RECT 211.505 13.735 211.675 14.695 ;
        RECT 214.330 14.675 214.500 14.695 ;
        RECT 213.225 14.195 213.510 14.585 ;
        RECT 212.205 13.970 213.510 14.195 ;
        RECT 210.495 13.410 210.725 13.735 ;
        RECT 211.475 13.410 211.705 13.735 ;
        RECT 209.515 13.370 211.705 13.410 ;
        RECT 208.495 13.290 209.335 13.335 ;
        RECT 202.760 12.715 202.990 13.020 ;
        RECT 200.830 12.255 201.000 12.715 ;
        RECT 201.810 12.255 201.980 12.715 ;
        RECT 202.790 12.255 202.960 12.715 ;
        RECT 203.855 12.415 204.090 13.090 ;
        RECT 206.635 13.005 209.335 13.290 ;
        RECT 206.635 12.895 207.510 13.005 ;
        RECT 208.495 12.965 209.335 13.005 ;
        RECT 209.515 13.300 211.855 13.370 ;
        RECT 212.205 13.300 212.430 13.970 ;
        RECT 213.225 13.765 213.510 13.970 ;
        RECT 214.300 13.410 214.530 14.675 ;
        RECT 215.310 13.735 215.480 14.695 ;
        RECT 216.290 13.735 216.460 14.695 ;
        RECT 217.380 14.565 217.560 14.790 ;
        RECT 215.280 13.410 215.510 13.735 ;
        RECT 216.260 13.410 216.490 13.735 ;
        RECT 214.300 13.370 216.490 13.410 ;
        RECT 216.765 13.490 217.135 14.330 ;
        RECT 217.385 14.195 217.555 14.565 ;
        RECT 216.765 13.370 217.130 13.490 ;
        RECT 209.515 13.180 212.430 13.300 ;
        RECT 204.355 12.725 207.510 12.895 ;
        RECT 204.355 12.520 204.560 12.725 ;
        RECT 203.885 12.065 204.055 12.415 ;
        RECT 203.860 11.775 204.080 12.065 ;
        RECT 204.375 12.005 204.545 12.520 ;
        RECT 204.865 12.120 205.035 12.545 ;
        RECT 205.345 12.480 205.550 12.725 ;
        RECT 204.840 11.775 205.060 12.120 ;
        RECT 205.355 12.005 205.525 12.480 ;
        RECT 205.845 12.120 206.015 12.545 ;
        RECT 206.315 12.480 206.520 12.725 ;
        RECT 207.300 12.690 207.510 12.725 ;
        RECT 209.515 12.715 209.745 13.180 ;
        RECT 210.495 12.715 210.725 13.180 ;
        RECT 211.475 13.075 212.430 13.180 ;
        RECT 212.680 13.280 212.980 13.285 ;
        RECT 213.280 13.280 214.120 13.335 ;
        RECT 211.475 13.020 211.855 13.075 ;
        RECT 211.475 12.715 211.705 13.020 ;
        RECT 205.820 11.775 206.040 12.120 ;
        RECT 206.335 12.005 206.505 12.480 ;
        RECT 206.825 12.065 206.995 12.545 ;
        RECT 207.300 12.525 207.505 12.690 ;
        RECT 207.270 12.475 207.505 12.525 ;
        RECT 206.805 11.775 207.025 12.065 ;
        RECT 207.270 11.865 207.500 12.475 ;
        RECT 209.545 12.255 209.715 12.715 ;
        RECT 210.525 12.255 210.695 12.715 ;
        RECT 211.505 12.255 211.675 12.715 ;
        RECT 212.105 12.500 212.405 13.075 ;
        RECT 212.680 12.990 214.120 13.280 ;
        RECT 212.680 12.625 212.980 12.990 ;
        RECT 213.280 12.965 214.120 12.990 ;
        RECT 214.300 13.180 217.130 13.370 ;
        RECT 214.300 12.715 214.530 13.180 ;
        RECT 215.280 12.715 215.510 13.180 ;
        RECT 216.260 13.020 217.130 13.180 ;
        RECT 217.355 13.460 217.590 14.195 ;
        RECT 217.875 14.160 218.045 14.620 ;
        RECT 218.360 14.515 218.570 14.790 ;
        RECT 217.870 13.900 218.050 14.160 ;
        RECT 218.365 14.080 218.535 14.515 ;
        RECT 218.855 14.170 219.025 14.620 ;
        RECT 219.330 14.510 219.540 14.790 ;
        RECT 218.855 14.080 219.040 14.170 ;
        RECT 219.345 14.080 219.515 14.510 ;
        RECT 219.835 14.170 220.005 14.620 ;
        RECT 220.310 14.535 220.520 14.790 ;
        RECT 223.045 14.675 223.215 14.695 ;
        RECT 218.860 13.900 219.040 14.080 ;
        RECT 219.830 13.900 220.010 14.170 ;
        RECT 220.325 14.080 220.495 14.535 ;
        RECT 220.815 14.120 220.985 14.620 ;
        RECT 220.800 13.900 221.010 14.120 ;
        RECT 217.870 13.730 221.010 13.900 ;
        RECT 217.355 13.090 218.215 13.460 ;
        RECT 220.135 13.305 221.010 13.730 ;
        RECT 223.015 13.410 223.245 14.675 ;
        RECT 224.025 13.735 224.195 14.695 ;
        RECT 225.005 13.735 225.175 14.695 ;
        RECT 223.995 13.410 224.225 13.735 ;
        RECT 224.975 13.410 225.205 13.735 ;
        RECT 223.015 13.370 225.205 13.410 ;
        RECT 221.995 13.305 222.835 13.335 ;
        RECT 216.260 12.715 216.490 13.020 ;
        RECT 214.330 12.255 214.500 12.715 ;
        RECT 215.310 12.255 215.480 12.715 ;
        RECT 216.290 12.255 216.460 12.715 ;
        RECT 217.355 12.415 217.590 13.090 ;
        RECT 220.135 13.040 222.835 13.305 ;
        RECT 220.135 12.895 221.010 13.040 ;
        RECT 221.995 12.965 222.835 13.040 ;
        RECT 223.015 13.325 225.355 13.370 ;
        RECT 223.015 13.315 225.765 13.325 ;
        RECT 223.015 13.180 225.770 13.315 ;
        RECT 217.855 12.725 221.010 12.895 ;
        RECT 217.855 12.520 218.060 12.725 ;
        RECT 217.385 12.065 217.555 12.415 ;
        RECT 203.860 11.605 207.025 11.775 ;
        RECT 217.360 11.775 217.580 12.065 ;
        RECT 217.875 12.005 218.045 12.520 ;
        RECT 218.365 12.120 218.535 12.545 ;
        RECT 218.845 12.480 219.050 12.725 ;
        RECT 218.340 11.775 218.560 12.120 ;
        RECT 218.855 12.005 219.025 12.480 ;
        RECT 219.345 12.120 219.515 12.545 ;
        RECT 219.815 12.480 220.020 12.725 ;
        RECT 220.800 12.690 221.010 12.725 ;
        RECT 223.015 12.715 223.245 13.180 ;
        RECT 223.995 12.715 224.225 13.180 ;
        RECT 224.975 13.130 225.770 13.180 ;
        RECT 255.070 13.150 255.240 15.190 ;
        RECT 224.975 13.020 225.355 13.130 ;
        RECT 224.975 12.715 225.205 13.020 ;
        RECT 219.320 11.775 219.540 12.120 ;
        RECT 219.835 12.005 220.005 12.480 ;
        RECT 220.325 12.065 220.495 12.545 ;
        RECT 220.800 12.475 221.005 12.690 ;
        RECT 220.305 11.775 220.525 12.065 ;
        RECT 220.815 12.005 220.985 12.475 ;
        RECT 223.045 12.255 223.215 12.715 ;
        RECT 224.025 12.255 224.195 12.715 ;
        RECT 225.005 12.255 225.175 12.715 ;
        RECT 217.360 11.605 220.525 11.775 ;
        RECT 198.815 11.425 199.475 11.480 ;
        RECT 221.430 11.425 222.090 11.490 ;
        RECT 198.815 11.230 224.120 11.425 ;
        RECT 225.530 11.340 225.770 13.130 ;
        RECT 256.250 12.820 256.420 15.190 ;
        RECT 258.080 13.150 258.250 15.190 ;
        RECT 259.260 13.150 259.430 15.190 ;
        RECT 260.440 13.150 260.610 15.190 ;
        RECT 256.250 12.650 257.290 12.820 ;
        RECT 252.550 12.055 253.745 12.335 ;
        RECT 256.125 12.055 256.505 12.355 ;
        RECT 252.550 11.750 256.505 12.055 ;
        RECT 257.120 12.205 257.290 12.650 ;
        RECT 259.005 12.205 259.515 12.445 ;
        RECT 257.120 12.035 259.515 12.205 ;
        RECT 261.620 12.220 261.790 15.190 ;
        RECT 263.450 13.150 263.620 15.190 ;
        RECT 264.630 13.150 264.800 15.190 ;
        RECT 265.810 13.150 265.980 15.190 ;
        RECT 266.990 13.150 267.160 15.190 ;
        RECT 268.170 13.150 268.340 15.190 ;
        RECT 269.350 13.150 269.520 15.190 ;
        RECT 270.530 13.150 270.700 15.190 ;
        RECT 263.810 12.220 264.170 12.590 ;
        RECT 261.620 12.050 264.170 12.220 ;
        RECT 198.815 11.180 199.475 11.230 ;
        RECT 221.430 11.190 222.090 11.230 ;
        RECT 207.835 10.995 208.495 11.050 ;
        RECT 212.540 10.995 213.225 11.045 ;
        RECT 195.470 10.800 224.120 10.995 ;
        RECT 182.980 9.750 184.465 9.915 ;
        RECT 177.695 9.580 184.465 9.750 ;
        RECT 177.695 7.290 177.865 9.580 ;
        RECT 179.275 7.290 179.445 9.580 ;
        RECT 180.855 7.290 181.025 9.580 ;
        RECT 182.980 9.505 184.465 9.580 ;
        RECT 184.720 9.805 186.470 9.975 ;
        RECT 173.305 7.075 173.510 7.190 ;
        RECT 184.720 7.075 184.890 9.805 ;
        RECT 186.300 9.535 186.470 9.805 ;
        RECT 192.145 9.710 193.105 10.065 ;
        RECT 195.765 9.710 196.225 10.800 ;
        RECT 207.835 10.750 208.495 10.800 ;
        RECT 212.540 10.745 213.225 10.800 ;
        RECT 225.475 10.655 225.775 11.340 ;
        RECT 252.550 11.075 253.745 11.750 ;
        RECT 256.125 11.470 256.505 11.750 ;
        RECT 259.005 11.745 259.515 12.035 ;
        RECT 263.810 11.810 264.170 12.050 ;
        RECT 271.710 12.150 271.880 15.190 ;
        RECT 273.250 12.150 273.610 12.420 ;
        RECT 271.710 11.980 273.610 12.150 ;
        RECT 273.250 11.640 273.610 11.980 ;
        RECT 200.805 9.985 203.970 10.155 ;
        RECT 192.145 9.535 196.225 9.710 ;
        RECT 186.300 9.365 196.225 9.535 ;
        RECT 186.300 7.075 186.470 9.365 ;
        RECT 187.880 7.075 188.050 9.365 ;
        RECT 189.460 7.075 189.630 9.365 ;
        RECT 192.145 9.250 196.225 9.365 ;
        RECT 200.345 9.285 200.515 9.755 ;
        RECT 200.805 9.695 201.025 9.985 ;
        RECT 192.145 8.775 193.105 9.250 ;
        RECT 200.325 9.070 200.530 9.285 ;
        RECT 200.835 9.215 201.005 9.695 ;
        RECT 201.325 9.280 201.495 9.755 ;
        RECT 201.790 9.640 202.010 9.985 ;
        RECT 200.320 9.035 200.530 9.070 ;
        RECT 201.310 9.035 201.515 9.280 ;
        RECT 201.815 9.215 201.985 9.640 ;
        RECT 202.305 9.280 202.475 9.755 ;
        RECT 202.770 9.640 202.990 9.985 ;
        RECT 202.280 9.035 202.485 9.280 ;
        RECT 202.795 9.215 202.965 9.640 ;
        RECT 203.285 9.240 203.455 9.755 ;
        RECT 203.750 9.695 203.970 9.985 ;
        RECT 214.305 9.985 217.470 10.155 ;
        RECT 203.775 9.345 203.945 9.695 ;
        RECT 203.270 9.035 203.475 9.240 ;
        RECT 200.320 8.875 203.475 9.035 ;
        RECT 199.945 8.865 203.475 8.875 ;
        RECT 199.945 8.575 201.195 8.865 ;
        RECT 203.740 8.670 203.975 9.345 ;
        RECT 204.870 9.045 205.040 9.505 ;
        RECT 205.850 9.045 206.020 9.505 ;
        RECT 206.830 9.045 207.000 9.505 ;
        RECT 204.840 8.740 205.070 9.045 ;
        RECT 200.320 8.030 201.195 8.575 ;
        RECT 203.115 8.300 203.975 8.670 ;
        RECT 200.320 7.860 203.460 8.030 ;
        RECT 200.320 7.640 200.530 7.860 ;
        RECT 200.345 7.140 200.515 7.640 ;
        RECT 200.835 7.225 201.005 7.680 ;
        RECT 201.320 7.590 201.500 7.860 ;
        RECT 202.290 7.680 202.470 7.860 ;
        RECT 170.575 6.745 173.510 7.075 ;
        RECT 200.810 6.970 201.020 7.225 ;
        RECT 201.325 7.140 201.495 7.590 ;
        RECT 201.815 7.250 201.985 7.680 ;
        RECT 202.290 7.590 202.475 7.680 ;
        RECT 201.790 6.970 202.000 7.250 ;
        RECT 202.305 7.140 202.475 7.590 ;
        RECT 202.795 7.245 202.965 7.680 ;
        RECT 203.280 7.600 203.460 7.860 ;
        RECT 202.760 6.970 202.970 7.245 ;
        RECT 203.285 7.140 203.455 7.600 ;
        RECT 203.740 7.565 203.975 8.300 ;
        RECT 204.200 8.580 205.070 8.740 ;
        RECT 205.820 8.580 206.050 9.045 ;
        RECT 206.800 8.580 207.030 9.045 ;
        RECT 208.050 8.795 208.350 9.590 ;
        RECT 209.055 9.045 209.225 9.505 ;
        RECT 210.035 9.045 210.205 9.505 ;
        RECT 211.015 9.045 211.185 9.505 ;
        RECT 213.845 9.285 214.015 9.755 ;
        RECT 214.305 9.695 214.525 9.985 ;
        RECT 213.825 9.070 214.030 9.285 ;
        RECT 214.335 9.215 214.505 9.695 ;
        RECT 214.825 9.280 214.995 9.755 ;
        RECT 215.290 9.640 215.510 9.985 ;
        RECT 204.200 8.390 207.030 8.580 ;
        RECT 207.210 8.480 208.350 8.795 ;
        RECT 209.025 8.740 209.255 9.045 ;
        RECT 208.535 8.580 209.255 8.740 ;
        RECT 210.005 8.580 210.235 9.045 ;
        RECT 210.985 8.580 211.215 9.045 ;
        RECT 213.820 9.035 214.030 9.070 ;
        RECT 214.810 9.035 215.015 9.280 ;
        RECT 215.315 9.215 215.485 9.640 ;
        RECT 215.805 9.280 215.975 9.755 ;
        RECT 216.270 9.640 216.490 9.985 ;
        RECT 215.780 9.035 215.985 9.280 ;
        RECT 216.295 9.215 216.465 9.640 ;
        RECT 216.785 9.240 216.955 9.755 ;
        RECT 217.250 9.695 217.470 9.985 ;
        RECT 217.275 9.345 217.445 9.695 ;
        RECT 216.770 9.035 216.975 9.240 ;
        RECT 213.820 8.865 216.975 9.035 ;
        RECT 207.210 8.425 208.050 8.480 ;
        RECT 204.200 8.270 204.565 8.390 ;
        RECT 203.775 7.195 203.945 7.565 ;
        RECT 204.195 7.430 204.565 8.270 ;
        RECT 204.840 8.350 207.030 8.390 ;
        RECT 204.840 8.025 205.070 8.350 ;
        RECT 205.820 8.025 206.050 8.350 ;
        RECT 203.770 6.970 203.950 7.195 ;
        RECT 204.870 7.065 205.040 8.025 ;
        RECT 205.850 7.065 206.020 8.025 ;
        RECT 206.800 7.085 207.030 8.350 ;
        RECT 208.535 8.390 211.215 8.580 ;
        RECT 211.395 8.760 212.235 8.795 ;
        RECT 211.395 8.460 212.345 8.760 ;
        RECT 213.365 8.565 214.695 8.865 ;
        RECT 217.240 8.670 217.475 9.345 ;
        RECT 218.370 9.045 218.540 9.505 ;
        RECT 219.350 9.045 219.520 9.505 ;
        RECT 220.330 9.045 220.500 9.505 ;
        RECT 218.340 8.740 218.570 9.045 ;
        RECT 211.395 8.425 212.235 8.460 ;
        RECT 207.820 7.745 208.105 7.995 ;
        RECT 208.535 7.745 208.845 8.390 ;
        RECT 209.025 8.350 211.215 8.390 ;
        RECT 209.025 8.025 209.255 8.350 ;
        RECT 210.005 8.025 210.235 8.350 ;
        RECT 207.820 7.435 208.845 7.745 ;
        RECT 207.820 7.175 208.105 7.435 ;
        RECT 206.830 7.065 207.000 7.085 ;
        RECT 209.055 7.065 209.225 8.025 ;
        RECT 210.035 7.065 210.205 8.025 ;
        RECT 210.985 7.085 211.215 8.350 ;
        RECT 213.820 8.030 214.695 8.565 ;
        RECT 216.615 8.300 217.475 8.670 ;
        RECT 213.820 7.860 216.960 8.030 ;
        RECT 213.820 7.640 214.030 7.860 ;
        RECT 213.845 7.140 214.015 7.640 ;
        RECT 214.335 7.225 214.505 7.680 ;
        RECT 214.820 7.590 215.000 7.860 ;
        RECT 215.790 7.680 215.970 7.860 ;
        RECT 211.015 7.065 211.185 7.085 ;
        RECT 200.810 6.800 203.950 6.970 ;
        RECT 214.310 6.970 214.520 7.225 ;
        RECT 214.825 7.140 214.995 7.590 ;
        RECT 215.315 7.250 215.485 7.680 ;
        RECT 215.790 7.590 215.975 7.680 ;
        RECT 215.290 6.970 215.500 7.250 ;
        RECT 215.805 7.140 215.975 7.590 ;
        RECT 216.295 7.245 216.465 7.680 ;
        RECT 216.780 7.600 216.960 7.860 ;
        RECT 216.260 6.970 216.470 7.245 ;
        RECT 216.785 7.140 216.955 7.600 ;
        RECT 217.240 7.565 217.475 8.300 ;
        RECT 217.700 8.580 218.570 8.740 ;
        RECT 219.320 8.580 219.550 9.045 ;
        RECT 220.300 8.580 220.530 9.045 ;
        RECT 221.610 8.795 221.910 9.515 ;
        RECT 222.555 9.045 222.725 9.505 ;
        RECT 223.535 9.045 223.705 9.505 ;
        RECT 224.515 9.045 224.685 9.505 ;
        RECT 217.700 8.390 220.530 8.580 ;
        RECT 220.710 8.485 221.910 8.795 ;
        RECT 222.525 8.740 222.755 9.045 ;
        RECT 222.090 8.580 222.755 8.740 ;
        RECT 223.505 8.580 223.735 9.045 ;
        RECT 224.485 8.580 224.715 9.045 ;
        RECT 225.530 8.795 225.770 10.655 ;
        RECT 226.755 9.675 227.485 10.605 ;
        RECT 227.000 9.260 227.220 9.675 ;
        RECT 228.385 9.495 228.555 9.955 ;
        RECT 229.365 9.495 229.535 9.955 ;
        RECT 230.345 9.495 230.515 9.955 ;
        RECT 227.000 9.245 227.825 9.260 ;
        RECT 227.000 8.990 228.175 9.245 ;
        RECT 227.335 8.875 228.175 8.990 ;
        RECT 228.355 9.030 228.585 9.495 ;
        RECT 229.335 9.030 229.565 9.495 ;
        RECT 230.315 9.190 230.545 9.495 ;
        RECT 233.185 9.190 234.805 9.985 ;
        RECT 230.315 9.030 234.805 9.190 ;
        RECT 220.710 8.480 221.725 8.485 ;
        RECT 220.710 8.425 221.550 8.480 ;
        RECT 217.700 8.270 218.065 8.390 ;
        RECT 217.275 7.195 217.445 7.565 ;
        RECT 217.695 7.430 218.065 8.270 ;
        RECT 218.340 8.350 220.530 8.390 ;
        RECT 218.340 8.025 218.570 8.350 ;
        RECT 219.320 8.025 219.550 8.350 ;
        RECT 217.270 6.970 217.450 7.195 ;
        RECT 218.370 7.065 218.540 8.025 ;
        RECT 219.350 7.065 219.520 8.025 ;
        RECT 220.300 7.085 220.530 8.350 ;
        RECT 222.090 8.390 224.715 8.580 ;
        RECT 224.895 8.575 225.770 8.795 ;
        RECT 228.355 8.840 234.805 9.030 ;
        RECT 228.355 8.800 230.545 8.840 ;
        RECT 224.895 8.425 225.735 8.575 ;
        RECT 221.320 7.740 221.605 7.995 ;
        RECT 222.090 7.740 222.320 8.390 ;
        RECT 222.525 8.350 224.715 8.390 ;
        RECT 222.525 8.025 222.755 8.350 ;
        RECT 223.505 8.025 223.735 8.350 ;
        RECT 221.320 7.495 222.320 7.740 ;
        RECT 221.320 7.175 221.605 7.495 ;
        RECT 220.330 7.065 220.500 7.085 ;
        RECT 222.555 7.065 222.725 8.025 ;
        RECT 223.535 7.065 223.705 8.025 ;
        RECT 224.485 7.085 224.715 8.350 ;
        RECT 228.355 7.535 228.585 8.800 ;
        RECT 229.335 8.475 229.565 8.800 ;
        RECT 230.315 8.475 230.545 8.800 ;
        RECT 228.385 7.515 228.555 7.535 ;
        RECT 229.365 7.515 229.535 8.475 ;
        RECT 230.345 7.515 230.515 8.475 ;
        RECT 233.185 8.430 234.805 8.840 ;
        RECT 239.480 9.500 241.080 9.960 ;
        RECT 252.705 9.500 253.600 11.075 ;
        RECT 239.480 8.605 253.600 9.500 ;
        RECT 256.530 9.110 256.700 11.150 ;
        RECT 257.710 9.110 257.880 11.150 ;
        RECT 258.890 9.110 259.060 11.150 ;
        RECT 260.070 9.110 260.240 11.150 ;
        RECT 261.250 9.110 261.420 11.150 ;
        RECT 262.430 9.110 262.600 11.150 ;
        RECT 263.610 9.110 263.780 11.150 ;
        RECT 239.480 8.180 241.080 8.605 ;
        RECT 224.515 7.065 224.685 7.085 ;
        RECT 214.310 6.800 217.450 6.970 ;
        RECT 231.805 6.475 232.535 6.785 ;
        RECT 164.275 6.385 169.625 6.415 ;
        RECT 161.810 6.195 169.625 6.385 ;
        RECT 159.650 4.905 161.525 4.995 ;
        RECT 159.610 4.580 161.525 4.905 ;
        RECT 159.935 4.495 161.525 4.580 ;
        RECT 140.795 4.425 141.150 4.475 ;
        RECT 143.095 4.425 143.485 4.480 ;
        RECT 138.275 4.090 145.165 4.425 ;
        RECT 137.535 3.675 144.400 3.860 ;
        RECT 8.000 3.235 8.970 3.445 ;
        RECT 8.000 3.140 8.395 3.235 ;
        RECT 9.260 3.120 11.425 3.510 ;
        RECT 3.690 2.170 4.875 2.305 ;
        RECT 2.345 1.975 4.875 2.170 ;
        RECT 3.690 1.825 4.875 1.975 ;
        RECT 5.170 1.805 10.060 2.285 ;
        RECT 131.205 1.835 132.165 2.730 ;
        RECT 140.480 2.250 140.650 3.465 ;
        RECT 141.270 2.425 141.440 3.465 ;
        RECT 142.060 2.425 142.230 3.675 ;
        RECT 142.850 2.425 143.020 3.465 ;
        RECT 143.640 2.250 143.810 3.465 ;
        RECT 144.230 2.425 144.400 3.675 ;
        RECT 144.580 3.620 144.925 4.090 ;
        RECT 146.855 3.605 147.230 4.345 ;
        RECT 145.020 2.425 145.190 3.465 ;
        RECT 146.950 2.875 147.135 3.605 ;
        RECT 146.950 2.465 148.985 2.875 ;
        RECT 146.950 2.250 147.135 2.465 ;
        RECT 140.345 2.065 147.135 2.250 ;
        RECT 140.245 1.835 141.065 1.895 ;
        RECT 131.205 1.630 141.065 1.835 ;
        RECT 131.205 1.440 132.165 1.630 ;
        RECT 140.245 1.545 141.065 1.630 ;
        RECT 148.575 1.790 148.985 2.465 ;
        RECT 148.575 1.380 152.185 1.790 ;
        RECT 152.440 1.490 152.610 4.220 ;
        RECT 154.020 1.930 154.190 4.220 ;
        RECT 155.600 1.930 155.770 4.220 ;
        RECT 157.180 1.930 157.350 4.220 ;
        RECT 161.810 3.825 162.000 6.195 ;
        RECT 164.275 6.040 169.625 6.195 ;
        RECT 231.805 6.145 234.320 6.475 ;
        RECT 164.275 5.960 164.925 6.040 ;
        RECT 162.550 4.390 162.910 5.140 ;
        RECT 164.755 4.640 164.925 5.960 ;
        RECT 165.545 4.640 165.715 5.680 ;
        RECT 166.335 4.640 166.505 5.680 ;
        RECT 167.125 4.640 167.295 5.680 ;
        RECT 167.915 4.640 168.085 6.040 ;
        RECT 231.805 5.855 232.535 6.145 ;
        RECT 168.505 4.640 168.675 5.680 ;
        RECT 169.295 4.640 169.465 5.680 ;
        RECT 165.070 4.390 165.425 4.440 ;
        RECT 167.370 4.390 167.760 4.445 ;
        RECT 162.550 4.055 169.440 4.390 ;
        RECT 161.810 3.640 168.675 3.825 ;
        RECT 164.755 2.215 164.925 3.430 ;
        RECT 165.545 2.390 165.715 3.430 ;
        RECT 166.335 2.390 166.505 3.640 ;
        RECT 167.125 2.390 167.295 3.430 ;
        RECT 167.915 2.215 168.085 3.430 ;
        RECT 168.505 2.390 168.675 3.640 ;
        RECT 168.855 3.585 169.200 4.055 ;
        RECT 171.130 3.570 171.505 4.310 ;
        RECT 169.295 2.390 169.465 3.430 ;
        RECT 171.225 2.735 171.410 3.570 ;
        RECT 171.225 2.325 173.080 2.735 ;
        RECT 171.225 2.215 171.410 2.325 ;
        RECT 164.620 2.030 171.410 2.215 ;
        RECT 154.020 1.800 158.585 1.930 ;
        RECT 172.670 1.905 173.080 2.325 ;
        RECT 164.520 1.800 165.340 1.860 ;
        RECT 154.020 1.760 165.340 1.800 ;
        RECT 154.020 1.490 154.190 1.760 ;
        RECT 158.275 1.595 165.340 1.760 ;
        RECT 164.520 1.510 165.340 1.595 ;
        RECT 172.670 1.495 175.860 1.905 ;
        RECT 176.115 1.605 176.285 4.335 ;
        RECT 177.695 2.045 177.865 4.335 ;
        RECT 179.275 2.045 179.445 4.335 ;
        RECT 180.855 2.045 181.025 4.335 ;
        RECT 182.980 2.045 184.465 2.120 ;
        RECT 177.695 1.875 184.465 2.045 ;
        RECT 177.695 1.605 177.865 1.875 ;
        RECT 182.980 1.710 184.465 1.875 ;
        RECT 184.720 1.820 184.890 4.550 ;
        RECT 186.300 2.260 186.470 4.550 ;
        RECT 187.880 2.260 188.050 4.550 ;
        RECT 189.460 2.260 189.630 4.550 ;
        RECT 192.255 2.415 193.215 2.825 ;
        RECT 192.255 2.260 193.285 2.415 ;
        RECT 186.300 2.090 193.285 2.260 ;
        RECT 186.300 1.820 186.470 2.090 ;
        RECT 152.440 1.320 154.190 1.490 ;
        RECT 107.540 0.505 108.380 0.705 ;
        RECT 106.910 0.335 108.380 0.505 ;
        RECT 100.320 0.140 100.490 0.160 ;
        RECT -65.985 -1.370 -35.815 -0.675 ;
        RECT -17.550 -1.310 -16.710 -1.110 ;
        RECT -65.985 -1.890 -28.600 -1.370 ;
        RECT -18.180 -1.480 -16.710 -1.310 ;
        RECT 100.290 -1.125 100.520 0.140 ;
        RECT 101.300 -0.800 101.470 0.160 ;
        RECT 102.280 -0.800 102.450 0.160 ;
        RECT 104.570 0.140 104.740 0.160 ;
        RECT 101.270 -1.125 101.500 -0.800 ;
        RECT 102.250 -1.125 102.480 -0.800 ;
        RECT 100.290 -1.165 102.480 -1.125 ;
        RECT 104.540 -1.125 104.770 0.140 ;
        RECT 105.550 -0.800 105.720 0.160 ;
        RECT 106.530 -0.800 106.700 0.160 ;
        RECT 105.520 -1.125 105.750 -0.800 ;
        RECT 106.500 -1.125 106.730 -0.800 ;
        RECT 104.540 -1.165 106.730 -1.125 ;
        RECT 106.910 -1.165 107.080 0.335 ;
        RECT 100.290 -1.240 103.310 -1.165 ;
        RECT 103.520 -1.240 104.360 -1.200 ;
        RECT 100.290 -1.355 104.360 -1.240 ;
        RECT -24.770 -1.675 -24.600 -1.655 ;
        RECT -65.985 -2.265 -35.815 -1.890 ;
        RECT -24.800 -2.940 -24.570 -1.675 ;
        RECT -23.790 -2.615 -23.620 -1.655 ;
        RECT -22.810 -2.615 -22.640 -1.655 ;
        RECT -20.520 -1.675 -20.350 -1.655 ;
        RECT -23.820 -2.940 -23.590 -2.615 ;
        RECT -22.840 -2.940 -22.610 -2.615 ;
        RECT -24.800 -2.980 -22.610 -2.940 ;
        RECT -20.550 -2.940 -20.320 -1.675 ;
        RECT -19.540 -2.615 -19.370 -1.655 ;
        RECT -18.560 -2.615 -18.390 -1.655 ;
        RECT -19.570 -2.940 -19.340 -2.615 ;
        RECT -18.590 -2.940 -18.360 -2.615 ;
        RECT -20.550 -2.980 -18.360 -2.940 ;
        RECT -18.180 -2.980 -18.010 -1.480 ;
        RECT -24.800 -3.055 -21.780 -2.980 ;
        RECT -21.570 -3.055 -20.730 -3.015 ;
        RECT -24.800 -3.170 -20.730 -3.055 ;
        RECT -127.765 -4.030 -125.825 -3.270 ;
        RECT -29.880 -4.030 -29.000 -3.920 ;
        RECT -127.765 -4.715 -29.000 -4.030 ;
        RECT -25.260 -4.345 -25.090 -3.555 ;
        RECT -24.800 -3.635 -24.570 -3.170 ;
        RECT -24.770 -4.095 -24.600 -3.635 ;
        RECT -24.280 -4.345 -24.110 -3.555 ;
        RECT -23.820 -3.635 -23.590 -3.170 ;
        RECT -22.840 -3.315 -20.730 -3.170 ;
        RECT -22.840 -3.330 -21.780 -3.315 ;
        RECT -23.790 -4.095 -23.620 -3.635 ;
        RECT -23.300 -4.345 -23.130 -3.555 ;
        RECT -22.840 -3.635 -22.610 -3.330 ;
        RECT -21.570 -3.385 -20.730 -3.315 ;
        RECT -20.550 -3.170 -18.010 -2.980 ;
        RECT -22.810 -4.095 -22.640 -3.635 ;
        RECT -25.260 -4.350 -22.840 -4.345 ;
        RECT -21.010 -4.350 -20.840 -3.555 ;
        RECT -20.550 -3.635 -20.320 -3.170 ;
        RECT -20.520 -4.095 -20.350 -3.635 ;
        RECT -20.030 -4.350 -19.860 -3.555 ;
        RECT -19.570 -3.635 -19.340 -3.170 ;
        RECT -18.590 -3.330 -18.010 -3.170 ;
        RECT -17.780 -2.940 -17.610 -1.655 ;
        RECT -17.290 -2.695 -17.120 -1.655 ;
        RECT -16.800 -2.940 -16.630 -1.655 ;
        RECT -16.310 -2.695 -16.140 -1.655 ;
        RECT -15.820 -2.940 -15.650 -1.655 ;
        RECT -15.330 -2.695 -15.160 -1.655 ;
        RECT -14.840 -2.940 -14.670 -1.655 ;
        RECT -14.350 -2.695 -14.180 -1.655 ;
        RECT -13.860 -2.940 -13.690 -1.655 ;
        RECT 100.290 -1.820 100.520 -1.355 ;
        RECT 101.270 -1.820 101.500 -1.355 ;
        RECT 102.250 -1.500 104.360 -1.355 ;
        RECT 102.250 -1.515 103.310 -1.500 ;
        RECT 102.250 -1.820 102.480 -1.515 ;
        RECT 103.520 -1.570 104.360 -1.500 ;
        RECT 104.540 -1.355 107.080 -1.165 ;
        RECT 104.540 -1.820 104.770 -1.355 ;
        RECT 105.520 -1.820 105.750 -1.355 ;
        RECT 106.500 -1.515 107.080 -1.355 ;
        RECT 107.310 -1.125 107.480 0.160 ;
        RECT 107.800 -0.880 107.970 0.160 ;
        RECT 108.290 -1.125 108.460 0.160 ;
        RECT 108.780 -0.880 108.950 0.160 ;
        RECT 109.270 -1.125 109.440 0.160 ;
        RECT 109.760 -0.880 109.930 0.160 ;
        RECT 110.250 -1.125 110.420 0.160 ;
        RECT 110.740 -0.880 110.910 0.160 ;
        RECT 111.230 -1.125 111.400 0.160 ;
        RECT 139.045 -0.125 139.215 0.915 ;
        RECT 140.625 -0.125 140.795 0.915 ;
        RECT 142.205 -0.125 142.375 0.915 ;
        RECT 143.785 -0.125 143.955 0.915 ;
        RECT 145.365 -0.125 145.535 0.915 ;
        RECT 146.945 -0.125 147.115 0.915 ;
        RECT 152.440 -1.100 152.610 1.320 ;
        RECT 154.020 -1.100 154.190 1.320 ;
        RECT 176.115 1.435 177.865 1.605 ;
        RECT 163.320 -0.160 163.490 0.880 ;
        RECT 164.900 -0.160 165.070 0.880 ;
        RECT 166.480 -0.160 166.650 0.880 ;
        RECT 168.060 -0.160 168.230 0.880 ;
        RECT 169.640 -0.160 169.810 0.880 ;
        RECT 171.220 -0.160 171.390 0.880 ;
        RECT 176.115 -0.985 176.285 1.435 ;
        RECT 177.695 -0.985 177.865 1.435 ;
        RECT 184.720 1.650 186.470 1.820 ;
        RECT 184.720 -0.770 184.890 1.650 ;
        RECT 186.300 -0.770 186.470 1.650 ;
        RECT 192.255 1.900 193.285 2.090 ;
        RECT 192.255 1.535 193.215 1.900 ;
        RECT 107.310 -1.295 111.400 -1.125 ;
        RECT 106.500 -1.820 106.730 -1.515 ;
        RECT 30.360 -2.020 31.200 -1.820 ;
        RECT 29.730 -2.190 31.200 -2.020 ;
        RECT 23.140 -2.385 23.310 -2.365 ;
        RECT -17.780 -3.110 -13.690 -2.940 ;
        RECT -19.540 -4.095 -19.370 -3.635 ;
        RECT -19.050 -4.350 -18.880 -3.555 ;
        RECT -18.590 -3.635 -18.360 -3.330 ;
        RECT -18.560 -4.095 -18.390 -3.635 ;
        RECT -25.305 -4.690 -18.385 -4.350 ;
        RECT -17.780 -4.425 -17.610 -3.110 ;
        RECT -17.290 -4.425 -17.120 -3.385 ;
        RECT -16.800 -4.425 -16.630 -3.110 ;
        RECT -16.310 -4.425 -16.140 -3.385 ;
        RECT -15.820 -4.425 -15.650 -3.110 ;
        RECT -15.330 -4.425 -15.160 -3.385 ;
        RECT -14.840 -4.425 -14.670 -3.110 ;
        RECT -14.350 -4.425 -14.180 -3.385 ;
        RECT -13.860 -4.425 -13.690 -3.110 ;
        RECT 23.110 -3.650 23.340 -2.385 ;
        RECT 24.120 -3.325 24.290 -2.365 ;
        RECT 25.100 -3.325 25.270 -2.365 ;
        RECT 27.390 -2.385 27.560 -2.365 ;
        RECT 24.090 -3.650 24.320 -3.325 ;
        RECT 25.070 -3.650 25.300 -3.325 ;
        RECT 23.110 -3.690 25.300 -3.650 ;
        RECT 27.360 -3.650 27.590 -2.385 ;
        RECT 28.370 -3.325 28.540 -2.365 ;
        RECT 29.350 -3.325 29.520 -2.365 ;
        RECT 28.340 -3.650 28.570 -3.325 ;
        RECT 29.320 -3.650 29.550 -3.325 ;
        RECT 27.360 -3.690 29.550 -3.650 ;
        RECT 29.730 -3.690 29.900 -2.190 ;
        RECT 100.320 -2.280 100.490 -1.820 ;
        RECT 101.300 -2.280 101.470 -1.820 ;
        RECT 102.280 -2.280 102.450 -1.820 ;
        RECT 104.570 -2.280 104.740 -1.820 ;
        RECT 105.550 -2.280 105.720 -1.820 ;
        RECT 106.530 -2.280 106.700 -1.820 ;
        RECT 23.110 -3.765 26.130 -3.690 ;
        RECT 26.340 -3.765 27.180 -3.725 ;
        RECT 23.110 -3.880 27.180 -3.765 ;
        RECT 23.110 -4.345 23.340 -3.880 ;
        RECT 24.090 -4.345 24.320 -3.880 ;
        RECT 25.070 -4.025 27.180 -3.880 ;
        RECT 25.070 -4.040 26.130 -4.025 ;
        RECT 25.070 -4.345 25.300 -4.040 ;
        RECT 26.340 -4.095 27.180 -4.025 ;
        RECT 27.360 -3.880 29.900 -3.690 ;
        RECT 27.360 -4.345 27.590 -3.880 ;
        RECT 28.340 -4.345 28.570 -3.880 ;
        RECT 29.320 -4.040 29.900 -3.880 ;
        RECT 30.130 -3.650 30.300 -2.365 ;
        RECT 30.620 -3.405 30.790 -2.365 ;
        RECT 31.110 -3.650 31.280 -2.365 ;
        RECT 31.600 -3.405 31.770 -2.365 ;
        RECT 32.090 -3.650 32.260 -2.365 ;
        RECT 32.580 -3.405 32.750 -2.365 ;
        RECT 33.070 -3.650 33.240 -2.365 ;
        RECT 33.560 -3.405 33.730 -2.365 ;
        RECT 34.050 -3.650 34.220 -2.365 ;
        RECT 30.130 -3.820 34.220 -3.650 ;
        RECT 29.320 -4.345 29.550 -4.040 ;
        RECT -127.765 -5.250 -125.825 -4.715 ;
        RECT -29.880 -5.025 -29.000 -4.715 ;
        RECT -21.055 -5.375 -18.385 -4.690 ;
        RECT 23.140 -4.805 23.310 -4.345 ;
        RECT 24.120 -4.805 24.290 -4.345 ;
        RECT 25.100 -4.805 25.270 -4.345 ;
        RECT 27.390 -4.805 27.560 -4.345 ;
        RECT 28.370 -4.805 28.540 -4.345 ;
        RECT 29.350 -4.805 29.520 -4.345 ;
        RECT 30.130 -5.135 30.300 -3.820 ;
        RECT 30.620 -5.135 30.790 -4.095 ;
        RECT 31.110 -5.135 31.280 -3.820 ;
        RECT 31.600 -5.135 31.770 -4.095 ;
        RECT 32.090 -5.135 32.260 -3.820 ;
        RECT 32.580 -5.135 32.750 -4.095 ;
        RECT 33.070 -5.135 33.240 -3.820 ;
        RECT 33.560 -5.135 33.730 -4.095 ;
        RECT 34.050 -5.135 34.220 -3.820 ;
        RECT 38.475 -4.515 38.645 -2.475 ;
        RECT 39.655 -4.845 39.825 -2.475 ;
        RECT 41.485 -4.515 41.655 -2.475 ;
        RECT 42.665 -4.515 42.835 -2.475 ;
        RECT 43.845 -4.515 44.015 -2.475 ;
        RECT 39.655 -5.015 40.695 -4.845 ;
        RECT -21.010 -6.170 -20.840 -5.375 ;
        RECT -20.520 -6.090 -20.350 -5.630 ;
        RECT -20.550 -6.555 -20.320 -6.090 ;
        RECT -20.030 -6.170 -19.860 -5.375 ;
        RECT -19.540 -6.090 -19.370 -5.630 ;
        RECT -19.570 -6.555 -19.340 -6.090 ;
        RECT -19.050 -6.170 -18.880 -5.375 ;
        RECT -18.560 -6.090 -18.390 -5.630 ;
        RECT -18.590 -6.395 -18.360 -6.090 ;
        RECT -18.590 -6.555 -18.010 -6.395 ;
        RECT -20.550 -6.745 -18.010 -6.555 ;
        RECT -20.550 -6.785 -18.360 -6.745 ;
        RECT -20.550 -8.050 -20.320 -6.785 ;
        RECT -19.570 -7.110 -19.340 -6.785 ;
        RECT -18.590 -7.110 -18.360 -6.785 ;
        RECT -20.520 -8.070 -20.350 -8.050 ;
        RECT -19.540 -8.070 -19.370 -7.110 ;
        RECT -18.560 -8.070 -18.390 -7.110 ;
        RECT -18.180 -8.245 -18.010 -6.745 ;
        RECT -17.780 -6.615 -17.610 -5.300 ;
        RECT -17.290 -6.340 -17.120 -5.300 ;
        RECT -16.800 -6.615 -16.630 -5.300 ;
        RECT -16.310 -6.340 -16.140 -5.300 ;
        RECT -15.820 -6.615 -15.650 -5.300 ;
        RECT -15.330 -6.340 -15.160 -5.300 ;
        RECT -14.840 -6.615 -14.670 -5.300 ;
        RECT -14.350 -6.340 -14.180 -5.300 ;
        RECT -13.860 -6.615 -13.690 -5.300 ;
        RECT 36.670 -5.610 37.215 -5.465 ;
        RECT 39.530 -5.610 39.910 -5.310 ;
        RECT 36.670 -5.915 39.910 -5.610 ;
        RECT 40.525 -5.460 40.695 -5.015 ;
        RECT 42.410 -5.460 42.920 -5.220 ;
        RECT 40.525 -5.630 42.920 -5.460 ;
        RECT 45.025 -5.445 45.195 -2.475 ;
        RECT 46.855 -4.515 47.025 -2.475 ;
        RECT 48.035 -4.515 48.205 -2.475 ;
        RECT 49.215 -4.515 49.385 -2.475 ;
        RECT 50.395 -4.515 50.565 -2.475 ;
        RECT 51.575 -4.515 51.745 -2.475 ;
        RECT 52.755 -4.515 52.925 -2.475 ;
        RECT 53.935 -4.515 54.105 -2.475 ;
        RECT 47.215 -5.445 47.575 -5.075 ;
        RECT 45.025 -5.615 47.575 -5.445 ;
        RECT -17.780 -6.785 -13.690 -6.615 ;
        RECT -17.780 -8.070 -17.610 -6.785 ;
        RECT -17.290 -8.070 -17.120 -7.030 ;
        RECT -16.800 -8.070 -16.630 -6.785 ;
        RECT -16.310 -8.070 -16.140 -7.030 ;
        RECT -15.820 -8.070 -15.650 -6.785 ;
        RECT -15.330 -8.070 -15.160 -7.030 ;
        RECT -14.840 -8.070 -14.670 -6.785 ;
        RECT -14.350 -8.070 -14.180 -7.030 ;
        RECT -13.860 -8.070 -13.690 -6.785 ;
        RECT 27.390 -6.800 27.560 -6.340 ;
        RECT 28.370 -6.800 28.540 -6.340 ;
        RECT 29.350 -6.800 29.520 -6.340 ;
        RECT 27.360 -7.265 27.590 -6.800 ;
        RECT 28.340 -7.265 28.570 -6.800 ;
        RECT 29.320 -7.105 29.550 -6.800 ;
        RECT 30.620 -7.050 30.790 -6.010 ;
        RECT 31.600 -7.050 31.770 -6.010 ;
        RECT 32.580 -7.050 32.750 -6.010 ;
        RECT 33.560 -7.050 33.730 -6.010 ;
        RECT 36.670 -6.035 37.215 -5.915 ;
        RECT 39.530 -6.195 39.910 -5.915 ;
        RECT 42.410 -5.920 42.920 -5.630 ;
        RECT 47.215 -5.855 47.575 -5.615 ;
        RECT 55.115 -5.515 55.285 -2.475 ;
        RECT 107.310 -2.610 107.480 -1.295 ;
        RECT 107.800 -2.610 107.970 -1.570 ;
        RECT 108.290 -2.610 108.460 -1.295 ;
        RECT 108.780 -2.610 108.950 -1.570 ;
        RECT 109.270 -2.610 109.440 -1.295 ;
        RECT 109.760 -2.610 109.930 -1.570 ;
        RECT 110.250 -2.610 110.420 -1.295 ;
        RECT 110.740 -2.610 110.910 -1.570 ;
        RECT 111.230 -2.610 111.400 -1.295 ;
        RECT 254.055 -1.405 254.225 0.635 ;
        RECT 255.235 -1.735 255.405 0.635 ;
        RECT 257.065 -1.405 257.235 0.635 ;
        RECT 258.245 -1.405 258.415 0.635 ;
        RECT 259.425 -1.405 259.595 0.635 ;
        RECT 255.235 -1.905 256.275 -1.735 ;
        RECT 252.170 -2.500 253.625 -2.390 ;
        RECT 255.110 -2.500 255.490 -2.200 ;
        RECT 252.170 -2.805 255.490 -2.500 ;
        RECT 256.105 -2.350 256.275 -1.905 ;
        RECT 257.990 -2.350 258.500 -2.110 ;
        RECT 256.105 -2.520 258.500 -2.350 ;
        RECT 260.605 -2.335 260.775 0.635 ;
        RECT 262.435 -1.405 262.605 0.635 ;
        RECT 263.615 -1.405 263.785 0.635 ;
        RECT 264.795 -1.405 264.965 0.635 ;
        RECT 265.975 -1.405 266.145 0.635 ;
        RECT 267.155 -1.405 267.325 0.635 ;
        RECT 268.335 -1.405 268.505 0.635 ;
        RECT 269.515 -1.405 269.685 0.635 ;
        RECT 262.795 -2.335 263.155 -1.965 ;
        RECT 260.605 -2.505 263.155 -2.335 ;
        RECT 252.170 -2.860 253.625 -2.805 ;
        RECT 238.790 -3.160 253.625 -2.860 ;
        RECT 255.110 -3.085 255.490 -2.805 ;
        RECT 257.990 -2.810 258.500 -2.520 ;
        RECT 262.795 -2.745 263.155 -2.505 ;
        RECT 270.695 -2.405 270.865 0.635 ;
        RECT 272.235 -2.405 272.595 -2.135 ;
        RECT 270.695 -2.575 272.595 -2.405 ;
        RECT 272.235 -2.915 272.595 -2.575 ;
        RECT 104.570 -4.275 104.740 -3.815 ;
        RECT 105.550 -4.275 105.720 -3.815 ;
        RECT 106.530 -4.275 106.700 -3.815 ;
        RECT 104.540 -4.740 104.770 -4.275 ;
        RECT 105.520 -4.740 105.750 -4.275 ;
        RECT 106.500 -4.580 106.730 -4.275 ;
        RECT 107.800 -4.525 107.970 -3.485 ;
        RECT 108.780 -4.525 108.950 -3.485 ;
        RECT 109.760 -4.525 109.930 -3.485 ;
        RECT 110.740 -4.525 110.910 -3.485 ;
        RECT 238.790 -3.630 252.940 -3.160 ;
        RECT 238.790 -3.760 239.765 -3.630 ;
        RECT 106.500 -4.740 107.080 -4.580 ;
        RECT 104.540 -4.930 107.080 -4.740 ;
        RECT 104.540 -4.970 106.730 -4.930 ;
        RECT 56.655 -5.515 57.015 -5.245 ;
        RECT 55.115 -5.685 57.015 -5.515 ;
        RECT 56.655 -6.025 57.015 -5.685 ;
        RECT 104.540 -6.235 104.770 -4.970 ;
        RECT 105.520 -5.295 105.750 -4.970 ;
        RECT 106.500 -5.295 106.730 -4.970 ;
        RECT 104.570 -6.255 104.740 -6.235 ;
        RECT 105.550 -6.255 105.720 -5.295 ;
        RECT 106.530 -6.255 106.700 -5.295 ;
        RECT 106.910 -6.430 107.080 -4.930 ;
        RECT 107.800 -6.255 107.970 -5.215 ;
        RECT 108.780 -6.255 108.950 -5.215 ;
        RECT 109.760 -6.255 109.930 -5.215 ;
        RECT 110.740 -6.255 110.910 -5.215 ;
        RECT 255.515 -5.445 255.685 -3.405 ;
        RECT 256.695 -5.445 256.865 -3.405 ;
        RECT 257.875 -5.445 258.045 -3.405 ;
        RECT 259.055 -5.445 259.225 -3.405 ;
        RECT 260.235 -5.445 260.405 -3.405 ;
        RECT 261.415 -5.445 261.585 -3.405 ;
        RECT 262.595 -5.445 262.765 -3.405 ;
        RECT 29.320 -7.265 29.900 -7.105 ;
        RECT 27.360 -7.455 29.900 -7.265 ;
        RECT 27.360 -7.495 29.550 -7.455 ;
        RECT -18.180 -8.415 -16.710 -8.245 ;
        RECT -17.550 -8.615 -16.710 -8.415 ;
        RECT 27.360 -8.760 27.590 -7.495 ;
        RECT 28.340 -7.820 28.570 -7.495 ;
        RECT 29.320 -7.820 29.550 -7.495 ;
        RECT 27.390 -8.780 27.560 -8.760 ;
        RECT 28.370 -8.780 28.540 -7.820 ;
        RECT 29.350 -8.780 29.520 -7.820 ;
        RECT 29.730 -8.955 29.900 -7.455 ;
        RECT 30.620 -8.780 30.790 -7.740 ;
        RECT 31.600 -8.780 31.770 -7.740 ;
        RECT 32.580 -8.780 32.750 -7.740 ;
        RECT 33.560 -8.780 33.730 -7.740 ;
        RECT 39.935 -8.555 40.105 -6.515 ;
        RECT 41.115 -8.555 41.285 -6.515 ;
        RECT 42.295 -8.555 42.465 -6.515 ;
        RECT 43.475 -8.555 43.645 -6.515 ;
        RECT 44.655 -8.555 44.825 -6.515 ;
        RECT 45.835 -8.555 46.005 -6.515 ;
        RECT 47.015 -8.555 47.185 -6.515 ;
        RECT 106.910 -6.600 108.380 -6.430 ;
        RECT 107.540 -6.800 108.380 -6.600 ;
        RECT 29.730 -9.125 31.200 -8.955 ;
        RECT 30.360 -9.325 31.200 -9.125 ;
        RECT 319.675 -13.825 320.515 -13.625 ;
        RECT 319.045 -13.995 320.515 -13.825 ;
        RECT 312.455 -14.190 312.625 -14.170 ;
        RECT 254.055 -16.640 254.225 -14.600 ;
        RECT 244.830 -17.735 246.385 -16.855 ;
        RECT 255.235 -16.970 255.405 -14.600 ;
        RECT 257.065 -16.640 257.235 -14.600 ;
        RECT 258.245 -16.640 258.415 -14.600 ;
        RECT 259.425 -16.640 259.595 -14.600 ;
        RECT 255.235 -17.140 256.275 -16.970 ;
        RECT 255.110 -17.735 255.490 -17.435 ;
        RECT 244.830 -18.040 255.490 -17.735 ;
        RECT 256.105 -17.585 256.275 -17.140 ;
        RECT 257.990 -17.585 258.500 -17.345 ;
        RECT 256.105 -17.755 258.500 -17.585 ;
        RECT 260.605 -17.570 260.775 -14.600 ;
        RECT 262.435 -16.640 262.605 -14.600 ;
        RECT 263.615 -16.640 263.785 -14.600 ;
        RECT 264.795 -16.640 264.965 -14.600 ;
        RECT 265.975 -16.640 266.145 -14.600 ;
        RECT 267.155 -16.640 267.325 -14.600 ;
        RECT 268.335 -16.640 268.505 -14.600 ;
        RECT 269.515 -16.640 269.685 -14.600 ;
        RECT 262.795 -17.570 263.155 -17.200 ;
        RECT 260.605 -17.740 263.155 -17.570 ;
        RECT 244.830 -18.485 246.385 -18.040 ;
        RECT 255.110 -18.320 255.490 -18.040 ;
        RECT 257.990 -18.045 258.500 -17.755 ;
        RECT 262.795 -17.980 263.155 -17.740 ;
        RECT 270.695 -17.640 270.865 -14.600 ;
        RECT 271.935 -16.640 272.105 -14.600 ;
        RECT 273.115 -16.640 273.285 -14.600 ;
        RECT 274.295 -16.640 274.465 -14.600 ;
        RECT 275.475 -16.640 275.645 -14.600 ;
        RECT 276.655 -16.640 276.825 -14.600 ;
        RECT 277.835 -16.640 278.005 -14.600 ;
        RECT 279.015 -16.640 279.185 -14.600 ;
        RECT 280.195 -16.640 280.365 -14.600 ;
        RECT 281.375 -16.640 281.545 -14.600 ;
        RECT 282.555 -16.640 282.725 -14.600 ;
        RECT 283.735 -16.640 283.905 -14.600 ;
        RECT 284.915 -16.640 285.085 -14.600 ;
        RECT 286.095 -16.640 286.265 -14.600 ;
        RECT 287.275 -16.640 287.445 -14.600 ;
        RECT 288.455 -16.640 288.625 -14.600 ;
        RECT 289.635 -16.640 289.805 -14.600 ;
        RECT 290.815 -17.160 290.985 -14.600 ;
        RECT 312.425 -15.455 312.655 -14.190 ;
        RECT 313.435 -15.130 313.605 -14.170 ;
        RECT 314.415 -15.130 314.585 -14.170 ;
        RECT 316.705 -14.190 316.875 -14.170 ;
        RECT 313.405 -15.455 313.635 -15.130 ;
        RECT 314.385 -15.455 314.615 -15.130 ;
        RECT 312.425 -15.495 314.615 -15.455 ;
        RECT 316.675 -15.455 316.905 -14.190 ;
        RECT 317.685 -15.130 317.855 -14.170 ;
        RECT 318.665 -15.130 318.835 -14.170 ;
        RECT 317.655 -15.455 317.885 -15.130 ;
        RECT 318.635 -15.455 318.865 -15.130 ;
        RECT 316.675 -15.495 318.865 -15.455 ;
        RECT 319.045 -15.495 319.215 -13.995 ;
        RECT 312.425 -15.570 315.445 -15.495 ;
        RECT 315.655 -15.570 316.495 -15.530 ;
        RECT 312.425 -15.685 316.495 -15.570 ;
        RECT 312.425 -16.150 312.655 -15.685 ;
        RECT 313.405 -16.150 313.635 -15.685 ;
        RECT 314.385 -15.830 316.495 -15.685 ;
        RECT 314.385 -15.845 315.445 -15.830 ;
        RECT 314.385 -16.150 314.615 -15.845 ;
        RECT 315.655 -15.900 316.495 -15.830 ;
        RECT 316.675 -15.685 319.215 -15.495 ;
        RECT 316.675 -16.150 316.905 -15.685 ;
        RECT 317.655 -16.150 317.885 -15.685 ;
        RECT 318.635 -15.845 319.215 -15.685 ;
        RECT 319.445 -15.455 319.615 -14.170 ;
        RECT 319.935 -15.210 320.105 -14.170 ;
        RECT 320.425 -15.455 320.595 -14.170 ;
        RECT 320.915 -15.210 321.085 -14.170 ;
        RECT 321.405 -15.455 321.575 -14.170 ;
        RECT 321.895 -15.210 322.065 -14.170 ;
        RECT 322.385 -15.455 322.555 -14.170 ;
        RECT 322.875 -15.210 323.045 -14.170 ;
        RECT 323.365 -15.455 323.535 -14.170 ;
        RECT 319.445 -15.625 323.535 -15.455 ;
        RECT 318.635 -16.150 318.865 -15.845 ;
        RECT 312.455 -16.610 312.625 -16.150 ;
        RECT 313.435 -16.610 313.605 -16.150 ;
        RECT 314.415 -16.610 314.585 -16.150 ;
        RECT 316.705 -16.610 316.875 -16.150 ;
        RECT 317.685 -16.610 317.855 -16.150 ;
        RECT 318.665 -16.610 318.835 -16.150 ;
        RECT 319.445 -16.940 319.615 -15.625 ;
        RECT 319.935 -16.940 320.105 -15.900 ;
        RECT 320.425 -16.940 320.595 -15.625 ;
        RECT 320.915 -16.940 321.085 -15.900 ;
        RECT 321.405 -16.940 321.575 -15.625 ;
        RECT 321.895 -16.940 322.065 -15.900 ;
        RECT 322.385 -16.940 322.555 -15.625 ;
        RECT 322.875 -16.940 323.045 -15.900 ;
        RECT 323.365 -16.940 323.535 -15.625 ;
        RECT 438.925 -16.440 441.050 -15.945 ;
        RECT 309.365 -17.160 310.335 -17.035 ;
        RECT 290.815 -17.370 310.335 -17.160 ;
        RECT 272.235 -17.640 272.595 -17.370 ;
        RECT 290.815 -17.540 310.480 -17.370 ;
        RECT 325.635 -17.535 441.050 -16.440 ;
        RECT 309.365 -17.580 310.335 -17.540 ;
        RECT 270.695 -17.810 272.595 -17.640 ;
        RECT 272.235 -18.150 272.595 -17.810 ;
        RECT 316.705 -18.605 316.875 -18.145 ;
        RECT 317.685 -18.605 317.855 -18.145 ;
        RECT 318.665 -18.605 318.835 -18.145 ;
        RECT 255.515 -20.680 255.685 -18.640 ;
        RECT 256.695 -20.680 256.865 -18.640 ;
        RECT 257.875 -20.680 258.045 -18.640 ;
        RECT 259.055 -20.680 259.225 -18.640 ;
        RECT 260.235 -20.680 260.405 -18.640 ;
        RECT 261.415 -20.680 261.585 -18.640 ;
        RECT 262.595 -20.680 262.765 -18.640 ;
        RECT 263.775 -20.680 263.945 -18.640 ;
        RECT 264.955 -20.680 265.125 -18.640 ;
        RECT 266.135 -20.680 266.305 -18.640 ;
        RECT 267.315 -20.680 267.485 -18.640 ;
        RECT 268.495 -20.680 268.665 -18.640 ;
        RECT 269.675 -20.680 269.845 -18.640 ;
        RECT 270.855 -20.680 271.025 -18.640 ;
        RECT 272.035 -20.680 272.205 -18.640 ;
        RECT 316.675 -19.070 316.905 -18.605 ;
        RECT 317.655 -19.070 317.885 -18.605 ;
        RECT 318.635 -18.910 318.865 -18.605 ;
        RECT 319.935 -18.855 320.105 -17.815 ;
        RECT 320.915 -18.855 321.085 -17.815 ;
        RECT 321.895 -18.855 322.065 -17.815 ;
        RECT 322.875 -18.855 323.045 -17.815 ;
        RECT 438.925 -17.905 441.050 -17.535 ;
        RECT 318.635 -19.070 319.215 -18.910 ;
        RECT 316.675 -19.260 319.215 -19.070 ;
        RECT 316.675 -19.300 318.865 -19.260 ;
        RECT 316.675 -20.565 316.905 -19.300 ;
        RECT 317.655 -19.625 317.885 -19.300 ;
        RECT 318.635 -19.625 318.865 -19.300 ;
        RECT 316.705 -20.585 316.875 -20.565 ;
        RECT 317.685 -20.585 317.855 -19.625 ;
        RECT 318.665 -20.585 318.835 -19.625 ;
        RECT 319.045 -20.760 319.215 -19.260 ;
        RECT 319.935 -20.585 320.105 -19.545 ;
        RECT 320.915 -20.585 321.085 -19.545 ;
        RECT 321.895 -20.585 322.065 -19.545 ;
        RECT 322.875 -20.585 323.045 -19.545 ;
        RECT 319.045 -20.930 320.515 -20.760 ;
        RECT 319.675 -21.130 320.515 -20.930 ;
        RECT -134.535 -55.440 -129.915 -54.900 ;
        RECT -121.865 -55.440 -116.390 -54.795 ;
        RECT -134.535 -58.660 -116.390 -55.440 ;
        RECT -134.535 -59.520 -129.915 -58.660 ;
        RECT -121.865 -59.200 -116.390 -58.660 ;
        RECT -129.655 -70.940 -124.350 -70.540 ;
        RECT -129.655 -74.040 -35.925 -70.940 ;
        RECT -129.655 -74.380 -124.350 -74.040 ;
        RECT -64.370 -75.595 -39.350 -74.845 ;
        RECT -74.910 -76.195 -38.975 -75.595 ;
        RECT -74.755 -78.660 -74.585 -76.620 ;
        RECT -74.165 -78.660 -73.995 -76.620 ;
        RECT -73.575 -78.660 -73.405 -76.620 ;
        RECT -72.985 -78.660 -72.815 -76.620 ;
        RECT -72.395 -78.660 -72.225 -76.620 ;
        RECT -71.805 -78.660 -71.635 -76.620 ;
        RECT -71.215 -78.660 -71.045 -76.620 ;
        RECT -70.625 -78.660 -70.455 -76.620 ;
        RECT -70.035 -78.660 -69.865 -76.620 ;
        RECT -69.445 -78.660 -69.275 -76.620 ;
        RECT -68.855 -78.660 -68.685 -76.620 ;
        RECT -68.265 -78.660 -68.095 -76.620 ;
        RECT -67.675 -78.660 -67.505 -76.620 ;
        RECT -67.085 -78.660 -66.915 -76.620 ;
        RECT -66.495 -78.660 -66.325 -76.620 ;
        RECT -65.905 -78.660 -65.735 -76.620 ;
        RECT -65.315 -78.660 -65.145 -76.620 ;
        RECT -64.725 -78.660 -64.555 -76.620 ;
        RECT -64.135 -78.660 -63.965 -76.620 ;
        RECT -63.545 -78.660 -63.375 -76.620 ;
        RECT -62.955 -78.660 -62.785 -76.620 ;
        RECT -62.365 -78.660 -62.195 -76.620 ;
        RECT -61.775 -78.660 -61.605 -76.620 ;
        RECT -61.185 -78.660 -61.015 -76.620 ;
        RECT -60.595 -78.660 -60.425 -76.620 ;
        RECT -60.005 -78.660 -59.835 -76.620 ;
        RECT -59.415 -78.660 -59.245 -76.620 ;
        RECT -58.825 -78.660 -58.655 -76.620 ;
        RECT -58.235 -78.660 -58.065 -76.620 ;
        RECT -57.645 -78.660 -57.475 -76.620 ;
        RECT -57.055 -78.660 -56.885 -76.195 ;
        RECT -55.875 -78.660 -55.705 -76.195 ;
        RECT -54.695 -78.660 -54.525 -76.195 ;
        RECT -53.515 -78.660 -53.345 -76.195 ;
        RECT -52.335 -78.660 -52.165 -76.195 ;
        RECT -51.155 -78.660 -50.985 -76.195 ;
        RECT -49.975 -78.660 -49.805 -76.195 ;
        RECT -48.795 -78.660 -48.625 -76.195 ;
        RECT -47.615 -78.660 -47.445 -76.195 ;
        RECT -47.025 -78.660 -46.855 -76.620 ;
        RECT -46.435 -78.660 -46.265 -76.195 ;
        RECT -45.845 -78.660 -45.675 -76.620 ;
        RECT -45.255 -78.660 -45.085 -76.195 ;
        RECT -44.665 -78.660 -44.495 -76.620 ;
        RECT -44.075 -78.660 -43.905 -76.195 ;
        RECT -43.485 -78.660 -43.315 -76.620 ;
        RECT -42.895 -78.660 -42.725 -76.195 ;
        RECT -42.305 -78.660 -42.135 -76.620 ;
        RECT -41.715 -78.660 -41.545 -76.195 ;
        RECT -41.125 -78.660 -40.955 -76.620 ;
        RECT -40.535 -78.660 -40.365 -76.195 ;
        RECT -39.945 -78.660 -39.775 -76.620 ;
        RECT -39.355 -78.660 -39.185 -76.195 ;
        RECT -74.885 -78.980 -56.735 -78.660 ;
        RECT -74.885 -79.120 -57.475 -78.980 ;
        RECT -56.855 -79.490 -56.495 -79.150 ;
        RECT -56.855 -79.660 -54.955 -79.490 ;
        RECT -56.855 -79.930 -56.495 -79.660 ;
        RECT -55.125 -82.700 -54.955 -79.660 ;
        RECT -47.415 -79.560 -47.055 -79.320 ;
        RECT -42.760 -79.545 -42.250 -79.255 ;
        RECT -39.750 -79.260 -39.370 -78.980 ;
        RECT -37.680 -79.260 -35.925 -74.040 ;
        RECT -47.415 -79.730 -44.865 -79.560 ;
        RECT -47.415 -80.100 -47.055 -79.730 ;
        RECT -53.945 -82.700 -53.775 -80.660 ;
        RECT -52.765 -82.700 -52.595 -80.660 ;
        RECT -51.585 -82.700 -51.415 -80.660 ;
        RECT -50.405 -82.700 -50.235 -80.660 ;
        RECT -49.225 -82.700 -49.055 -80.660 ;
        RECT -48.045 -82.700 -47.875 -80.660 ;
        RECT -46.865 -82.700 -46.695 -80.660 ;
        RECT -45.035 -82.700 -44.865 -79.730 ;
        RECT -42.760 -79.715 -40.365 -79.545 ;
        RECT -42.760 -79.955 -42.250 -79.715 ;
        RECT -40.535 -80.160 -40.365 -79.715 ;
        RECT -39.750 -79.565 -35.925 -79.260 ;
        RECT -39.750 -79.865 -39.370 -79.565 ;
        RECT -40.535 -80.330 -39.495 -80.160 ;
        RECT -43.855 -82.700 -43.685 -80.660 ;
        RECT -42.675 -82.700 -42.505 -80.660 ;
        RECT -41.495 -82.700 -41.325 -80.660 ;
        RECT -39.665 -82.700 -39.495 -80.330 ;
        RECT -38.485 -82.700 -38.315 -80.660 ;
        RECT 37.715 -88.055 94.055 -86.390 ;
        RECT -67.970 -91.870 -64.830 -91.700 ;
        RECT -75.205 -91.985 -75.035 -91.965 ;
        RECT -75.235 -93.250 -75.005 -91.985 ;
        RECT -74.225 -92.925 -74.055 -91.965 ;
        RECT -73.245 -92.925 -73.075 -91.965 ;
        RECT -71.020 -91.985 -70.850 -91.965 ;
        RECT -72.125 -92.395 -71.840 -92.075 ;
        RECT -72.840 -92.640 -71.840 -92.395 ;
        RECT -74.255 -93.250 -74.025 -92.925 ;
        RECT -73.275 -93.250 -73.045 -92.925 ;
        RECT -75.235 -93.290 -73.045 -93.250 ;
        RECT -72.840 -93.290 -72.610 -92.640 ;
        RECT -72.125 -92.895 -71.840 -92.640 ;
        RECT -76.255 -93.475 -75.415 -93.325 ;
        RECT -76.290 -93.695 -75.415 -93.475 ;
        RECT -75.235 -93.480 -72.610 -93.290 ;
        RECT -71.050 -93.250 -70.820 -91.985 ;
        RECT -70.040 -92.925 -69.870 -91.965 ;
        RECT -69.060 -92.925 -68.890 -91.965 ;
        RECT -67.970 -92.095 -67.790 -91.870 ;
        RECT -70.070 -93.250 -69.840 -92.925 ;
        RECT -69.090 -93.250 -68.860 -92.925 ;
        RECT -71.050 -93.290 -68.860 -93.250 ;
        RECT -68.585 -93.170 -68.215 -92.330 ;
        RECT -67.965 -92.465 -67.795 -92.095 ;
        RECT -68.585 -93.290 -68.220 -93.170 ;
        RECT -72.070 -93.380 -71.230 -93.325 ;
        RECT -72.245 -93.385 -71.230 -93.380 ;
        RECT -76.290 -95.555 -76.050 -93.695 ;
        RECT -75.695 -94.660 -75.525 -93.865 ;
        RECT -75.235 -93.945 -75.005 -93.480 ;
        RECT -75.205 -94.405 -75.035 -93.945 ;
        RECT -74.715 -94.660 -74.545 -93.865 ;
        RECT -74.255 -93.945 -74.025 -93.480 ;
        RECT -73.275 -93.640 -72.610 -93.480 ;
        RECT -74.225 -94.405 -74.055 -93.945 ;
        RECT -73.735 -94.660 -73.565 -93.865 ;
        RECT -73.275 -93.945 -73.045 -93.640 ;
        RECT -72.430 -93.695 -71.230 -93.385 ;
        RECT -71.050 -93.480 -68.220 -93.290 ;
        RECT -73.245 -94.405 -73.075 -93.945 ;
        RECT -72.430 -94.415 -72.130 -93.695 ;
        RECT -71.510 -94.660 -71.340 -93.865 ;
        RECT -71.050 -93.945 -70.820 -93.480 ;
        RECT -71.020 -94.405 -70.850 -93.945 ;
        RECT -70.530 -94.660 -70.360 -93.865 ;
        RECT -70.070 -93.945 -69.840 -93.480 ;
        RECT -69.090 -93.640 -68.220 -93.480 ;
        RECT -67.995 -93.200 -67.760 -92.465 ;
        RECT -67.475 -92.500 -67.305 -92.040 ;
        RECT -66.990 -92.145 -66.780 -91.870 ;
        RECT -67.480 -92.760 -67.300 -92.500 ;
        RECT -66.985 -92.580 -66.815 -92.145 ;
        RECT -66.495 -92.490 -66.325 -92.040 ;
        RECT -66.020 -92.150 -65.810 -91.870 ;
        RECT -66.495 -92.580 -66.310 -92.490 ;
        RECT -66.005 -92.580 -65.835 -92.150 ;
        RECT -65.515 -92.490 -65.345 -92.040 ;
        RECT -65.040 -92.125 -64.830 -91.870 ;
        RECT -54.470 -91.870 -51.330 -91.700 ;
        RECT -61.705 -91.985 -61.535 -91.965 ;
        RECT -66.490 -92.760 -66.310 -92.580 ;
        RECT -65.520 -92.760 -65.340 -92.490 ;
        RECT -65.025 -92.580 -64.855 -92.125 ;
        RECT -64.535 -92.540 -64.365 -92.040 ;
        RECT -64.550 -92.760 -64.340 -92.540 ;
        RECT -67.480 -92.930 -64.340 -92.760 ;
        RECT -67.995 -93.570 -67.135 -93.200 ;
        RECT -65.215 -93.465 -64.340 -92.930 ;
        RECT -61.735 -93.250 -61.505 -91.985 ;
        RECT -60.725 -92.925 -60.555 -91.965 ;
        RECT -59.745 -92.925 -59.575 -91.965 ;
        RECT -57.520 -91.985 -57.350 -91.965 ;
        RECT -58.625 -92.335 -58.340 -92.075 ;
        RECT -59.365 -92.645 -58.340 -92.335 ;
        RECT -60.755 -93.250 -60.525 -92.925 ;
        RECT -59.775 -93.250 -59.545 -92.925 ;
        RECT -61.735 -93.290 -59.545 -93.250 ;
        RECT -59.365 -93.290 -59.055 -92.645 ;
        RECT -58.625 -92.895 -58.340 -92.645 ;
        RECT -62.755 -93.360 -61.915 -93.325 ;
        RECT -70.040 -94.405 -69.870 -93.945 ;
        RECT -69.550 -94.660 -69.380 -93.865 ;
        RECT -69.090 -93.945 -68.860 -93.640 ;
        RECT -69.060 -94.405 -68.890 -93.945 ;
        RECT -67.995 -94.245 -67.760 -93.570 ;
        RECT -65.215 -93.765 -63.885 -93.465 ;
        RECT -62.865 -93.660 -61.915 -93.360 ;
        RECT -62.755 -93.695 -61.915 -93.660 ;
        RECT -61.735 -93.480 -59.055 -93.290 ;
        RECT -57.550 -93.250 -57.320 -91.985 ;
        RECT -56.540 -92.925 -56.370 -91.965 ;
        RECT -55.560 -92.925 -55.390 -91.965 ;
        RECT -54.470 -92.095 -54.290 -91.870 ;
        RECT -56.570 -93.250 -56.340 -92.925 ;
        RECT -55.590 -93.250 -55.360 -92.925 ;
        RECT -57.550 -93.290 -55.360 -93.250 ;
        RECT -55.085 -93.170 -54.715 -92.330 ;
        RECT -54.465 -92.465 -54.295 -92.095 ;
        RECT -55.085 -93.290 -54.720 -93.170 ;
        RECT -58.570 -93.380 -57.730 -93.325 ;
        RECT -67.495 -93.935 -64.340 -93.765 ;
        RECT -67.495 -94.140 -67.290 -93.935 ;
        RECT -67.965 -94.595 -67.795 -94.245 ;
        RECT -75.740 -95.000 -68.885 -94.660 ;
        RECT -67.990 -94.885 -67.770 -94.595 ;
        RECT -67.475 -94.655 -67.305 -94.140 ;
        RECT -66.985 -94.540 -66.815 -94.115 ;
        RECT -66.505 -94.180 -66.300 -93.935 ;
        RECT -67.010 -94.885 -66.790 -94.540 ;
        RECT -66.495 -94.655 -66.325 -94.180 ;
        RECT -66.005 -94.540 -65.835 -94.115 ;
        RECT -65.535 -94.180 -65.330 -93.935 ;
        RECT -64.550 -93.970 -64.340 -93.935 ;
        RECT -66.030 -94.885 -65.810 -94.540 ;
        RECT -65.515 -94.655 -65.345 -94.180 ;
        RECT -65.025 -94.595 -64.855 -94.115 ;
        RECT -64.550 -94.185 -64.345 -93.970 ;
        RECT -65.045 -94.885 -64.825 -94.595 ;
        RECT -64.535 -94.655 -64.365 -94.185 ;
        RECT -62.195 -94.660 -62.025 -93.865 ;
        RECT -61.735 -93.945 -61.505 -93.480 ;
        RECT -61.705 -94.405 -61.535 -93.945 ;
        RECT -61.215 -94.660 -61.045 -93.865 ;
        RECT -60.755 -93.945 -60.525 -93.480 ;
        RECT -59.775 -93.640 -59.055 -93.480 ;
        RECT -60.725 -94.405 -60.555 -93.945 ;
        RECT -60.235 -94.660 -60.065 -93.865 ;
        RECT -59.775 -93.945 -59.545 -93.640 ;
        RECT -58.870 -93.695 -57.730 -93.380 ;
        RECT -57.550 -93.480 -54.720 -93.290 ;
        RECT -59.745 -94.405 -59.575 -93.945 ;
        RECT -58.870 -94.490 -58.570 -93.695 ;
        RECT -58.010 -94.660 -57.840 -93.865 ;
        RECT -57.550 -93.945 -57.320 -93.480 ;
        RECT -57.520 -94.405 -57.350 -93.945 ;
        RECT -57.030 -94.660 -56.860 -93.865 ;
        RECT -56.570 -93.945 -56.340 -93.480 ;
        RECT -55.590 -93.640 -54.720 -93.480 ;
        RECT -54.495 -93.200 -54.260 -92.465 ;
        RECT -53.975 -92.500 -53.805 -92.040 ;
        RECT -53.490 -92.145 -53.280 -91.870 ;
        RECT -53.980 -92.760 -53.800 -92.500 ;
        RECT -53.485 -92.580 -53.315 -92.145 ;
        RECT -52.995 -92.490 -52.825 -92.040 ;
        RECT -52.520 -92.150 -52.310 -91.870 ;
        RECT -52.995 -92.580 -52.810 -92.490 ;
        RECT -52.505 -92.580 -52.335 -92.150 ;
        RECT -52.015 -92.490 -51.845 -92.040 ;
        RECT -51.540 -92.125 -51.330 -91.870 ;
        RECT -43.345 -91.845 -42.145 -91.675 ;
        RECT -52.990 -92.760 -52.810 -92.580 ;
        RECT -52.020 -92.760 -51.840 -92.490 ;
        RECT -51.525 -92.580 -51.355 -92.125 ;
        RECT -51.035 -92.540 -50.865 -92.040 ;
        RECT -51.050 -92.760 -50.840 -92.540 ;
        RECT -53.980 -92.930 -50.840 -92.760 ;
        RECT -54.495 -93.570 -53.635 -93.200 ;
        RECT -51.715 -93.475 -50.840 -92.930 ;
        RECT -56.540 -94.405 -56.370 -93.945 ;
        RECT -56.050 -94.660 -55.880 -93.865 ;
        RECT -55.590 -93.945 -55.360 -93.640 ;
        RECT -55.560 -94.405 -55.390 -93.945 ;
        RECT -54.495 -94.245 -54.260 -93.570 ;
        RECT -51.715 -93.765 -50.465 -93.475 ;
        RECT -53.995 -93.775 -50.465 -93.765 ;
        RECT -53.995 -93.935 -50.840 -93.775 ;
        RECT -53.995 -94.140 -53.790 -93.935 ;
        RECT -54.465 -94.595 -54.295 -94.245 ;
        RECT -74.500 -95.200 -73.945 -95.000 ;
        RECT -74.555 -95.240 -73.870 -95.200 ;
        RECT -70.445 -95.240 -69.890 -95.000 ;
        RECT -67.990 -95.055 -64.825 -94.885 ;
        RECT -62.240 -94.670 -59.570 -94.660 ;
        RECT -58.055 -94.670 -55.385 -94.660 ;
        RECT -62.240 -95.000 -55.385 -94.670 ;
        RECT -54.490 -94.885 -54.270 -94.595 ;
        RECT -53.975 -94.655 -53.805 -94.140 ;
        RECT -53.485 -94.540 -53.315 -94.115 ;
        RECT -53.005 -94.180 -52.800 -93.935 ;
        RECT -53.510 -94.885 -53.290 -94.540 ;
        RECT -52.995 -94.655 -52.825 -94.180 ;
        RECT -52.505 -94.540 -52.335 -94.115 ;
        RECT -52.035 -94.180 -51.830 -93.935 ;
        RECT -51.050 -93.970 -50.840 -93.935 ;
        RECT -52.530 -94.885 -52.310 -94.540 ;
        RECT -52.015 -94.655 -51.845 -94.180 ;
        RECT -51.525 -94.595 -51.355 -94.115 ;
        RECT -51.050 -94.185 -50.845 -93.970 ;
        RECT -51.545 -94.885 -51.325 -94.595 ;
        RECT -51.035 -94.655 -50.865 -94.185 ;
        RECT -61.455 -95.230 -60.900 -95.000 ;
        RECT -60.540 -95.010 -57.940 -95.000 ;
        RECT -61.570 -95.240 -60.885 -95.230 ;
        RECT -57.065 -95.240 -56.510 -95.000 ;
        RECT -54.490 -95.055 -51.325 -94.885 ;
        RECT -44.375 -94.985 -44.205 -92.015 ;
        RECT -43.345 -92.065 -43.135 -91.845 ;
        RECT -48.380 -95.240 -47.720 -95.230 ;
        RECT -74.640 -95.435 -47.715 -95.240 ;
        RECT -74.555 -95.500 -73.870 -95.435 ;
        RECT -61.570 -95.530 -60.885 -95.435 ;
        RECT -48.380 -95.530 -47.720 -95.435 ;
        RECT -113.200 -97.120 -113.030 -95.900 ;
        RECT -112.220 -97.120 -112.050 -95.900 ;
        RECT -111.240 -97.120 -111.070 -95.900 ;
        RECT -113.200 -97.305 -110.425 -97.120 ;
        RECT -110.610 -97.995 -110.425 -97.305 ;
        RECT -108.400 -97.995 -107.725 -97.945 ;
        RECT -110.610 -98.180 -107.725 -97.995 ;
        RECT -110.610 -98.450 -110.425 -98.180 ;
        RECT -108.400 -98.215 -107.725 -98.180 ;
        RECT -113.690 -98.620 -111.475 -98.450 ;
        RECT -110.610 -98.620 -109.445 -98.450 ;
        RECT -113.690 -100.475 -113.520 -98.620 ;
        RECT -112.710 -98.625 -111.475 -98.620 ;
        RECT -113.200 -101.420 -113.030 -98.935 ;
        RECT -112.710 -100.475 -112.540 -98.625 ;
        RECT -111.650 -98.940 -111.475 -98.625 ;
        RECT -112.140 -100.435 -111.970 -98.940 ;
        RECT -112.140 -100.955 -111.965 -100.435 ;
        RECT -111.650 -100.480 -111.480 -98.940 ;
        RECT -111.160 -100.425 -110.990 -98.940 ;
        RECT -111.160 -100.955 -110.985 -100.425 ;
        RECT -110.595 -100.480 -110.425 -98.620 ;
        RECT -112.140 -100.970 -110.985 -100.955 ;
        RECT -110.105 -100.970 -109.935 -98.940 ;
        RECT -109.615 -100.480 -109.445 -98.620 ;
        RECT -112.140 -101.140 -109.935 -100.970 ;
        RECT -108.040 -100.975 -107.870 -99.440 ;
        RECT -107.550 -100.480 -107.380 -95.900 ;
        RECT -103.205 -98.230 -103.035 -96.510 ;
        RECT -102.225 -98.230 -102.055 -96.510 ;
        RECT -100.160 -97.045 -99.990 -96.505 ;
        RECT -99.180 -97.045 -99.010 -96.505 ;
        RECT -100.750 -97.280 -100.385 -97.215 ;
        RECT -101.250 -97.420 -100.385 -97.280 ;
        RECT -101.360 -97.485 -100.385 -97.420 ;
        RECT -101.360 -98.230 -101.055 -97.485 ;
        RECT -100.750 -97.515 -100.385 -97.485 ;
        RECT -98.200 -97.365 -98.030 -96.505 ;
        RECT -91.460 -96.685 -84.075 -96.120 ;
        RECT -76.295 -96.240 -75.995 -95.555 ;
        RECT -63.745 -95.700 -63.060 -95.645 ;
        RECT -59.015 -95.700 -58.355 -95.650 ;
        RECT -74.640 -95.895 -45.990 -95.700 ;
        RECT -63.745 -95.945 -63.060 -95.895 ;
        RECT -59.015 -95.950 -58.355 -95.895 ;
        RECT -72.610 -96.130 -71.950 -96.090 ;
        RECT -49.995 -96.130 -49.335 -96.080 ;
        RECT -98.200 -97.370 -96.180 -97.365 ;
        RECT -98.200 -97.660 -95.860 -97.370 ;
        RECT -103.205 -98.380 -101.055 -98.230 ;
        RECT -103.205 -98.420 -101.110 -98.380 ;
        RECT -100.160 -98.440 -99.990 -97.660 ;
        RECT -99.670 -98.200 -99.500 -97.660 ;
        RECT -99.180 -98.440 -99.010 -97.660 ;
        RECT -98.690 -98.200 -98.520 -97.660 ;
        RECT -98.200 -97.715 -96.180 -97.660 ;
        RECT -95.615 -98.160 -93.370 -98.070 ;
        RECT -91.460 -98.160 -91.155 -96.685 ;
        RECT -87.825 -97.275 -87.590 -96.685 ;
        RECT -97.995 -98.440 -91.155 -98.160 ;
        RECT -100.860 -98.465 -91.155 -98.440 ;
        RECT -100.860 -98.870 -97.690 -98.465 ;
        RECT -95.030 -98.635 -94.855 -98.465 ;
        RECT -103.695 -100.735 -103.525 -99.195 ;
        RECT -103.205 -100.735 -103.035 -99.195 ;
        RECT -102.715 -100.735 -102.545 -99.195 ;
        RECT -102.225 -100.735 -102.055 -99.195 ;
        RECT -101.735 -100.735 -101.565 -99.195 ;
        RECT -103.210 -100.975 -103.035 -100.735 ;
        RECT -99.640 -100.905 -99.335 -98.870 ;
        RECT -97.995 -98.880 -97.690 -98.870 ;
        RECT -95.515 -100.175 -95.345 -98.635 ;
        RECT -95.025 -100.175 -94.855 -98.635 ;
        RECT -94.535 -100.175 -94.365 -98.635 ;
        RECT -94.045 -100.175 -93.875 -98.635 ;
        RECT -93.555 -100.175 -93.385 -98.635 ;
        RECT -95.675 -100.390 -95.320 -100.385 ;
        RECT -93.615 -100.390 -93.245 -100.360 ;
        RECT -95.675 -100.395 -93.245 -100.390 ;
        RECT -96.805 -100.585 -93.245 -100.395 ;
        RECT -91.460 -100.500 -91.155 -98.465 ;
        RECT -87.790 -98.745 -87.620 -97.275 ;
        RECT -87.300 -98.665 -87.130 -97.205 ;
        RECT -86.845 -97.280 -86.610 -96.685 ;
        RECT -88.335 -98.975 -87.560 -98.915 ;
        RECT -88.520 -99.145 -87.560 -98.975 ;
        RECT -88.335 -99.190 -87.560 -99.145 ;
        RECT -87.330 -99.015 -87.105 -98.665 ;
        RECT -86.810 -98.745 -86.640 -97.280 ;
        RECT -85.635 -97.330 -85.400 -96.685 ;
        RECT -85.600 -98.745 -85.430 -97.330 ;
        RECT -85.110 -98.700 -84.940 -97.205 ;
        RECT -76.290 -98.030 -76.050 -96.240 ;
        RECT -74.640 -96.325 -49.335 -96.130 ;
        RECT -46.185 -96.205 -45.990 -95.895 ;
        RECT -44.415 -96.205 -44.200 -94.985 ;
        RECT -43.315 -95.055 -43.145 -92.065 ;
        RECT -42.825 -94.955 -42.655 -92.015 ;
        RECT -42.355 -92.055 -42.145 -91.845 ;
        RECT -42.845 -95.225 -42.635 -94.955 ;
        RECT -42.335 -94.965 -42.165 -92.055 ;
        RECT -41.280 -94.935 -41.110 -92.015 ;
        RECT -37.225 -92.475 -33.585 -92.305 ;
        RECT -37.225 -94.035 -37.055 -92.475 ;
        RECT -36.735 -94.215 -36.565 -92.995 ;
        RECT -36.245 -94.035 -36.075 -92.475 ;
        RECT -35.645 -92.820 -33.935 -92.650 ;
        RECT -35.645 -94.035 -35.475 -92.820 ;
        RECT -35.155 -94.215 -34.985 -92.995 ;
        RECT -34.665 -94.035 -34.495 -92.820 ;
        RECT -37.780 -94.385 -34.410 -94.215 ;
        RECT -43.340 -95.420 -42.635 -95.225 ;
        RECT -42.360 -95.230 -42.150 -94.965 ;
        RECT -41.300 -95.230 -41.090 -94.935 ;
        RECT -42.360 -95.410 -41.090 -95.230 ;
        RECT -43.340 -95.480 -43.125 -95.420 ;
        RECT -44.030 -95.755 -43.125 -95.480 ;
        RECT -43.340 -96.105 -43.125 -95.755 ;
        RECT -42.690 -95.640 -41.915 -95.590 ;
        RECT -39.990 -95.640 -39.330 -95.285 ;
        RECT -42.690 -95.820 -39.330 -95.640 ;
        RECT -42.690 -95.865 -41.915 -95.820 ;
        RECT -72.610 -96.390 -71.950 -96.325 ;
        RECT -49.995 -96.380 -49.335 -96.325 ;
        RECT -46.205 -96.405 -43.530 -96.205 ;
        RECT -43.340 -96.305 -41.570 -96.105 ;
        RECT -46.205 -96.420 -43.770 -96.405 ;
        RECT -75.700 -96.900 -73.030 -96.560 ;
        RECT -71.045 -96.675 -67.880 -96.505 ;
        RECT -75.695 -97.615 -75.525 -97.155 ;
        RECT -75.725 -97.920 -75.495 -97.615 ;
        RECT -75.205 -97.695 -75.035 -96.900 ;
        RECT -74.715 -97.615 -74.545 -97.155 ;
        RECT -75.875 -98.030 -75.495 -97.920 ;
        RECT -76.290 -98.080 -75.495 -98.030 ;
        RECT -74.745 -98.080 -74.515 -97.615 ;
        RECT -74.225 -97.695 -74.055 -96.900 ;
        RECT -73.735 -97.615 -73.565 -97.155 ;
        RECT -73.765 -98.080 -73.535 -97.615 ;
        RECT -73.245 -97.695 -73.075 -96.900 ;
        RECT -71.505 -97.375 -71.335 -96.905 ;
        RECT -71.045 -96.965 -70.825 -96.675 ;
        RECT -71.525 -97.590 -71.320 -97.375 ;
        RECT -71.015 -97.445 -70.845 -96.965 ;
        RECT -70.525 -97.380 -70.355 -96.905 ;
        RECT -70.060 -97.020 -69.840 -96.675 ;
        RECT -71.530 -97.625 -71.320 -97.590 ;
        RECT -70.540 -97.625 -70.335 -97.380 ;
        RECT -70.035 -97.445 -69.865 -97.020 ;
        RECT -69.545 -97.380 -69.375 -96.905 ;
        RECT -69.080 -97.020 -68.860 -96.675 ;
        RECT -69.570 -97.625 -69.365 -97.380 ;
        RECT -69.055 -97.445 -68.885 -97.020 ;
        RECT -68.565 -97.420 -68.395 -96.905 ;
        RECT -68.100 -96.965 -67.880 -96.675 ;
        RECT -66.985 -96.900 -59.530 -96.560 ;
        RECT -57.545 -96.675 -54.380 -96.505 ;
        RECT -68.075 -97.315 -67.905 -96.965 ;
        RECT -68.580 -97.625 -68.375 -97.420 ;
        RECT -71.530 -97.795 -68.375 -97.625 ;
        RECT -76.290 -98.215 -73.535 -98.080 ;
        RECT -76.285 -98.225 -73.535 -98.215 ;
        RECT -75.875 -98.270 -73.535 -98.225 ;
        RECT -73.355 -97.940 -72.515 -97.865 ;
        RECT -71.530 -97.940 -70.655 -97.795 ;
        RECT -73.355 -98.205 -70.655 -97.940 ;
        RECT -68.110 -97.990 -67.875 -97.315 ;
        RECT -66.980 -97.615 -66.810 -97.155 ;
        RECT -67.010 -97.920 -66.780 -97.615 ;
        RECT -66.490 -97.695 -66.320 -96.900 ;
        RECT -66.000 -97.615 -65.830 -97.155 ;
        RECT -73.355 -98.235 -72.515 -98.205 ;
        RECT -75.725 -98.310 -73.535 -98.270 ;
        RECT -75.725 -98.635 -75.495 -98.310 ;
        RECT -74.745 -98.635 -74.515 -98.310 ;
        RECT -85.130 -98.900 -84.910 -98.700 ;
        RECT -85.130 -98.915 -79.430 -98.900 ;
        RECT -87.330 -99.215 -85.560 -99.015 ;
        RECT -85.370 -99.115 -79.430 -98.915 ;
        RECT -89.010 -99.500 -88.660 -99.490 ;
        RECT -86.985 -99.500 -86.210 -99.455 ;
        RECT -89.010 -99.680 -86.210 -99.500 ;
        RECT -96.805 -100.595 -95.670 -100.585 ;
        RECT -93.615 -100.715 -93.245 -100.585 ;
        RECT -95.940 -100.875 -95.265 -100.835 ;
        RECT -96.040 -100.885 -95.265 -100.875 ;
        RECT -101.585 -100.975 -99.335 -100.905 ;
        RECT -108.965 -101.420 -99.185 -100.975 ;
        RECT -97.995 -101.065 -95.265 -100.885 ;
        RECT -92.680 -100.930 -89.605 -100.500 ;
        RECT -113.690 -101.735 -99.185 -101.420 ;
        RECT -113.690 -101.745 -107.320 -101.735 ;
        RECT -120.160 -103.645 -119.655 -102.780 ;
        RECT -97.610 -103.645 -97.325 -101.065 ;
        RECT -96.040 -101.075 -95.265 -101.065 ;
        RECT -95.940 -101.105 -95.265 -101.075 ;
        RECT -95.025 -100.990 -92.930 -100.950 ;
        RECT -95.025 -101.140 -92.875 -100.990 ;
        RECT -95.025 -102.860 -94.855 -101.140 ;
        RECT -94.045 -102.860 -93.875 -101.140 ;
        RECT -93.180 -101.885 -92.875 -101.140 ;
        RECT -91.980 -101.710 -91.810 -100.930 ;
        RECT -91.490 -101.710 -91.320 -101.170 ;
        RECT -91.000 -101.710 -90.830 -100.930 ;
        RECT -90.510 -101.710 -90.340 -101.170 ;
        RECT -89.010 -101.655 -88.660 -99.680 ;
        RECT -86.985 -99.730 -86.210 -99.680 ;
        RECT -85.775 -99.565 -85.560 -99.215 ;
        RECT -85.775 -99.840 -84.870 -99.565 ;
        RECT -85.775 -99.900 -85.560 -99.840 ;
        RECT -87.810 -100.090 -86.540 -99.910 ;
        RECT -87.810 -100.385 -87.600 -100.090 ;
        RECT -86.750 -100.355 -86.540 -100.090 ;
        RECT -86.265 -100.095 -85.560 -99.900 ;
        RECT -92.570 -101.885 -92.205 -101.855 ;
        RECT -93.180 -101.950 -92.205 -101.885 ;
        RECT -93.070 -102.090 -92.205 -101.950 ;
        RECT -92.570 -102.155 -92.205 -102.090 ;
        RECT -90.020 -102.005 -88.630 -101.655 ;
        RECT -91.980 -102.865 -91.810 -102.325 ;
        RECT -91.000 -102.865 -90.830 -102.325 ;
        RECT -90.020 -102.865 -89.850 -102.005 ;
        RECT -87.790 -103.305 -87.620 -100.385 ;
        RECT -86.735 -103.265 -86.565 -100.355 ;
        RECT -86.265 -100.365 -86.055 -100.095 ;
        RECT -86.755 -103.475 -86.545 -103.265 ;
        RECT -86.245 -103.305 -86.075 -100.365 ;
        RECT -85.755 -103.255 -85.585 -100.265 ;
        RECT -84.700 -100.335 -84.485 -99.115 ;
        RECT -83.570 -99.990 -83.045 -99.630 ;
        RECT -85.765 -103.475 -85.555 -103.255 ;
        RECT -84.695 -103.305 -84.525 -100.335 ;
        RECT -86.755 -103.645 -85.555 -103.475 ;
        RECT -120.160 -103.960 -97.325 -103.645 ;
        RECT -120.160 -103.995 -119.655 -103.960 ;
        RECT -112.915 -107.775 -112.745 -106.055 ;
        RECT -111.935 -107.775 -111.765 -106.055 ;
        RECT -109.870 -106.590 -109.700 -106.050 ;
        RECT -108.890 -106.590 -108.720 -106.050 ;
        RECT -110.460 -106.825 -110.095 -106.760 ;
        RECT -110.960 -106.965 -110.095 -106.825 ;
        RECT -111.070 -107.030 -110.095 -106.965 ;
        RECT -111.070 -107.775 -110.765 -107.030 ;
        RECT -110.460 -107.060 -110.095 -107.030 ;
        RECT -107.910 -106.910 -107.740 -106.050 ;
        RECT -104.050 -106.800 -103.880 -105.580 ;
        RECT -103.070 -106.800 -102.900 -105.580 ;
        RECT -102.090 -106.800 -101.920 -105.580 ;
        RECT -104.925 -106.855 -104.250 -106.815 ;
        RECT -106.725 -106.910 -104.250 -106.855 ;
        RECT -107.910 -107.030 -104.250 -106.910 ;
        RECT -104.050 -106.985 -101.275 -106.800 ;
        RECT -112.915 -107.925 -110.765 -107.775 ;
        RECT -112.915 -107.965 -110.820 -107.925 ;
        RECT -109.870 -107.985 -109.700 -107.205 ;
        RECT -109.380 -107.745 -109.210 -107.205 ;
        RECT -108.890 -107.985 -108.720 -107.205 ;
        RECT -108.400 -107.745 -108.230 -107.205 ;
        RECT -107.910 -107.260 -106.520 -107.030 ;
        RECT -105.020 -107.040 -104.250 -107.030 ;
        RECT -104.925 -107.085 -104.250 -107.040 ;
        RECT -105.500 -107.270 -105.210 -107.230 ;
        RECT -103.245 -107.270 -102.570 -107.225 ;
        RECT -105.630 -107.460 -102.570 -107.270 ;
        RECT -110.570 -108.415 -107.495 -107.985 ;
        RECT -113.405 -110.280 -113.235 -108.740 ;
        RECT -112.915 -110.280 -112.745 -108.740 ;
        RECT -112.425 -110.280 -112.255 -108.740 ;
        RECT -111.935 -110.280 -111.765 -108.740 ;
        RECT -111.445 -110.280 -111.275 -108.740 ;
        RECT -112.920 -110.540 -112.745 -110.280 ;
        RECT -109.350 -110.450 -109.045 -108.415 ;
        RECT -107.055 -109.055 -106.765 -108.370 ;
        RECT -105.985 -108.385 -105.695 -107.885 ;
        RECT -105.500 -107.915 -105.210 -107.460 ;
        RECT -103.245 -107.495 -102.570 -107.460 ;
        RECT -102.305 -107.680 -101.630 -107.615 ;
        RECT -105.010 -107.850 -101.630 -107.680 ;
        RECT -105.010 -108.385 -104.840 -107.850 ;
        RECT -102.305 -107.885 -101.630 -107.850 ;
        RECT -101.460 -107.675 -101.275 -106.985 ;
        RECT -99.250 -107.675 -98.575 -107.625 ;
        RECT -101.460 -107.860 -98.575 -107.675 ;
        RECT -101.460 -108.130 -101.275 -107.860 ;
        RECT -99.250 -107.895 -98.575 -107.860 ;
        RECT -98.400 -107.985 -98.230 -105.580 ;
        RECT -94.895 -107.505 -94.725 -106.465 ;
        RECT -93.915 -107.505 -93.745 -106.465 ;
        RECT -92.935 -107.505 -92.765 -106.465 ;
        RECT -90.030 -107.540 -89.860 -105.820 ;
        RECT -89.050 -107.540 -88.880 -105.820 ;
        RECT -86.985 -106.355 -86.815 -105.815 ;
        RECT -86.005 -106.355 -85.835 -105.815 ;
        RECT -87.575 -106.590 -87.210 -106.525 ;
        RECT -88.075 -106.730 -87.210 -106.590 ;
        RECT -88.185 -106.795 -87.210 -106.730 ;
        RECT -88.185 -107.540 -87.880 -106.795 ;
        RECT -87.575 -106.825 -87.210 -106.795 ;
        RECT -85.025 -106.675 -84.855 -105.815 ;
        RECT -83.515 -106.675 -83.165 -99.990 ;
        RECT -90.945 -107.605 -90.270 -107.575 ;
        RECT -91.045 -107.615 -90.270 -107.605 ;
        RECT -96.355 -107.740 -95.705 -107.655 ;
        RECT -95.485 -107.740 -95.120 -107.675 ;
        RECT -96.355 -107.945 -95.120 -107.740 ;
        RECT -92.080 -107.795 -90.270 -107.615 ;
        RECT -90.030 -107.690 -87.880 -107.540 ;
        RECT -90.030 -107.730 -87.935 -107.690 ;
        RECT -86.985 -107.750 -86.815 -106.970 ;
        RECT -86.495 -107.510 -86.325 -106.970 ;
        RECT -86.005 -107.750 -85.835 -106.970 ;
        RECT -85.515 -107.510 -85.345 -106.970 ;
        RECT -85.025 -107.025 -83.165 -106.675 ;
        RECT -91.045 -107.805 -90.270 -107.795 ;
        RECT -90.945 -107.845 -90.270 -107.805 ;
        RECT -96.355 -107.985 -95.705 -107.945 ;
        RECT -95.485 -107.975 -95.120 -107.945 ;
        RECT -105.985 -108.555 -104.840 -108.385 ;
        RECT -104.540 -108.300 -102.325 -108.130 ;
        RECT -101.460 -108.300 -100.295 -108.130 ;
        RECT -105.985 -108.570 -105.695 -108.555 ;
        RECT -104.540 -110.155 -104.370 -108.300 ;
        RECT -103.560 -108.305 -102.325 -108.300 ;
        RECT -111.295 -110.540 -105.450 -110.450 ;
        RECT -113.505 -110.845 -105.450 -110.540 ;
        RECT -111.300 -111.025 -105.450 -110.845 ;
        RECT -106.025 -111.115 -105.450 -111.025 ;
        RECT -104.050 -111.100 -103.880 -108.615 ;
        RECT -103.560 -110.155 -103.390 -108.305 ;
        RECT -102.500 -108.620 -102.325 -108.305 ;
        RECT -102.990 -110.115 -102.820 -108.620 ;
        RECT -102.990 -110.635 -102.815 -110.115 ;
        RECT -102.500 -110.160 -102.330 -108.620 ;
        RECT -102.010 -110.105 -101.840 -108.620 ;
        RECT -102.010 -110.635 -101.835 -110.105 ;
        RECT -101.445 -110.160 -101.275 -108.300 ;
        RECT -102.990 -110.650 -101.835 -110.635 ;
        RECT -100.955 -110.650 -100.785 -108.620 ;
        RECT -100.465 -110.160 -100.295 -108.300 ;
        RECT -98.400 -108.155 -95.705 -107.985 ;
        RECT -93.420 -108.095 -90.675 -108.085 ;
        RECT -88.620 -108.095 -88.250 -107.965 ;
        RECT -93.420 -108.115 -88.250 -108.095 ;
        RECT -102.990 -110.820 -100.785 -110.650 ;
        RECT -98.890 -110.965 -98.720 -109.120 ;
        RECT -98.400 -110.160 -98.230 -108.155 ;
        RECT -96.355 -108.405 -95.705 -108.155 ;
        RECT -94.895 -109.395 -94.725 -108.115 ;
        RECT -94.405 -109.155 -94.235 -108.115 ;
        RECT -93.915 -109.395 -93.745 -108.115 ;
        RECT -93.425 -108.285 -88.250 -108.115 ;
        RECT -87.685 -108.180 -83.760 -107.750 ;
        RECT -93.425 -109.155 -93.255 -108.285 ;
        RECT -90.680 -108.290 -88.250 -108.285 ;
        RECT -90.680 -108.295 -90.325 -108.290 ;
        RECT -88.620 -108.320 -88.250 -108.290 ;
        RECT -95.595 -109.825 -90.905 -109.395 ;
        RECT -91.335 -110.230 -90.905 -109.825 ;
        RECT -90.520 -110.045 -90.350 -108.505 ;
        RECT -90.030 -110.045 -89.860 -108.505 ;
        RECT -89.540 -110.045 -89.370 -108.505 ;
        RECT -89.050 -110.045 -88.880 -108.505 ;
        RECT -88.560 -110.045 -88.390 -108.505 ;
        RECT -90.035 -110.230 -89.860 -110.045 ;
        RECT -86.465 -110.215 -86.160 -108.180 ;
        RECT -88.410 -110.230 -86.160 -110.215 ;
        RECT -91.335 -110.520 -86.160 -110.230 ;
        RECT -91.335 -110.660 -88.010 -110.520 ;
        RECT -91.155 -110.965 -90.105 -110.660 ;
        RECT -99.895 -111.100 -90.105 -110.965 ;
        RECT -104.540 -111.115 -90.105 -111.100 ;
        RECT -106.025 -111.740 -90.105 -111.115 ;
        RECT -85.495 -110.910 -84.155 -110.660 ;
        RECT -80.345 -110.910 -79.430 -99.115 ;
        RECT -75.695 -99.595 -75.525 -98.635 ;
        RECT -74.715 -99.595 -74.545 -98.635 ;
        RECT -73.765 -99.575 -73.535 -98.310 ;
        RECT -71.530 -98.630 -70.655 -98.205 ;
        RECT -68.735 -98.360 -67.875 -97.990 ;
        RECT -71.530 -98.800 -68.390 -98.630 ;
        RECT -71.530 -99.020 -71.320 -98.800 ;
        RECT -71.505 -99.520 -71.335 -99.020 ;
        RECT -71.015 -99.435 -70.845 -98.980 ;
        RECT -70.530 -99.070 -70.350 -98.800 ;
        RECT -69.560 -98.980 -69.380 -98.800 ;
        RECT -73.735 -99.595 -73.565 -99.575 ;
        RECT -71.040 -99.690 -70.830 -99.435 ;
        RECT -70.525 -99.520 -70.355 -99.070 ;
        RECT -70.035 -99.410 -69.865 -98.980 ;
        RECT -69.560 -99.070 -69.375 -98.980 ;
        RECT -70.060 -99.690 -69.850 -99.410 ;
        RECT -69.545 -99.520 -69.375 -99.070 ;
        RECT -69.055 -99.415 -68.885 -98.980 ;
        RECT -68.570 -99.060 -68.390 -98.800 ;
        RECT -69.090 -99.690 -68.880 -99.415 ;
        RECT -68.565 -99.520 -68.395 -99.060 ;
        RECT -68.110 -99.095 -67.875 -98.360 ;
        RECT -67.650 -98.080 -66.780 -97.920 ;
        RECT -66.030 -98.080 -65.800 -97.615 ;
        RECT -65.510 -97.695 -65.340 -96.900 ;
        RECT -65.020 -97.615 -64.850 -97.155 ;
        RECT -65.050 -98.080 -64.820 -97.615 ;
        RECT -64.530 -97.695 -64.360 -96.900 ;
        RECT -67.650 -98.270 -64.820 -98.080 ;
        RECT -64.640 -97.890 -63.800 -97.865 ;
        RECT -63.500 -97.890 -63.200 -97.525 ;
        RECT -64.640 -98.180 -63.200 -97.890 ;
        RECT -62.925 -97.975 -62.625 -97.400 ;
        RECT -62.195 -97.615 -62.025 -97.155 ;
        RECT -62.225 -97.920 -61.995 -97.615 ;
        RECT -61.705 -97.695 -61.535 -96.900 ;
        RECT -61.215 -97.615 -61.045 -97.155 ;
        RECT -62.375 -97.975 -61.995 -97.920 ;
        RECT -64.640 -98.235 -63.800 -98.180 ;
        RECT -63.500 -98.185 -63.200 -98.180 ;
        RECT -62.950 -98.080 -61.995 -97.975 ;
        RECT -61.245 -98.080 -61.015 -97.615 ;
        RECT -60.725 -97.695 -60.555 -96.900 ;
        RECT -60.235 -97.615 -60.065 -97.155 ;
        RECT -60.265 -98.080 -60.035 -97.615 ;
        RECT -59.745 -97.695 -59.575 -96.900 ;
        RECT -58.020 -97.375 -57.790 -96.765 ;
        RECT -57.545 -96.965 -57.325 -96.675 ;
        RECT -58.025 -97.425 -57.790 -97.375 ;
        RECT -58.025 -97.590 -57.820 -97.425 ;
        RECT -57.515 -97.445 -57.345 -96.965 ;
        RECT -57.025 -97.380 -56.855 -96.905 ;
        RECT -56.560 -97.020 -56.340 -96.675 ;
        RECT -58.030 -97.625 -57.820 -97.590 ;
        RECT -57.040 -97.625 -56.835 -97.380 ;
        RECT -56.535 -97.445 -56.365 -97.020 ;
        RECT -56.045 -97.380 -55.875 -96.905 ;
        RECT -55.580 -97.020 -55.360 -96.675 ;
        RECT -56.070 -97.625 -55.865 -97.380 ;
        RECT -55.555 -97.445 -55.385 -97.020 ;
        RECT -55.065 -97.420 -54.895 -96.905 ;
        RECT -54.600 -96.965 -54.380 -96.675 ;
        RECT -53.485 -96.900 -46.405 -96.560 ;
        RECT -54.575 -97.315 -54.405 -96.965 ;
        RECT -55.080 -97.625 -54.875 -97.420 ;
        RECT -58.030 -97.795 -54.875 -97.625 ;
        RECT -62.950 -98.200 -60.035 -98.080 ;
        RECT -67.650 -98.390 -67.285 -98.270 ;
        RECT -68.075 -99.465 -67.905 -99.095 ;
        RECT -67.655 -99.230 -67.285 -98.390 ;
        RECT -67.010 -98.310 -64.820 -98.270 ;
        RECT -67.010 -98.635 -66.780 -98.310 ;
        RECT -66.030 -98.635 -65.800 -98.310 ;
        RECT -68.080 -99.690 -67.900 -99.465 ;
        RECT -66.980 -99.595 -66.810 -98.635 ;
        RECT -66.000 -99.595 -65.830 -98.635 ;
        RECT -65.050 -99.575 -64.820 -98.310 ;
        RECT -64.030 -98.870 -63.745 -98.665 ;
        RECT -62.950 -98.870 -62.725 -98.200 ;
        RECT -62.375 -98.270 -60.035 -98.200 ;
        RECT -59.855 -97.905 -59.015 -97.865 ;
        RECT -58.030 -97.905 -57.155 -97.795 ;
        RECT -59.855 -98.190 -57.155 -97.905 ;
        RECT -54.610 -97.990 -54.375 -97.315 ;
        RECT -53.480 -97.615 -53.310 -97.155 ;
        RECT -53.510 -97.920 -53.280 -97.615 ;
        RECT -52.990 -97.695 -52.820 -96.900 ;
        RECT -52.500 -97.615 -52.330 -97.155 ;
        RECT -59.855 -98.235 -59.015 -98.190 ;
        RECT -62.225 -98.310 -60.035 -98.270 ;
        RECT -62.225 -98.635 -61.995 -98.310 ;
        RECT -61.245 -98.635 -61.015 -98.310 ;
        RECT -64.030 -99.095 -62.725 -98.870 ;
        RECT -64.030 -99.485 -63.745 -99.095 ;
        RECT -65.020 -99.595 -64.850 -99.575 ;
        RECT -62.195 -99.595 -62.025 -98.635 ;
        RECT -61.215 -99.595 -61.045 -98.635 ;
        RECT -60.265 -99.575 -60.035 -98.310 ;
        RECT -58.030 -98.630 -57.155 -98.190 ;
        RECT -55.235 -98.360 -54.375 -97.990 ;
        RECT -58.030 -98.800 -54.890 -98.630 ;
        RECT -58.030 -99.020 -57.820 -98.800 ;
        RECT -58.005 -99.520 -57.835 -99.020 ;
        RECT -57.515 -99.435 -57.345 -98.980 ;
        RECT -57.030 -99.070 -56.850 -98.800 ;
        RECT -56.060 -98.980 -55.880 -98.800 ;
        RECT -60.235 -99.595 -60.065 -99.575 ;
        RECT -71.040 -99.860 -67.900 -99.690 ;
        RECT -57.540 -99.690 -57.330 -99.435 ;
        RECT -57.025 -99.520 -56.855 -99.070 ;
        RECT -56.535 -99.410 -56.365 -98.980 ;
        RECT -56.060 -99.070 -55.875 -98.980 ;
        RECT -56.560 -99.690 -56.350 -99.410 ;
        RECT -56.045 -99.520 -55.875 -99.070 ;
        RECT -55.555 -99.415 -55.385 -98.980 ;
        RECT -55.070 -99.060 -54.890 -98.800 ;
        RECT -55.590 -99.690 -55.380 -99.415 ;
        RECT -55.065 -99.520 -54.895 -99.060 ;
        RECT -54.610 -99.095 -54.375 -98.360 ;
        RECT -54.150 -98.080 -53.280 -97.920 ;
        RECT -52.530 -98.080 -52.300 -97.615 ;
        RECT -52.010 -97.695 -51.840 -96.900 ;
        RECT -51.520 -97.615 -51.350 -97.155 ;
        RECT -51.550 -98.080 -51.320 -97.615 ;
        RECT -51.030 -97.695 -50.860 -96.900 ;
        RECT -54.150 -98.270 -51.320 -98.080 ;
        RECT -51.140 -97.890 -50.300 -97.865 ;
        RECT -51.140 -97.950 -50.125 -97.890 ;
        RECT -49.840 -97.950 -49.540 -97.520 ;
        RECT -49.070 -97.615 -48.900 -97.155 ;
        RECT -49.100 -97.920 -48.870 -97.615 ;
        RECT -48.580 -97.695 -48.410 -96.900 ;
        RECT -48.090 -97.615 -47.920 -97.155 ;
        RECT -49.250 -97.950 -48.870 -97.920 ;
        RECT -51.140 -98.080 -48.870 -97.950 ;
        RECT -48.120 -98.080 -47.890 -97.615 ;
        RECT -47.600 -97.695 -47.430 -96.900 ;
        RECT -47.110 -97.615 -46.940 -97.155 ;
        RECT -47.140 -98.080 -46.910 -97.615 ;
        RECT -46.620 -97.695 -46.450 -96.900 ;
        RECT -46.185 -97.865 -45.990 -96.420 ;
        RECT -43.990 -96.620 -43.770 -96.420 ;
        RECT -51.140 -98.160 -46.910 -98.080 ;
        RECT -51.140 -98.180 -50.125 -98.160 ;
        RECT -49.840 -98.180 -49.540 -98.160 ;
        RECT -51.140 -98.235 -50.300 -98.180 ;
        RECT -49.250 -98.270 -46.910 -98.160 ;
        RECT -46.730 -98.235 -45.890 -97.865 ;
        RECT -43.960 -98.115 -43.790 -96.620 ;
        RECT -43.470 -97.990 -43.300 -96.575 ;
        RECT -54.150 -98.390 -53.785 -98.270 ;
        RECT -54.575 -99.465 -54.405 -99.095 ;
        RECT -54.155 -99.230 -53.785 -98.390 ;
        RECT -53.510 -98.310 -51.320 -98.270 ;
        RECT -53.510 -98.635 -53.280 -98.310 ;
        RECT -52.530 -98.635 -52.300 -98.310 ;
        RECT -54.580 -99.690 -54.400 -99.465 ;
        RECT -53.480 -99.595 -53.310 -98.635 ;
        RECT -52.500 -99.595 -52.330 -98.635 ;
        RECT -51.550 -99.575 -51.320 -98.310 ;
        RECT -49.100 -98.310 -46.910 -98.270 ;
        RECT -49.100 -98.635 -48.870 -98.310 ;
        RECT -48.120 -98.635 -47.890 -98.310 ;
        RECT -50.530 -99.485 -50.245 -98.665 ;
        RECT -51.520 -99.595 -51.350 -99.575 ;
        RECT -49.070 -99.595 -48.900 -98.635 ;
        RECT -48.090 -99.595 -47.920 -98.635 ;
        RECT -47.140 -99.575 -46.910 -98.310 ;
        RECT -45.620 -98.640 -44.230 -98.635 ;
        RECT -43.500 -98.640 -43.265 -97.990 ;
        RECT -42.260 -98.040 -42.090 -96.575 ;
        RECT -41.795 -96.655 -41.570 -96.305 ;
        RECT -41.340 -96.175 -40.565 -96.130 ;
        RECT -41.340 -96.345 -38.530 -96.175 ;
        RECT -41.340 -96.405 -40.565 -96.345 ;
        RECT -42.290 -98.640 -42.055 -98.040 ;
        RECT -41.770 -98.115 -41.600 -96.655 ;
        RECT -41.280 -98.045 -41.110 -96.575 ;
        RECT -41.310 -98.640 -41.075 -98.045 ;
        RECT -45.620 -99.050 -40.665 -98.640 ;
        RECT -47.110 -99.595 -46.940 -99.575 ;
        RECT -57.540 -99.860 -54.400 -99.690 ;
        RECT -66.515 -101.565 -59.130 -101.000 ;
        RECT -70.670 -103.040 -68.425 -102.950 ;
        RECT -66.515 -103.040 -66.210 -101.565 ;
        RECT -62.880 -102.155 -62.645 -101.565 ;
        RECT -70.670 -103.255 -66.210 -103.040 ;
        RECT -70.085 -103.515 -69.910 -103.255 ;
        RECT -68.460 -103.345 -66.210 -103.255 ;
        RECT -70.570 -105.055 -70.400 -103.515 ;
        RECT -70.080 -105.055 -69.910 -103.515 ;
        RECT -69.590 -105.055 -69.420 -103.515 ;
        RECT -69.100 -105.055 -68.930 -103.515 ;
        RECT -68.610 -105.055 -68.440 -103.515 ;
        RECT -66.515 -105.380 -66.210 -103.345 ;
        RECT -62.845 -103.625 -62.675 -102.155 ;
        RECT -62.355 -103.545 -62.185 -102.085 ;
        RECT -61.900 -102.160 -61.665 -101.565 ;
        RECT -63.390 -103.855 -62.615 -103.795 ;
        RECT -63.575 -104.025 -62.615 -103.855 ;
        RECT -63.390 -104.070 -62.615 -104.025 ;
        RECT -62.385 -103.895 -62.160 -103.545 ;
        RECT -61.865 -103.625 -61.695 -102.160 ;
        RECT -60.690 -102.210 -60.455 -101.565 ;
        RECT -60.655 -103.625 -60.485 -102.210 ;
        RECT -60.165 -103.580 -59.995 -102.085 ;
        RECT -60.185 -103.780 -59.965 -103.580 ;
        RECT -60.185 -103.795 -44.785 -103.780 ;
        RECT -62.385 -104.095 -60.615 -103.895 ;
        RECT -60.425 -103.995 -44.785 -103.795 ;
        RECT -64.065 -104.380 -63.715 -104.370 ;
        RECT -62.040 -104.380 -61.265 -104.335 ;
        RECT -64.065 -104.560 -61.265 -104.380 ;
        RECT -73.295 -105.765 -72.365 -105.480 ;
        RECT -70.995 -105.755 -70.320 -105.715 ;
        RECT -71.095 -105.765 -70.320 -105.755 ;
        RECT -73.295 -105.945 -70.320 -105.765 ;
        RECT -67.735 -105.810 -64.660 -105.380 ;
        RECT -73.295 -106.250 -72.365 -105.945 ;
        RECT -71.095 -105.955 -70.320 -105.945 ;
        RECT -70.995 -105.985 -70.320 -105.955 ;
        RECT -70.080 -105.870 -67.985 -105.830 ;
        RECT -70.080 -106.020 -67.930 -105.870 ;
        RECT -70.080 -107.740 -69.910 -106.020 ;
        RECT -69.100 -107.740 -68.930 -106.020 ;
        RECT -68.235 -106.765 -67.930 -106.020 ;
        RECT -67.035 -106.590 -66.865 -105.810 ;
        RECT -66.545 -106.590 -66.375 -106.050 ;
        RECT -66.055 -106.590 -65.885 -105.810 ;
        RECT -65.565 -106.590 -65.395 -106.050 ;
        RECT -64.065 -106.535 -63.715 -104.560 ;
        RECT -62.040 -104.610 -61.265 -104.560 ;
        RECT -60.830 -104.445 -60.615 -104.095 ;
        RECT -60.830 -104.720 -59.925 -104.445 ;
        RECT -60.830 -104.780 -60.615 -104.720 ;
        RECT -62.865 -104.970 -61.595 -104.790 ;
        RECT -62.865 -105.265 -62.655 -104.970 ;
        RECT -61.805 -105.235 -61.595 -104.970 ;
        RECT -61.320 -104.975 -60.615 -104.780 ;
        RECT -67.625 -106.765 -67.260 -106.735 ;
        RECT -68.235 -106.830 -67.260 -106.765 ;
        RECT -68.125 -106.970 -67.260 -106.830 ;
        RECT -67.625 -107.035 -67.260 -106.970 ;
        RECT -65.075 -106.885 -63.685 -106.535 ;
        RECT -67.035 -107.745 -66.865 -107.205 ;
        RECT -66.055 -107.745 -65.885 -107.205 ;
        RECT -65.075 -107.745 -64.905 -106.885 ;
        RECT -62.845 -108.185 -62.675 -105.265 ;
        RECT -61.790 -108.145 -61.620 -105.235 ;
        RECT -61.320 -105.245 -61.110 -104.975 ;
        RECT -61.810 -108.355 -61.600 -108.145 ;
        RECT -61.300 -108.185 -61.130 -105.245 ;
        RECT -60.810 -108.135 -60.640 -105.145 ;
        RECT -59.755 -105.215 -59.540 -103.995 ;
        RECT -45.665 -104.390 -44.785 -103.995 ;
        RECT -58.625 -104.870 -58.100 -104.510 ;
        RECT -60.820 -108.355 -60.610 -108.135 ;
        RECT -59.750 -108.185 -59.580 -105.215 ;
        RECT -61.810 -108.525 -60.610 -108.355 ;
        RECT -85.495 -111.825 -79.430 -110.910 ;
        RECT -85.495 -111.985 -84.155 -111.825 ;
        RECT -69.950 -112.385 -69.780 -111.345 ;
        RECT -68.970 -112.385 -68.800 -111.345 ;
        RECT -67.990 -112.385 -67.820 -111.345 ;
        RECT -65.085 -112.420 -64.915 -110.700 ;
        RECT -64.105 -112.420 -63.935 -110.700 ;
        RECT -62.040 -111.235 -61.870 -110.695 ;
        RECT -61.060 -111.235 -60.890 -110.695 ;
        RECT -62.630 -111.470 -62.265 -111.405 ;
        RECT -63.130 -111.610 -62.265 -111.470 ;
        RECT -63.240 -111.675 -62.265 -111.610 ;
        RECT -63.240 -112.420 -62.935 -111.675 ;
        RECT -62.630 -111.705 -62.265 -111.675 ;
        RECT -60.080 -111.555 -59.910 -110.695 ;
        RECT -58.570 -111.555 -58.220 -104.870 ;
        RECT -38.700 -107.640 -38.530 -96.345 ;
        RECT -37.780 -102.085 -37.610 -94.385 ;
        RECT -37.230 -95.055 -36.535 -94.785 ;
        RECT -34.580 -94.960 -34.410 -94.385 ;
        RECT -34.105 -94.580 -33.935 -92.820 ;
        RECT -33.755 -94.210 -33.585 -92.475 ;
        RECT -24.725 -92.475 -21.085 -92.305 ;
        RECT -32.855 -94.210 -32.685 -92.995 ;
        RECT -33.755 -94.380 -32.685 -94.210 ;
        RECT -31.875 -94.580 -31.705 -92.995 ;
        RECT -30.325 -93.960 -30.155 -92.995 ;
        RECT -28.780 -93.950 -28.610 -92.995 ;
        RECT -34.105 -94.750 -31.705 -94.580 ;
        RECT -31.440 -94.835 -30.745 -94.565 ;
        RECT -34.580 -95.130 -33.850 -94.960 ;
        RECT -37.235 -95.645 -35.580 -95.460 ;
        RECT -35.320 -95.575 -34.625 -95.305 ;
        RECT -34.020 -95.440 -33.850 -95.130 ;
        RECT -33.485 -95.205 -32.790 -94.935 ;
        RECT -34.020 -95.610 -31.215 -95.440 ;
        RECT -37.235 -96.060 -37.050 -95.645 ;
        RECT -35.765 -95.765 -35.580 -95.645 ;
        RECT -35.765 -95.950 -34.985 -95.765 ;
        RECT -37.225 -97.005 -37.055 -96.060 ;
        RECT -37.245 -97.620 -37.050 -97.005 ;
        RECT -36.735 -97.250 -36.565 -96.025 ;
        RECT -35.170 -96.055 -34.985 -95.950 ;
        RECT -35.155 -97.065 -34.985 -96.055 ;
        RECT -34.675 -96.070 -33.175 -95.875 ;
        RECT -34.665 -97.065 -34.495 -96.070 ;
        RECT -33.345 -97.065 -33.175 -96.070 ;
        RECT -32.855 -97.065 -32.685 -95.610 ;
        RECT -31.875 -96.980 -31.705 -96.025 ;
        RECT -31.875 -97.250 -31.695 -96.980 ;
        RECT -31.385 -97.065 -31.215 -95.610 ;
        RECT -30.350 -95.655 -30.135 -93.960 ;
        RECT -28.800 -94.935 -28.585 -93.950 ;
        RECT -24.725 -94.035 -24.555 -92.475 ;
        RECT -24.235 -94.215 -24.065 -92.995 ;
        RECT -23.745 -94.035 -23.575 -92.475 ;
        RECT -23.145 -92.820 -21.435 -92.650 ;
        RECT -23.145 -94.035 -22.975 -92.820 ;
        RECT -22.655 -94.215 -22.485 -92.995 ;
        RECT -22.165 -94.035 -21.995 -92.820 ;
        RECT -25.565 -94.385 -21.910 -94.215 ;
        RECT -28.365 -94.865 -27.670 -94.595 ;
        RECT -29.300 -95.165 -28.585 -94.935 ;
        RECT -29.930 -95.605 -29.235 -95.335 ;
        RECT -30.830 -95.885 -30.135 -95.655 ;
        RECT -30.350 -96.110 -30.135 -95.885 ;
        RECT -30.325 -97.065 -30.155 -96.110 ;
        RECT -29.835 -97.030 -29.665 -96.025 ;
        RECT -28.800 -96.120 -28.585 -95.165 ;
        RECT -36.735 -97.430 -31.695 -97.250 ;
        RECT -29.860 -97.450 -29.645 -97.030 ;
        RECT -28.780 -97.065 -28.610 -96.120 ;
        RECT -28.290 -97.020 -28.120 -96.025 ;
        RECT -25.565 -96.200 -25.395 -94.385 ;
        RECT -24.730 -95.055 -24.035 -94.785 ;
        RECT -22.080 -94.960 -21.910 -94.385 ;
        RECT -21.605 -94.580 -21.435 -92.820 ;
        RECT -21.255 -94.210 -21.085 -92.475 ;
        RECT -12.225 -92.475 -8.585 -92.305 ;
        RECT -20.355 -94.210 -20.185 -92.995 ;
        RECT -21.255 -94.380 -20.185 -94.210 ;
        RECT -19.375 -94.580 -19.205 -92.995 ;
        RECT -17.825 -93.960 -17.655 -92.995 ;
        RECT -16.280 -93.950 -16.110 -92.995 ;
        RECT -21.605 -94.750 -19.205 -94.580 ;
        RECT -18.940 -94.835 -18.245 -94.565 ;
        RECT -22.080 -95.130 -21.350 -94.960 ;
        RECT -21.520 -95.440 -21.350 -95.130 ;
        RECT -20.985 -95.205 -20.290 -94.935 ;
        RECT -24.735 -95.645 -23.080 -95.460 ;
        RECT -21.520 -95.610 -18.715 -95.440 ;
        RECT -24.735 -96.060 -24.550 -95.645 ;
        RECT -23.265 -95.765 -23.080 -95.645 ;
        RECT -23.265 -95.950 -22.485 -95.765 ;
        RECT -25.595 -96.880 -25.365 -96.200 ;
        RECT -24.725 -97.005 -24.555 -96.060 ;
        RECT -28.315 -97.445 -28.100 -97.020 ;
        RECT -24.745 -97.445 -24.550 -97.005 ;
        RECT -24.235 -97.250 -24.065 -96.025 ;
        RECT -22.670 -96.055 -22.485 -95.950 ;
        RECT -22.655 -97.065 -22.485 -96.055 ;
        RECT -22.175 -96.070 -20.675 -95.875 ;
        RECT -22.165 -97.065 -21.995 -96.070 ;
        RECT -20.845 -97.065 -20.675 -96.070 ;
        RECT -20.355 -97.065 -20.185 -95.610 ;
        RECT -19.375 -96.980 -19.205 -96.025 ;
        RECT -19.375 -97.250 -19.195 -96.980 ;
        RECT -18.885 -97.065 -18.715 -95.610 ;
        RECT -17.850 -95.655 -17.635 -93.960 ;
        RECT -16.300 -94.935 -16.085 -93.950 ;
        RECT -12.225 -94.035 -12.055 -92.475 ;
        RECT -11.735 -94.215 -11.565 -92.995 ;
        RECT -11.245 -94.035 -11.075 -92.475 ;
        RECT -10.645 -92.820 -8.935 -92.650 ;
        RECT -10.645 -94.035 -10.475 -92.820 ;
        RECT -10.155 -94.215 -9.985 -92.995 ;
        RECT -9.665 -94.035 -9.495 -92.820 ;
        RECT -12.825 -94.385 -9.410 -94.215 ;
        RECT -15.865 -94.865 -15.170 -94.595 ;
        RECT -16.800 -95.165 -16.085 -94.935 ;
        RECT -18.330 -95.885 -17.635 -95.655 ;
        RECT -17.850 -96.110 -17.635 -95.885 ;
        RECT -17.825 -97.065 -17.655 -96.110 ;
        RECT -17.335 -97.030 -17.165 -96.025 ;
        RECT -16.300 -96.120 -16.085 -95.165 ;
        RECT -24.235 -97.430 -19.195 -97.250 ;
        RECT -28.685 -97.450 -24.550 -97.445 ;
        RECT -17.360 -97.450 -17.145 -97.030 ;
        RECT -16.280 -97.065 -16.110 -96.120 ;
        RECT -15.790 -97.020 -15.620 -96.025 ;
        RECT -12.825 -96.220 -12.655 -94.385 ;
        RECT -12.230 -95.055 -11.535 -94.785 ;
        RECT -9.580 -94.960 -9.410 -94.385 ;
        RECT -9.105 -94.580 -8.935 -92.820 ;
        RECT -8.755 -94.210 -8.585 -92.475 ;
        RECT 0.275 -92.475 3.915 -92.305 ;
        RECT -7.855 -94.210 -7.685 -92.995 ;
        RECT -8.755 -94.380 -7.685 -94.210 ;
        RECT -6.875 -94.580 -6.705 -92.995 ;
        RECT -5.325 -93.960 -5.155 -92.995 ;
        RECT -3.780 -93.950 -3.610 -92.995 ;
        RECT -9.105 -94.750 -6.705 -94.580 ;
        RECT -6.440 -94.835 -5.745 -94.565 ;
        RECT -9.580 -95.130 -8.850 -94.960 ;
        RECT -9.020 -95.440 -8.850 -95.130 ;
        RECT -8.485 -95.205 -7.790 -94.935 ;
        RECT -12.235 -95.645 -10.580 -95.460 ;
        RECT -9.020 -95.610 -6.215 -95.440 ;
        RECT -12.235 -96.060 -12.050 -95.645 ;
        RECT -10.765 -95.765 -10.580 -95.645 ;
        RECT -10.765 -95.950 -9.985 -95.765 ;
        RECT -12.855 -96.900 -12.625 -96.220 ;
        RECT -12.225 -97.005 -12.055 -96.060 ;
        RECT -15.815 -97.450 -15.600 -97.020 ;
        RECT -31.240 -97.620 -24.550 -97.450 ;
        RECT -18.740 -97.620 -15.580 -97.450 ;
        RECT -12.245 -97.620 -12.050 -97.005 ;
        RECT -11.735 -97.250 -11.565 -96.025 ;
        RECT -10.170 -96.055 -9.985 -95.950 ;
        RECT -10.155 -97.065 -9.985 -96.055 ;
        RECT -9.675 -96.070 -8.175 -95.875 ;
        RECT -9.665 -97.065 -9.495 -96.070 ;
        RECT -8.345 -97.065 -8.175 -96.070 ;
        RECT -7.855 -97.065 -7.685 -95.610 ;
        RECT -6.875 -96.980 -6.705 -96.025 ;
        RECT -6.875 -97.250 -6.695 -96.980 ;
        RECT -6.385 -97.065 -6.215 -95.610 ;
        RECT -5.350 -95.655 -5.135 -93.960 ;
        RECT -3.800 -94.935 -3.585 -93.950 ;
        RECT 0.275 -94.035 0.445 -92.475 ;
        RECT -0.425 -94.215 -0.255 -94.210 ;
        RECT 0.765 -94.215 0.935 -92.995 ;
        RECT 1.255 -94.035 1.425 -92.475 ;
        RECT 1.855 -92.820 3.565 -92.650 ;
        RECT 1.855 -94.035 2.025 -92.820 ;
        RECT 2.345 -94.215 2.515 -92.995 ;
        RECT 2.835 -94.035 3.005 -92.820 ;
        RECT -0.425 -94.385 3.090 -94.215 ;
        RECT -3.365 -94.865 -2.670 -94.595 ;
        RECT -4.300 -95.165 -3.585 -94.935 ;
        RECT -5.830 -95.885 -5.135 -95.655 ;
        RECT -5.350 -96.110 -5.135 -95.885 ;
        RECT -5.325 -97.065 -5.155 -96.110 ;
        RECT -4.835 -97.030 -4.665 -96.025 ;
        RECT -3.800 -96.120 -3.585 -95.165 ;
        RECT -11.735 -97.430 -6.695 -97.250 ;
        RECT -4.860 -97.450 -4.645 -97.030 ;
        RECT -3.780 -97.065 -3.610 -96.120 ;
        RECT -3.290 -97.020 -3.120 -96.025 ;
        RECT -0.425 -96.220 -0.255 -94.385 ;
        RECT 0.270 -95.055 0.965 -94.785 ;
        RECT 2.920 -94.960 3.090 -94.385 ;
        RECT 3.395 -94.580 3.565 -92.820 ;
        RECT 3.745 -94.210 3.915 -92.475 ;
        RECT 12.775 -92.475 16.415 -92.305 ;
        RECT 4.645 -94.210 4.815 -92.995 ;
        RECT 3.745 -94.380 4.815 -94.210 ;
        RECT 5.625 -94.580 5.795 -92.995 ;
        RECT 7.175 -93.960 7.345 -92.995 ;
        RECT 8.720 -93.950 8.890 -92.995 ;
        RECT 3.395 -94.750 5.795 -94.580 ;
        RECT 6.060 -94.835 6.755 -94.565 ;
        RECT 2.920 -95.130 3.650 -94.960 ;
        RECT 3.480 -95.440 3.650 -95.130 ;
        RECT 4.015 -95.205 4.710 -94.935 ;
        RECT 0.265 -95.645 1.920 -95.460 ;
        RECT 3.480 -95.610 6.285 -95.440 ;
        RECT 0.265 -96.060 0.450 -95.645 ;
        RECT 1.735 -95.765 1.920 -95.645 ;
        RECT 1.735 -95.950 2.515 -95.765 ;
        RECT -0.455 -96.900 -0.225 -96.220 ;
        RECT 0.275 -97.005 0.445 -96.060 ;
        RECT -3.315 -97.450 -3.100 -97.020 ;
        RECT -6.240 -97.620 -3.080 -97.450 ;
        RECT 0.255 -97.620 0.450 -97.005 ;
        RECT 0.765 -97.250 0.935 -96.025 ;
        RECT 2.330 -96.055 2.515 -95.950 ;
        RECT 2.345 -97.065 2.515 -96.055 ;
        RECT 2.825 -96.070 4.325 -95.875 ;
        RECT 2.835 -97.065 3.005 -96.070 ;
        RECT 4.155 -97.065 4.325 -96.070 ;
        RECT 4.645 -97.065 4.815 -95.610 ;
        RECT 5.625 -96.980 5.795 -96.025 ;
        RECT 5.625 -97.250 5.805 -96.980 ;
        RECT 6.115 -97.065 6.285 -95.610 ;
        RECT 7.150 -95.655 7.365 -93.960 ;
        RECT 8.700 -94.935 8.915 -93.950 ;
        RECT 12.775 -94.035 12.945 -92.475 ;
        RECT 13.265 -94.215 13.435 -92.995 ;
        RECT 13.755 -94.035 13.925 -92.475 ;
        RECT 14.355 -92.820 16.065 -92.650 ;
        RECT 14.355 -94.035 14.525 -92.820 ;
        RECT 14.845 -94.215 15.015 -92.995 ;
        RECT 15.335 -94.035 15.505 -92.820 ;
        RECT 11.655 -94.385 15.590 -94.215 ;
        RECT 9.135 -94.865 9.830 -94.595 ;
        RECT 8.200 -95.165 8.915 -94.935 ;
        RECT 6.670 -95.885 7.365 -95.655 ;
        RECT 7.150 -96.110 7.365 -95.885 ;
        RECT 7.175 -97.065 7.345 -96.110 ;
        RECT 7.665 -97.030 7.835 -96.025 ;
        RECT 8.700 -96.120 8.915 -95.165 ;
        RECT 0.765 -97.430 5.805 -97.250 ;
        RECT 7.640 -97.450 7.855 -97.030 ;
        RECT 8.720 -97.065 8.890 -96.120 ;
        RECT 9.210 -97.020 9.380 -96.025 ;
        RECT 11.655 -96.215 11.825 -94.385 ;
        RECT 12.770 -95.055 13.465 -94.785 ;
        RECT 15.420 -94.960 15.590 -94.385 ;
        RECT 15.895 -94.580 16.065 -92.820 ;
        RECT 16.245 -94.210 16.415 -92.475 ;
        RECT 27.775 -92.475 31.415 -92.305 ;
        RECT 17.145 -94.210 17.315 -92.995 ;
        RECT 16.245 -94.380 17.315 -94.210 ;
        RECT 18.125 -94.580 18.295 -92.995 ;
        RECT 19.675 -93.960 19.845 -92.995 ;
        RECT 21.220 -93.950 21.390 -92.995 ;
        RECT 15.895 -94.750 18.295 -94.580 ;
        RECT 18.560 -94.835 19.255 -94.565 ;
        RECT 15.420 -95.130 16.150 -94.960 ;
        RECT 15.980 -95.440 16.150 -95.130 ;
        RECT 16.515 -95.205 17.210 -94.935 ;
        RECT 12.765 -95.645 14.420 -95.460 ;
        RECT 15.980 -95.610 18.785 -95.440 ;
        RECT 12.765 -96.060 12.950 -95.645 ;
        RECT 14.235 -95.765 14.420 -95.645 ;
        RECT 14.235 -95.950 15.015 -95.765 ;
        RECT 11.655 -96.220 11.830 -96.215 ;
        RECT 11.630 -96.900 11.860 -96.220 ;
        RECT 12.775 -97.005 12.945 -96.060 ;
        RECT 9.185 -97.450 9.400 -97.020 ;
        RECT 6.260 -97.620 9.420 -97.450 ;
        RECT 12.755 -97.620 12.950 -97.005 ;
        RECT 13.265 -97.250 13.435 -96.025 ;
        RECT 14.830 -96.055 15.015 -95.950 ;
        RECT 14.845 -97.065 15.015 -96.055 ;
        RECT 15.325 -96.070 16.825 -95.875 ;
        RECT 15.335 -97.065 15.505 -96.070 ;
        RECT 16.655 -97.065 16.825 -96.070 ;
        RECT 17.145 -97.065 17.315 -95.610 ;
        RECT 18.125 -96.980 18.295 -96.025 ;
        RECT 18.125 -97.250 18.305 -96.980 ;
        RECT 18.615 -97.065 18.785 -95.610 ;
        RECT 19.650 -95.655 19.865 -93.960 ;
        RECT 21.200 -94.935 21.415 -93.950 ;
        RECT 27.775 -94.035 27.945 -92.475 ;
        RECT 28.265 -94.215 28.435 -92.995 ;
        RECT 28.755 -94.035 28.925 -92.475 ;
        RECT 29.355 -92.820 31.065 -92.650 ;
        RECT 29.355 -94.035 29.525 -92.820 ;
        RECT 29.845 -94.215 30.015 -92.995 ;
        RECT 30.335 -94.035 30.505 -92.820 ;
        RECT 26.185 -94.385 30.590 -94.215 ;
        RECT 21.635 -94.865 22.330 -94.595 ;
        RECT 20.700 -95.165 21.415 -94.935 ;
        RECT 19.170 -95.885 19.865 -95.655 ;
        RECT 19.650 -96.110 19.865 -95.885 ;
        RECT 19.675 -97.065 19.845 -96.110 ;
        RECT 20.165 -97.030 20.335 -96.025 ;
        RECT 21.200 -96.120 21.415 -95.165 ;
        RECT 13.265 -97.430 18.305 -97.250 ;
        RECT 20.140 -97.450 20.355 -97.030 ;
        RECT 21.220 -97.065 21.390 -96.120 ;
        RECT 21.710 -97.020 21.880 -96.025 ;
        RECT 26.185 -96.220 26.355 -94.385 ;
        RECT 27.770 -95.055 28.465 -94.785 ;
        RECT 30.420 -94.960 30.590 -94.385 ;
        RECT 30.895 -94.580 31.065 -92.820 ;
        RECT 31.245 -94.210 31.415 -92.475 ;
        RECT 32.145 -94.210 32.315 -92.995 ;
        RECT 31.245 -94.380 32.315 -94.210 ;
        RECT 33.125 -94.580 33.295 -92.995 ;
        RECT 34.675 -93.960 34.845 -92.995 ;
        RECT 36.220 -93.950 36.390 -92.995 ;
        RECT 30.895 -94.750 33.295 -94.580 ;
        RECT 33.560 -94.835 34.255 -94.565 ;
        RECT 30.420 -95.130 31.150 -94.960 ;
        RECT 30.980 -95.440 31.150 -95.130 ;
        RECT 31.515 -95.205 32.210 -94.935 ;
        RECT 27.765 -95.645 29.420 -95.460 ;
        RECT 30.980 -95.610 33.785 -95.440 ;
        RECT 27.765 -96.060 27.950 -95.645 ;
        RECT 29.235 -95.765 29.420 -95.645 ;
        RECT 29.235 -95.950 30.015 -95.765 ;
        RECT 26.155 -96.900 26.385 -96.220 ;
        RECT 27.775 -97.005 27.945 -96.060 ;
        RECT 21.685 -97.450 21.900 -97.020 ;
        RECT 18.760 -97.620 21.920 -97.450 ;
        RECT 27.755 -97.620 27.950 -97.005 ;
        RECT 28.265 -97.250 28.435 -96.025 ;
        RECT 29.830 -96.055 30.015 -95.950 ;
        RECT 29.845 -97.065 30.015 -96.055 ;
        RECT 30.325 -96.070 31.825 -95.875 ;
        RECT 30.335 -97.065 30.505 -96.070 ;
        RECT 31.655 -97.065 31.825 -96.070 ;
        RECT 32.145 -97.065 32.315 -95.610 ;
        RECT 33.125 -96.980 33.295 -96.025 ;
        RECT 33.125 -97.250 33.305 -96.980 ;
        RECT 33.615 -97.065 33.785 -95.610 ;
        RECT 34.650 -95.655 34.865 -93.960 ;
        RECT 36.200 -94.935 36.415 -93.950 ;
        RECT 36.635 -94.865 37.330 -94.595 ;
        RECT 35.700 -95.165 36.415 -94.935 ;
        RECT 34.170 -95.885 34.865 -95.655 ;
        RECT 34.650 -96.110 34.865 -95.885 ;
        RECT 34.675 -97.065 34.845 -96.110 ;
        RECT 35.165 -97.030 35.335 -96.025 ;
        RECT 36.200 -96.120 36.415 -95.165 ;
        RECT 28.265 -97.430 33.305 -97.250 ;
        RECT 35.140 -97.360 35.355 -97.030 ;
        RECT 36.220 -97.065 36.390 -96.120 ;
        RECT 36.710 -97.020 36.880 -96.025 ;
        RECT 36.685 -97.360 36.900 -97.020 ;
        RECT 37.715 -97.360 39.020 -88.055 ;
        RECT 80.790 -89.675 81.775 -88.770 ;
        RECT 79.070 -92.050 80.475 -91.005 ;
        RECT 40.140 -93.065 41.140 -92.895 ;
        RECT 77.270 -93.065 79.080 -92.835 ;
        RECT 40.140 -93.925 79.080 -93.065 ;
        RECT 40.140 -94.750 41.140 -93.925 ;
        RECT 77.270 -94.190 79.080 -93.925 ;
        RECT 33.680 -97.620 39.020 -97.360 ;
        RECT 76.070 -97.555 77.530 -97.550 ;
        RECT -37.245 -97.880 39.020 -97.620 ;
        RECT -37.245 -97.885 -28.080 -97.880 ;
        RECT -24.745 -97.885 39.020 -97.880 ;
        RECT -35.085 -97.985 -32.415 -97.885 ;
        RECT -31.240 -97.930 -28.080 -97.885 ;
        RECT -18.740 -97.930 -15.580 -97.885 ;
        RECT -6.240 -97.930 -3.080 -97.885 ;
        RECT 6.260 -97.930 9.420 -97.885 ;
        RECT 18.760 -97.930 21.920 -97.885 ;
        RECT -35.040 -98.780 -34.870 -97.985 ;
        RECT -34.550 -98.700 -34.380 -98.240 ;
        RECT -34.580 -99.165 -34.350 -98.700 ;
        RECT -34.060 -98.780 -33.890 -97.985 ;
        RECT -33.570 -98.700 -33.400 -98.240 ;
        RECT -33.600 -99.165 -33.370 -98.700 ;
        RECT -33.080 -98.780 -32.910 -97.985 ;
        RECT 33.680 -97.995 39.020 -97.885 ;
        RECT -32.590 -98.700 -32.420 -98.240 ;
        RECT -12.030 -98.310 -11.350 -98.080 ;
        RECT 0.455 -98.160 1.135 -98.145 ;
        RECT -11.595 -98.550 -11.350 -98.310 ;
        RECT 0.290 -98.330 11.145 -98.160 ;
        RECT 0.455 -98.375 1.135 -98.330 ;
        RECT -32.620 -99.005 -32.390 -98.700 ;
        RECT -27.505 -99.005 -27.275 -98.675 ;
        RECT -11.595 -98.730 10.665 -98.550 ;
        RECT -32.620 -99.165 -27.275 -99.005 ;
        RECT -34.580 -99.355 -27.275 -99.165 ;
        RECT 10.485 -99.290 10.665 -98.730 ;
        RECT 10.975 -98.950 11.145 -98.330 ;
        RECT 25.895 -98.410 26.575 -98.380 ;
        RECT 11.370 -98.505 12.050 -98.460 ;
        RECT 11.370 -98.675 25.375 -98.505 ;
        RECT 25.895 -98.580 27.255 -98.410 ;
        RECT 25.895 -98.610 26.575 -98.580 ;
        RECT 11.370 -98.690 12.050 -98.675 ;
        RECT 25.205 -98.870 25.375 -98.675 ;
        RECT 10.975 -99.120 18.485 -98.950 ;
        RECT 25.205 -99.040 26.905 -98.870 ;
        RECT -34.580 -99.395 -32.390 -99.355 ;
        RECT -34.580 -100.660 -34.350 -99.395 ;
        RECT -33.600 -99.720 -33.370 -99.395 ;
        RECT -32.620 -99.720 -32.390 -99.395 ;
        RECT 10.485 -99.470 18.090 -99.290 ;
        RECT -34.550 -100.680 -34.380 -100.660 ;
        RECT -33.570 -100.680 -33.400 -99.720 ;
        RECT -32.590 -100.680 -32.420 -99.720 ;
        RECT -25.595 -100.410 -25.365 -99.730 ;
        RECT -25.580 -101.675 -25.380 -100.410 ;
        RECT -25.580 -101.905 -24.900 -101.675 ;
        RECT 9.665 -101.895 10.345 -101.665 ;
        RECT -37.980 -102.315 -37.300 -102.085 ;
        RECT 9.145 -102.315 9.920 -102.085 ;
        RECT -6.815 -102.770 -6.130 -102.515 ;
        RECT -31.670 -104.060 -28.530 -103.890 ;
        RECT -36.325 -105.115 -36.155 -104.155 ;
        RECT -35.345 -105.115 -35.175 -104.155 ;
        RECT -34.365 -104.175 -34.195 -104.155 ;
        RECT -36.355 -105.440 -36.125 -105.115 ;
        RECT -35.375 -105.440 -35.145 -105.115 ;
        RECT -34.395 -105.440 -34.165 -104.175 ;
        RECT -32.135 -104.730 -31.965 -104.230 ;
        RECT -31.670 -104.315 -31.460 -104.060 ;
        RECT -36.355 -105.480 -34.165 -105.440 ;
        RECT -36.505 -105.525 -34.165 -105.480 ;
        RECT -32.160 -104.950 -31.950 -104.730 ;
        RECT -31.645 -104.770 -31.475 -104.315 ;
        RECT -31.155 -104.680 -30.985 -104.230 ;
        RECT -30.690 -104.340 -30.480 -104.060 ;
        RECT -31.160 -104.950 -30.980 -104.680 ;
        RECT -30.665 -104.770 -30.495 -104.340 ;
        RECT -30.175 -104.680 -30.005 -104.230 ;
        RECT -29.720 -104.335 -29.510 -104.060 ;
        RECT -30.190 -104.770 -30.005 -104.680 ;
        RECT -29.685 -104.770 -29.515 -104.335 ;
        RECT -29.195 -104.690 -29.025 -104.230 ;
        RECT -28.710 -104.285 -28.530 -104.060 ;
        RECT -18.170 -104.060 -15.030 -103.890 ;
        RECT -28.705 -104.655 -28.535 -104.285 ;
        RECT -30.190 -104.950 -30.010 -104.770 ;
        RECT -29.200 -104.950 -29.020 -104.690 ;
        RECT -32.160 -105.120 -29.020 -104.950 ;
        RECT -36.915 -105.535 -34.165 -105.525 ;
        RECT -36.920 -105.670 -34.165 -105.535 ;
        RECT -36.920 -105.720 -36.125 -105.670 ;
        RECT -36.920 -107.510 -36.680 -105.720 ;
        RECT -36.505 -105.830 -36.125 -105.720 ;
        RECT -36.355 -106.135 -36.125 -105.830 ;
        RECT -36.325 -106.595 -36.155 -106.135 ;
        RECT -35.835 -106.850 -35.665 -106.055 ;
        RECT -35.375 -106.135 -35.145 -105.670 ;
        RECT -35.345 -106.595 -35.175 -106.135 ;
        RECT -34.855 -106.850 -34.685 -106.055 ;
        RECT -34.395 -106.135 -34.165 -105.670 ;
        RECT -33.985 -105.545 -33.145 -105.515 ;
        RECT -32.160 -105.545 -31.285 -105.120 ;
        RECT -28.740 -105.390 -28.505 -104.655 ;
        RECT -28.285 -105.360 -27.915 -104.520 ;
        RECT -27.610 -105.115 -27.440 -104.155 ;
        RECT -26.630 -105.115 -26.460 -104.155 ;
        RECT -25.650 -104.175 -25.480 -104.155 ;
        RECT -33.985 -105.810 -31.285 -105.545 ;
        RECT -29.365 -105.760 -28.505 -105.390 ;
        RECT -33.985 -105.885 -33.145 -105.810 ;
        RECT -32.160 -105.955 -31.285 -105.810 ;
        RECT -34.365 -106.595 -34.195 -106.135 ;
        RECT -33.875 -106.850 -33.705 -106.055 ;
        RECT -32.160 -106.125 -29.005 -105.955 ;
        RECT -32.160 -106.160 -31.950 -106.125 ;
        RECT -32.155 -106.375 -31.950 -106.160 ;
        RECT -32.135 -106.845 -31.965 -106.375 ;
        RECT -31.645 -106.785 -31.475 -106.305 ;
        RECT -31.170 -106.370 -30.965 -106.125 ;
        RECT -36.330 -107.190 -33.660 -106.850 ;
        RECT -31.675 -107.075 -31.455 -106.785 ;
        RECT -31.155 -106.845 -30.985 -106.370 ;
        RECT -30.665 -106.730 -30.495 -106.305 ;
        RECT -30.200 -106.370 -29.995 -106.125 ;
        RECT -30.690 -107.075 -30.470 -106.730 ;
        RECT -30.175 -106.845 -30.005 -106.370 ;
        RECT -29.685 -106.730 -29.515 -106.305 ;
        RECT -29.210 -106.330 -29.005 -106.125 ;
        RECT -29.710 -107.075 -29.490 -106.730 ;
        RECT -29.195 -106.845 -29.025 -106.330 ;
        RECT -28.740 -106.435 -28.505 -105.760 ;
        RECT -28.280 -105.480 -27.915 -105.360 ;
        RECT -27.640 -105.440 -27.410 -105.115 ;
        RECT -26.660 -105.440 -26.430 -105.115 ;
        RECT -25.680 -105.440 -25.450 -104.175 ;
        RECT -24.660 -104.655 -24.375 -104.265 ;
        RECT -24.660 -104.880 -23.355 -104.655 ;
        RECT -24.660 -105.085 -24.375 -104.880 ;
        RECT -27.640 -105.480 -25.450 -105.440 ;
        RECT -28.280 -105.670 -25.450 -105.480 ;
        RECT -28.280 -105.830 -27.410 -105.670 ;
        RECT -27.640 -106.135 -27.410 -105.830 ;
        RECT -28.705 -106.785 -28.535 -106.435 ;
        RECT -27.610 -106.595 -27.440 -106.135 ;
        RECT -28.730 -107.075 -28.510 -106.785 ;
        RECT -27.120 -106.850 -26.950 -106.055 ;
        RECT -26.660 -106.135 -26.430 -105.670 ;
        RECT -26.630 -106.595 -26.460 -106.135 ;
        RECT -26.140 -106.850 -25.970 -106.055 ;
        RECT -25.680 -106.135 -25.450 -105.670 ;
        RECT -25.270 -105.570 -24.430 -105.515 ;
        RECT -23.580 -105.550 -23.355 -104.880 ;
        RECT -22.825 -105.115 -22.655 -104.155 ;
        RECT -21.845 -105.115 -21.675 -104.155 ;
        RECT -20.865 -104.175 -20.695 -104.155 ;
        RECT -22.855 -105.440 -22.625 -105.115 ;
        RECT -21.875 -105.440 -21.645 -105.115 ;
        RECT -20.895 -105.440 -20.665 -104.175 ;
        RECT -18.635 -104.730 -18.465 -104.230 ;
        RECT -18.170 -104.315 -17.960 -104.060 ;
        RECT -22.855 -105.480 -20.665 -105.440 ;
        RECT -23.005 -105.550 -20.665 -105.480 ;
        RECT -18.660 -104.950 -18.450 -104.730 ;
        RECT -18.145 -104.770 -17.975 -104.315 ;
        RECT -17.655 -104.680 -17.485 -104.230 ;
        RECT -17.190 -104.340 -16.980 -104.060 ;
        RECT -17.660 -104.950 -17.480 -104.680 ;
        RECT -17.165 -104.770 -16.995 -104.340 ;
        RECT -16.675 -104.680 -16.505 -104.230 ;
        RECT -16.220 -104.335 -16.010 -104.060 ;
        RECT -16.690 -104.770 -16.505 -104.680 ;
        RECT -16.185 -104.770 -16.015 -104.335 ;
        RECT -15.695 -104.690 -15.525 -104.230 ;
        RECT -15.210 -104.285 -15.030 -104.060 ;
        RECT -15.205 -104.655 -15.035 -104.285 ;
        RECT -16.690 -104.950 -16.510 -104.770 ;
        RECT -15.700 -104.950 -15.520 -104.690 ;
        RECT -18.660 -105.120 -15.520 -104.950 ;
        RECT -24.130 -105.570 -23.830 -105.565 ;
        RECT -25.270 -105.860 -23.830 -105.570 ;
        RECT -23.580 -105.670 -20.665 -105.550 ;
        RECT -23.580 -105.775 -22.625 -105.670 ;
        RECT -25.270 -105.885 -24.430 -105.860 ;
        RECT -25.650 -106.595 -25.480 -106.135 ;
        RECT -25.160 -106.850 -24.990 -106.055 ;
        RECT -24.130 -106.225 -23.830 -105.860 ;
        RECT -23.555 -106.350 -23.255 -105.775 ;
        RECT -23.005 -105.830 -22.625 -105.775 ;
        RECT -22.855 -106.135 -22.625 -105.830 ;
        RECT -22.825 -106.595 -22.655 -106.135 ;
        RECT -22.335 -106.850 -22.165 -106.055 ;
        RECT -21.875 -106.135 -21.645 -105.670 ;
        RECT -21.845 -106.595 -21.675 -106.135 ;
        RECT -21.355 -106.850 -21.185 -106.055 ;
        RECT -20.895 -106.135 -20.665 -105.670 ;
        RECT -20.485 -105.560 -19.645 -105.515 ;
        RECT -18.660 -105.560 -17.785 -105.120 ;
        RECT -15.240 -105.390 -15.005 -104.655 ;
        RECT -14.785 -105.360 -14.415 -104.520 ;
        RECT -14.110 -105.115 -13.940 -104.155 ;
        RECT -13.130 -105.115 -12.960 -104.155 ;
        RECT -12.150 -104.175 -11.980 -104.155 ;
        RECT -20.485 -105.845 -17.785 -105.560 ;
        RECT -15.865 -105.760 -15.005 -105.390 ;
        RECT -20.485 -105.885 -19.645 -105.845 ;
        RECT -18.660 -105.955 -17.785 -105.845 ;
        RECT -20.865 -106.595 -20.695 -106.135 ;
        RECT -20.375 -106.850 -20.205 -106.055 ;
        RECT -18.660 -106.125 -15.505 -105.955 ;
        RECT -18.660 -106.160 -18.450 -106.125 ;
        RECT -18.655 -106.325 -18.450 -106.160 ;
        RECT -18.655 -106.375 -18.420 -106.325 ;
        RECT -31.675 -107.245 -28.510 -107.075 ;
        RECT -27.615 -107.190 -20.160 -106.850 ;
        RECT -18.650 -106.985 -18.420 -106.375 ;
        RECT -18.145 -106.785 -17.975 -106.305 ;
        RECT -17.670 -106.370 -17.465 -106.125 ;
        RECT -18.175 -107.075 -17.955 -106.785 ;
        RECT -17.655 -106.845 -17.485 -106.370 ;
        RECT -17.165 -106.730 -16.995 -106.305 ;
        RECT -16.700 -106.370 -16.495 -106.125 ;
        RECT -17.190 -107.075 -16.970 -106.730 ;
        RECT -16.675 -106.845 -16.505 -106.370 ;
        RECT -16.185 -106.730 -16.015 -106.305 ;
        RECT -15.710 -106.330 -15.505 -106.125 ;
        RECT -16.210 -107.075 -15.990 -106.730 ;
        RECT -15.695 -106.845 -15.525 -106.330 ;
        RECT -15.240 -106.435 -15.005 -105.760 ;
        RECT -14.780 -105.480 -14.415 -105.360 ;
        RECT -14.140 -105.440 -13.910 -105.115 ;
        RECT -13.160 -105.440 -12.930 -105.115 ;
        RECT -12.180 -105.440 -11.950 -104.175 ;
        RECT -11.160 -105.085 -10.875 -104.265 ;
        RECT -9.700 -105.115 -9.530 -104.155 ;
        RECT -8.720 -105.115 -8.550 -104.155 ;
        RECT -7.740 -104.175 -7.570 -104.155 ;
        RECT -14.140 -105.480 -11.950 -105.440 ;
        RECT -9.730 -105.440 -9.500 -105.115 ;
        RECT -8.750 -105.440 -8.520 -105.115 ;
        RECT -7.770 -105.440 -7.540 -104.175 ;
        RECT -9.730 -105.480 -7.540 -105.440 ;
        RECT -14.780 -105.670 -11.950 -105.480 ;
        RECT -14.780 -105.830 -13.910 -105.670 ;
        RECT -15.205 -106.785 -15.035 -106.435 ;
        RECT -15.230 -107.075 -15.010 -106.785 ;
        RECT -18.175 -107.245 -15.010 -107.075 ;
        RECT -14.785 -106.810 -14.415 -106.015 ;
        RECT -14.140 -106.135 -13.910 -105.830 ;
        RECT -14.110 -106.595 -13.940 -106.135 ;
        RECT -33.240 -107.425 -32.580 -107.360 ;
        RECT -14.785 -107.425 -14.410 -106.810 ;
        RECT -13.620 -106.850 -13.450 -106.055 ;
        RECT -13.160 -106.135 -12.930 -105.670 ;
        RECT -13.130 -106.595 -12.960 -106.135 ;
        RECT -12.640 -106.850 -12.470 -106.055 ;
        RECT -12.180 -106.135 -11.950 -105.670 ;
        RECT -11.770 -105.570 -10.930 -105.515 ;
        RECT -11.770 -105.860 -10.755 -105.570 ;
        RECT -10.470 -105.590 -10.170 -105.570 ;
        RECT -9.880 -105.590 -7.540 -105.480 ;
        RECT -6.815 -105.515 -6.620 -102.770 ;
        RECT -10.470 -105.670 -7.540 -105.590 ;
        RECT -10.470 -105.800 -9.500 -105.670 ;
        RECT -11.770 -105.885 -10.930 -105.860 ;
        RECT -12.150 -106.595 -11.980 -106.135 ;
        RECT -11.660 -106.850 -11.490 -106.055 ;
        RECT -10.470 -106.230 -10.170 -105.800 ;
        RECT -9.880 -105.830 -9.500 -105.800 ;
        RECT -9.730 -106.135 -9.500 -105.830 ;
        RECT -9.700 -106.595 -9.530 -106.135 ;
        RECT -9.210 -106.850 -9.040 -106.055 ;
        RECT -8.750 -106.135 -8.520 -105.670 ;
        RECT -8.720 -106.595 -8.550 -106.135 ;
        RECT -8.230 -106.850 -8.060 -106.055 ;
        RECT -7.770 -106.135 -7.540 -105.670 ;
        RECT -7.360 -105.885 -6.520 -105.515 ;
        RECT -7.740 -106.595 -7.570 -106.135 ;
        RECT -7.250 -106.850 -7.080 -106.055 ;
        RECT -14.115 -107.190 -7.035 -106.850 ;
        RECT -6.815 -107.425 -6.620 -105.885 ;
        RECT -5.050 -106.290 -4.880 -104.240 ;
        RECT -1.360 -105.460 -1.190 -104.240 ;
        RECT -0.380 -105.460 -0.210 -104.240 ;
        RECT 0.600 -105.460 0.770 -104.240 ;
        RECT -2.005 -105.645 0.770 -105.460 ;
        RECT 1.700 -105.475 1.930 -105.055 ;
        RECT 3.615 -105.165 3.785 -104.305 ;
        RECT 4.595 -104.845 4.765 -104.305 ;
        RECT 5.575 -104.845 5.745 -104.305 ;
        RECT -5.805 -106.555 -4.880 -106.290 ;
        RECT -4.705 -106.335 -4.030 -106.285 ;
        RECT -2.005 -106.335 -1.820 -105.645 ;
        RECT 0.970 -105.745 1.930 -105.475 ;
        RECT 2.930 -105.515 3.785 -105.165 ;
        RECT 5.970 -105.080 6.335 -105.015 ;
        RECT 5.970 -105.220 6.835 -105.080 ;
        RECT 5.970 -105.285 6.945 -105.220 ;
        RECT 5.970 -105.315 6.335 -105.285 ;
        RECT -0.710 -105.930 -0.035 -105.885 ;
        RECT 2.105 -105.930 2.785 -105.925 ;
        RECT -0.710 -106.120 2.785 -105.930 ;
        RECT -0.710 -106.155 -0.035 -106.120 ;
        RECT 2.105 -106.155 2.785 -106.120 ;
        RECT -4.705 -106.520 -1.820 -106.335 ;
        RECT -4.705 -106.555 -4.030 -106.520 ;
        RECT -38.700 -107.955 -37.780 -107.640 ;
        RECT -38.595 -107.960 -37.780 -107.955 ;
        RECT -36.925 -108.195 -36.625 -107.510 ;
        RECT -35.270 -107.620 -6.620 -107.425 ;
        RECT -33.240 -107.660 -32.580 -107.620 ;
        RECT -24.375 -107.855 -23.690 -107.805 ;
        RECT -19.645 -107.855 -18.985 -107.800 ;
        RECT -9.575 -107.855 -8.915 -107.805 ;
        RECT -35.270 -108.050 -8.915 -107.855 ;
        RECT -24.375 -108.105 -23.690 -108.050 ;
        RECT -19.645 -108.100 -18.985 -108.050 ;
        RECT -9.575 -108.105 -8.915 -108.050 ;
        RECT -36.920 -110.055 -36.680 -108.195 ;
        RECT -35.185 -108.315 -34.500 -108.250 ;
        RECT -22.200 -108.315 -21.515 -108.220 ;
        RECT -8.360 -108.315 -7.700 -108.220 ;
        RECT -35.270 -108.510 -7.695 -108.315 ;
        RECT -35.185 -108.550 -34.500 -108.510 ;
        RECT -35.130 -108.750 -34.575 -108.550 ;
        RECT -31.075 -108.750 -30.520 -108.510 ;
        RECT -22.200 -108.520 -21.515 -108.510 ;
        RECT -36.370 -109.090 -29.515 -108.750 ;
        RECT -28.620 -108.865 -25.455 -108.695 ;
        RECT -22.085 -108.750 -21.530 -108.520 ;
        RECT -21.170 -108.750 -18.570 -108.740 ;
        RECT -17.695 -108.750 -17.140 -108.510 ;
        RECT -36.325 -109.885 -36.155 -109.090 ;
        RECT -35.835 -109.805 -35.665 -109.345 ;
        RECT -36.920 -110.275 -36.045 -110.055 ;
        RECT -36.885 -110.425 -36.045 -110.275 ;
        RECT -35.865 -110.270 -35.635 -109.805 ;
        RECT -35.345 -109.885 -35.175 -109.090 ;
        RECT -34.855 -109.805 -34.685 -109.345 ;
        RECT -34.885 -110.270 -34.655 -109.805 ;
        RECT -34.365 -109.885 -34.195 -109.090 ;
        RECT -33.875 -109.805 -33.705 -109.345 ;
        RECT -33.905 -110.110 -33.675 -109.805 ;
        RECT -33.060 -110.055 -32.760 -109.335 ;
        RECT -32.140 -109.885 -31.970 -109.090 ;
        RECT -31.650 -109.805 -31.480 -109.345 ;
        RECT -33.905 -110.270 -33.240 -110.110 ;
        RECT -66.000 -112.485 -65.325 -112.455 ;
        RECT -66.100 -112.495 -65.325 -112.485 ;
        RECT -97.425 -113.695 -79.735 -112.665 ;
        RECT -67.135 -112.675 -65.325 -112.495 ;
        RECT -65.085 -112.570 -62.935 -112.420 ;
        RECT -65.085 -112.610 -62.990 -112.570 ;
        RECT -62.040 -112.630 -61.870 -111.850 ;
        RECT -61.550 -112.390 -61.380 -111.850 ;
        RECT -61.060 -112.630 -60.890 -111.850 ;
        RECT -60.570 -112.390 -60.400 -111.850 ;
        RECT -60.080 -111.905 -58.220 -111.555 ;
        RECT -35.865 -110.460 -33.240 -110.270 ;
        RECT -33.060 -110.365 -31.860 -110.055 ;
        RECT -32.875 -110.370 -31.860 -110.365 ;
        RECT -32.700 -110.425 -31.860 -110.370 ;
        RECT -31.680 -110.270 -31.450 -109.805 ;
        RECT -31.160 -109.885 -30.990 -109.090 ;
        RECT -30.670 -109.805 -30.500 -109.345 ;
        RECT -30.700 -110.270 -30.470 -109.805 ;
        RECT -30.180 -109.885 -30.010 -109.090 ;
        RECT -28.620 -109.155 -28.400 -108.865 ;
        RECT -29.690 -109.805 -29.520 -109.345 ;
        RECT -28.595 -109.505 -28.425 -109.155 ;
        RECT -29.720 -110.110 -29.490 -109.805 ;
        RECT -29.720 -110.270 -28.850 -110.110 ;
        RECT -35.865 -110.500 -33.675 -110.460 ;
        RECT -35.865 -111.765 -35.635 -110.500 ;
        RECT -34.885 -110.825 -34.655 -110.500 ;
        RECT -33.905 -110.825 -33.675 -110.500 ;
        RECT -35.835 -111.785 -35.665 -111.765 ;
        RECT -34.855 -111.785 -34.685 -110.825 ;
        RECT -33.875 -111.785 -33.705 -110.825 ;
        RECT -33.470 -111.110 -33.240 -110.460 ;
        RECT -31.680 -110.460 -28.850 -110.270 ;
        RECT -31.680 -110.500 -29.490 -110.460 ;
        RECT -32.755 -111.110 -32.470 -110.855 ;
        RECT -33.470 -111.355 -32.470 -111.110 ;
        RECT -32.755 -111.675 -32.470 -111.355 ;
        RECT -31.680 -111.765 -31.450 -110.500 ;
        RECT -30.700 -110.825 -30.470 -110.500 ;
        RECT -29.720 -110.825 -29.490 -110.500 ;
        RECT -29.215 -110.580 -28.850 -110.460 ;
        RECT -28.625 -110.180 -28.390 -109.505 ;
        RECT -28.105 -109.610 -27.935 -109.095 ;
        RECT -27.640 -109.210 -27.420 -108.865 ;
        RECT -28.125 -109.815 -27.920 -109.610 ;
        RECT -27.615 -109.635 -27.445 -109.210 ;
        RECT -27.125 -109.570 -26.955 -109.095 ;
        RECT -26.660 -109.210 -26.440 -108.865 ;
        RECT -27.135 -109.815 -26.930 -109.570 ;
        RECT -26.635 -109.635 -26.465 -109.210 ;
        RECT -26.145 -109.570 -25.975 -109.095 ;
        RECT -25.675 -109.155 -25.455 -108.865 ;
        RECT -22.870 -109.080 -16.015 -108.750 ;
        RECT -22.870 -109.090 -20.200 -109.080 ;
        RECT -18.685 -109.090 -16.015 -109.080 ;
        RECT -15.120 -108.865 -11.955 -108.695 ;
        RECT -26.165 -109.815 -25.960 -109.570 ;
        RECT -25.655 -109.635 -25.485 -109.155 ;
        RECT -25.165 -109.565 -24.995 -109.095 ;
        RECT -25.180 -109.780 -24.975 -109.565 ;
        RECT -25.180 -109.815 -24.970 -109.780 ;
        RECT -28.125 -109.985 -24.970 -109.815 ;
        RECT -22.825 -109.885 -22.655 -109.090 ;
        RECT -22.335 -109.805 -22.165 -109.345 ;
        RECT -28.625 -110.550 -27.765 -110.180 ;
        RECT -25.845 -110.285 -24.515 -109.985 ;
        RECT -23.385 -110.090 -22.545 -110.055 ;
        RECT -31.650 -111.785 -31.480 -111.765 ;
        RECT -30.670 -111.785 -30.500 -110.825 ;
        RECT -29.690 -111.785 -29.520 -110.825 ;
        RECT -29.215 -111.420 -28.845 -110.580 ;
        RECT -28.625 -111.285 -28.390 -110.550 ;
        RECT -25.845 -110.820 -24.970 -110.285 ;
        RECT -23.495 -110.390 -22.545 -110.090 ;
        RECT -23.385 -110.425 -22.545 -110.390 ;
        RECT -22.365 -110.270 -22.135 -109.805 ;
        RECT -21.845 -109.885 -21.675 -109.090 ;
        RECT -21.355 -109.805 -21.185 -109.345 ;
        RECT -21.385 -110.270 -21.155 -109.805 ;
        RECT -20.865 -109.885 -20.695 -109.090 ;
        RECT -20.375 -109.805 -20.205 -109.345 ;
        RECT -20.405 -110.110 -20.175 -109.805 ;
        RECT -19.500 -110.055 -19.200 -109.260 ;
        RECT -18.640 -109.885 -18.470 -109.090 ;
        RECT -18.150 -109.805 -17.980 -109.345 ;
        RECT -20.405 -110.270 -19.685 -110.110 ;
        RECT -28.110 -110.990 -24.970 -110.820 ;
        RECT -28.110 -111.250 -27.930 -110.990 ;
        RECT -27.120 -111.170 -26.940 -110.990 ;
        RECT -28.595 -111.655 -28.425 -111.285 ;
        RECT -28.600 -111.880 -28.420 -111.655 ;
        RECT -28.105 -111.710 -27.935 -111.250 ;
        RECT -27.615 -111.605 -27.445 -111.170 ;
        RECT -27.125 -111.260 -26.940 -111.170 ;
        RECT -27.620 -111.880 -27.410 -111.605 ;
        RECT -27.125 -111.710 -26.955 -111.260 ;
        RECT -26.635 -111.600 -26.465 -111.170 ;
        RECT -26.150 -111.260 -25.970 -110.990 ;
        RECT -26.650 -111.880 -26.440 -111.600 ;
        RECT -26.145 -111.710 -25.975 -111.260 ;
        RECT -25.655 -111.625 -25.485 -111.170 ;
        RECT -25.180 -111.210 -24.970 -110.990 ;
        RECT -22.365 -110.460 -19.685 -110.270 ;
        RECT -19.500 -110.370 -18.360 -110.055 ;
        RECT -19.200 -110.425 -18.360 -110.370 ;
        RECT -18.180 -110.270 -17.950 -109.805 ;
        RECT -17.660 -109.885 -17.490 -109.090 ;
        RECT -17.170 -109.805 -17.000 -109.345 ;
        RECT -17.200 -110.270 -16.970 -109.805 ;
        RECT -16.680 -109.885 -16.510 -109.090 ;
        RECT -15.120 -109.155 -14.900 -108.865 ;
        RECT -16.190 -109.805 -16.020 -109.345 ;
        RECT -15.095 -109.505 -14.925 -109.155 ;
        RECT -16.220 -110.110 -15.990 -109.805 ;
        RECT -16.220 -110.270 -15.350 -110.110 ;
        RECT -22.365 -110.500 -20.175 -110.460 ;
        RECT -25.670 -111.880 -25.460 -111.625 ;
        RECT -25.165 -111.710 -24.995 -111.210 ;
        RECT -22.365 -111.765 -22.135 -110.500 ;
        RECT -21.385 -110.825 -21.155 -110.500 ;
        RECT -20.405 -110.825 -20.175 -110.500 ;
        RECT -22.335 -111.785 -22.165 -111.765 ;
        RECT -21.355 -111.785 -21.185 -110.825 ;
        RECT -20.375 -111.785 -20.205 -110.825 ;
        RECT -19.995 -111.105 -19.685 -110.460 ;
        RECT -18.180 -110.460 -15.350 -110.270 ;
        RECT -18.180 -110.500 -15.990 -110.460 ;
        RECT -19.255 -111.105 -18.970 -110.855 ;
        RECT -19.995 -111.415 -18.970 -111.105 ;
        RECT -19.255 -111.675 -18.970 -111.415 ;
        RECT -18.180 -111.765 -17.950 -110.500 ;
        RECT -17.200 -110.825 -16.970 -110.500 ;
        RECT -16.220 -110.825 -15.990 -110.500 ;
        RECT -15.715 -110.580 -15.350 -110.460 ;
        RECT -15.125 -110.180 -14.890 -109.505 ;
        RECT -14.605 -109.610 -14.435 -109.095 ;
        RECT -14.140 -109.210 -13.920 -108.865 ;
        RECT -14.625 -109.815 -14.420 -109.610 ;
        RECT -14.115 -109.635 -13.945 -109.210 ;
        RECT -13.625 -109.570 -13.455 -109.095 ;
        RECT -13.160 -109.210 -12.940 -108.865 ;
        RECT -13.635 -109.815 -13.430 -109.570 ;
        RECT -13.135 -109.635 -12.965 -109.210 ;
        RECT -12.645 -109.570 -12.475 -109.095 ;
        RECT -12.175 -109.155 -11.955 -108.865 ;
        RECT -12.665 -109.815 -12.460 -109.570 ;
        RECT -12.155 -109.635 -11.985 -109.155 ;
        RECT -11.665 -109.565 -11.495 -109.095 ;
        RECT -11.680 -109.780 -11.475 -109.565 ;
        RECT -11.680 -109.815 -11.470 -109.780 ;
        RECT -14.625 -109.975 -11.470 -109.815 ;
        RECT -14.625 -109.985 -11.095 -109.975 ;
        RECT -15.125 -110.550 -14.265 -110.180 ;
        RECT -12.345 -110.275 -11.095 -109.985 ;
        RECT -18.150 -111.785 -17.980 -111.765 ;
        RECT -17.170 -111.785 -17.000 -110.825 ;
        RECT -16.190 -111.785 -16.020 -110.825 ;
        RECT -15.715 -111.420 -15.345 -110.580 ;
        RECT -15.125 -111.285 -14.890 -110.550 ;
        RECT -12.345 -110.820 -11.470 -110.275 ;
        RECT -14.610 -110.990 -11.470 -110.820 ;
        RECT -14.610 -111.250 -14.430 -110.990 ;
        RECT -13.620 -111.170 -13.440 -110.990 ;
        RECT -15.095 -111.655 -14.925 -111.285 ;
        RECT -28.600 -112.050 -25.460 -111.880 ;
        RECT -15.100 -111.880 -14.920 -111.655 ;
        RECT -14.605 -111.710 -14.435 -111.250 ;
        RECT -14.115 -111.605 -13.945 -111.170 ;
        RECT -13.625 -111.260 -13.440 -111.170 ;
        RECT -14.120 -111.880 -13.910 -111.605 ;
        RECT -13.625 -111.710 -13.455 -111.260 ;
        RECT -13.135 -111.600 -12.965 -111.170 ;
        RECT -12.650 -111.260 -12.470 -110.990 ;
        RECT -13.150 -111.880 -12.940 -111.600 ;
        RECT -12.645 -111.710 -12.475 -111.260 ;
        RECT -12.155 -111.625 -11.985 -111.170 ;
        RECT -11.680 -111.210 -11.470 -110.990 ;
        RECT -12.170 -111.880 -11.960 -111.625 ;
        RECT -11.665 -111.710 -11.495 -111.210 ;
        RECT -10.275 -111.410 -8.785 -108.510 ;
        RECT -8.360 -108.520 -7.700 -108.510 ;
        RECT -5.050 -108.820 -4.880 -106.555 ;
        RECT -2.005 -106.790 -1.820 -106.520 ;
        RECT -1.650 -106.340 -0.975 -106.275 ;
        RECT 2.960 -106.340 3.130 -105.515 ;
        RECT 4.105 -106.000 4.275 -105.460 ;
        RECT 4.595 -106.240 4.765 -105.460 ;
        RECT 5.085 -106.000 5.255 -105.460 ;
        RECT 5.575 -106.240 5.745 -105.460 ;
        RECT 6.640 -106.030 6.945 -105.285 ;
        RECT 7.640 -106.030 7.810 -104.310 ;
        RECT 8.620 -106.030 8.790 -104.310 ;
        RECT 6.640 -106.180 8.790 -106.030 ;
        RECT 9.740 -106.065 9.920 -102.315 ;
        RECT 6.695 -106.220 8.790 -106.180 ;
        RECT 9.030 -106.105 9.920 -106.065 ;
        RECT -1.650 -106.510 3.130 -106.340 ;
        RECT -1.650 -106.545 -0.975 -106.510 ;
        RECT 3.370 -106.670 6.445 -106.240 ;
        RECT 9.030 -106.285 9.965 -106.105 ;
        RECT 9.030 -106.305 9.855 -106.285 ;
        RECT 9.030 -106.335 9.705 -106.305 ;
        RECT 7.010 -106.585 7.380 -106.455 ;
        RECT 10.145 -106.575 10.345 -101.895 ;
        RECT 11.640 -105.175 11.810 -104.315 ;
        RECT 12.620 -104.855 12.790 -104.315 ;
        RECT 13.600 -104.855 13.770 -104.315 ;
        RECT 9.435 -106.585 10.345 -106.575 ;
        RECT -2.985 -106.960 -1.820 -106.790 ;
        RECT -0.955 -106.960 1.260 -106.790 ;
        RECT -4.560 -109.760 -4.390 -107.780 ;
        RECT -2.985 -108.820 -2.815 -106.960 ;
        RECT -2.495 -109.310 -2.325 -107.280 ;
        RECT -2.005 -108.820 -1.835 -106.960 ;
        RECT -0.955 -106.965 0.280 -106.960 ;
        RECT -0.955 -107.280 -0.780 -106.965 ;
        RECT -1.440 -108.765 -1.270 -107.280 ;
        RECT -1.445 -109.295 -1.270 -108.765 ;
        RECT -0.950 -108.820 -0.780 -107.280 ;
        RECT -0.460 -108.775 -0.290 -107.280 ;
        RECT -0.465 -109.295 -0.290 -108.775 ;
        RECT 0.110 -108.815 0.280 -106.965 ;
        RECT -1.445 -109.310 -0.290 -109.295 ;
        RECT -2.495 -109.480 -0.290 -109.310 ;
        RECT 0.600 -109.760 0.770 -107.275 ;
        RECT 1.090 -108.815 1.260 -106.960 ;
        RECT 4.920 -108.705 5.225 -106.670 ;
        RECT 7.010 -106.775 10.345 -106.585 ;
        RECT 10.820 -105.525 11.810 -105.175 ;
        RECT 13.995 -105.090 14.360 -105.025 ;
        RECT 13.995 -105.230 14.860 -105.090 ;
        RECT 13.995 -105.295 14.970 -105.230 ;
        RECT 13.995 -105.325 14.360 -105.295 ;
        RECT 7.010 -106.780 9.440 -106.775 ;
        RECT 7.010 -106.810 7.380 -106.780 ;
        RECT 9.085 -106.785 9.440 -106.780 ;
        RECT 7.150 -108.535 7.320 -106.995 ;
        RECT 7.640 -108.535 7.810 -106.995 ;
        RECT 8.130 -108.535 8.300 -106.995 ;
        RECT 8.620 -108.535 8.790 -106.995 ;
        RECT 9.110 -108.535 9.280 -106.995 ;
        RECT 4.920 -108.795 7.170 -108.705 ;
        RECT 8.620 -108.795 8.795 -108.535 ;
        RECT 4.920 -109.010 9.380 -108.795 ;
        RECT -5.110 -110.085 1.260 -109.760 ;
        RECT -5.045 -111.410 -4.395 -110.085 ;
        RECT -3.515 -111.410 -2.865 -110.085 ;
        RECT -1.930 -111.410 -1.280 -110.085 ;
        RECT 0.300 -111.410 0.950 -110.085 ;
        RECT 4.920 -111.410 5.675 -109.010 ;
        RECT 6.805 -109.100 9.380 -109.010 ;
        RECT 6.805 -111.410 7.425 -109.100 ;
        RECT 8.455 -111.410 9.075 -109.100 ;
        RECT 10.820 -109.200 11.170 -105.525 ;
        RECT 12.130 -106.010 12.300 -105.470 ;
        RECT 12.620 -106.250 12.790 -105.470 ;
        RECT 13.110 -106.010 13.280 -105.470 ;
        RECT 13.600 -106.250 13.770 -105.470 ;
        RECT 14.665 -106.040 14.970 -105.295 ;
        RECT 15.665 -106.040 15.835 -104.320 ;
        RECT 16.645 -106.040 16.815 -104.320 ;
        RECT 14.665 -106.190 16.815 -106.040 ;
        RECT 14.720 -106.230 16.815 -106.190 ;
        RECT 17.055 -106.105 17.730 -106.075 ;
        RECT 17.910 -106.105 18.090 -99.470 ;
        RECT 11.395 -106.680 14.470 -106.250 ;
        RECT 17.055 -106.295 18.090 -106.105 ;
        RECT 17.055 -106.305 17.990 -106.295 ;
        RECT 17.055 -106.345 17.730 -106.305 ;
        RECT 15.035 -106.595 15.405 -106.465 ;
        RECT 18.285 -106.585 18.485 -99.120 ;
        RECT 17.460 -106.595 18.485 -106.585 ;
        RECT 10.490 -109.430 11.170 -109.200 ;
        RECT 12.945 -108.715 13.250 -106.680 ;
        RECT 15.035 -106.785 18.485 -106.595 ;
        RECT 15.035 -106.790 17.465 -106.785 ;
        RECT 15.035 -106.820 15.405 -106.790 ;
        RECT 17.110 -106.795 17.465 -106.790 ;
        RECT 15.175 -108.545 15.345 -107.005 ;
        RECT 15.665 -108.545 15.835 -107.005 ;
        RECT 16.155 -108.545 16.325 -107.005 ;
        RECT 16.645 -108.545 16.815 -107.005 ;
        RECT 17.135 -108.545 17.305 -107.005 ;
        RECT 19.760 -107.195 19.930 -104.195 ;
        RECT 23.450 -105.415 23.620 -104.195 ;
        RECT 24.430 -105.415 24.600 -104.195 ;
        RECT 25.410 -105.415 25.580 -104.195 ;
        RECT 22.805 -105.600 25.580 -105.415 ;
        RECT 25.780 -105.470 26.455 -105.430 ;
        RECT 20.105 -106.290 20.780 -106.240 ;
        RECT 22.805 -106.290 22.990 -105.600 ;
        RECT 25.775 -105.655 26.550 -105.470 ;
        RECT 25.775 -105.700 26.455 -105.655 ;
        RECT 24.100 -105.885 24.775 -105.840 ;
        RECT 26.735 -105.885 26.905 -99.040 ;
        RECT 24.100 -106.075 26.905 -105.885 ;
        RECT 24.100 -106.110 24.775 -106.075 ;
        RECT 20.105 -106.475 22.990 -106.290 ;
        RECT 20.105 -106.510 20.780 -106.475 ;
        RECT 22.805 -106.745 22.990 -106.475 ;
        RECT 23.160 -106.295 23.835 -106.230 ;
        RECT 27.085 -106.295 27.255 -98.580 ;
        RECT 27.825 -103.730 31.465 -103.560 ;
        RECT 27.825 -105.290 27.995 -103.730 ;
        RECT 28.315 -105.470 28.485 -104.250 ;
        RECT 28.805 -105.290 28.975 -103.730 ;
        RECT 29.405 -104.075 31.115 -103.905 ;
        RECT 29.405 -105.290 29.575 -104.075 ;
        RECT 29.895 -105.470 30.065 -104.250 ;
        RECT 30.385 -105.290 30.555 -104.075 ;
        RECT 27.570 -105.640 30.640 -105.470 ;
        RECT 23.160 -106.465 27.255 -106.295 ;
        RECT 27.820 -106.310 28.515 -106.040 ;
        RECT 30.470 -106.215 30.640 -105.640 ;
        RECT 30.945 -105.835 31.115 -104.075 ;
        RECT 31.295 -105.465 31.465 -103.730 ;
        RECT 32.195 -105.465 32.365 -104.250 ;
        RECT 31.295 -105.635 32.365 -105.465 ;
        RECT 33.175 -105.835 33.345 -104.250 ;
        RECT 34.725 -105.215 34.895 -104.250 ;
        RECT 36.270 -105.205 36.440 -104.250 ;
        RECT 30.945 -106.005 33.345 -105.835 ;
        RECT 33.610 -106.090 34.305 -105.820 ;
        RECT 30.470 -106.385 31.200 -106.215 ;
        RECT 23.160 -106.500 23.835 -106.465 ;
        RECT 31.030 -106.695 31.200 -106.385 ;
        RECT 31.565 -106.460 32.260 -106.190 ;
        RECT 18.680 -107.485 19.930 -107.195 ;
        RECT 12.945 -108.805 15.195 -108.715 ;
        RECT 16.645 -108.805 16.820 -108.545 ;
        RECT 12.945 -109.020 17.405 -108.805 ;
        RECT 12.945 -111.410 13.700 -109.020 ;
        RECT 15.155 -109.110 17.405 -109.020 ;
        RECT 15.155 -111.410 15.910 -109.110 ;
        RECT 16.620 -111.410 17.375 -109.110 ;
        RECT 18.680 -109.760 19.005 -107.485 ;
        RECT 19.760 -108.775 19.930 -107.485 ;
        RECT 21.825 -106.915 22.990 -106.745 ;
        RECT 23.855 -106.915 26.070 -106.745 ;
        RECT 20.250 -109.715 20.420 -107.735 ;
        RECT 21.825 -108.775 21.995 -106.915 ;
        RECT 22.315 -109.265 22.485 -107.235 ;
        RECT 22.805 -108.775 22.975 -106.915 ;
        RECT 23.855 -106.920 25.090 -106.915 ;
        RECT 23.855 -107.235 24.030 -106.920 ;
        RECT 23.370 -108.720 23.540 -107.235 ;
        RECT 23.365 -109.250 23.540 -108.720 ;
        RECT 23.860 -108.775 24.030 -107.235 ;
        RECT 24.350 -108.730 24.520 -107.235 ;
        RECT 24.345 -109.250 24.520 -108.730 ;
        RECT 24.920 -108.770 25.090 -106.920 ;
        RECT 23.365 -109.265 24.520 -109.250 ;
        RECT 22.315 -109.435 24.520 -109.265 ;
        RECT 25.410 -109.715 25.580 -107.230 ;
        RECT 25.900 -108.770 26.070 -106.915 ;
        RECT 27.815 -106.900 29.470 -106.715 ;
        RECT 31.030 -106.865 33.835 -106.695 ;
        RECT 27.815 -107.315 28.000 -106.900 ;
        RECT 29.285 -107.020 29.470 -106.900 ;
        RECT 29.285 -107.205 30.065 -107.020 ;
        RECT 27.825 -108.260 27.995 -107.315 ;
        RECT 27.805 -108.875 28.000 -108.260 ;
        RECT 28.315 -108.505 28.485 -107.280 ;
        RECT 29.880 -107.310 30.065 -107.205 ;
        RECT 29.895 -108.320 30.065 -107.310 ;
        RECT 30.375 -107.325 31.875 -107.130 ;
        RECT 30.385 -108.320 30.555 -107.325 ;
        RECT 31.705 -108.320 31.875 -107.325 ;
        RECT 32.195 -108.320 32.365 -106.865 ;
        RECT 33.175 -108.235 33.345 -107.280 ;
        RECT 33.175 -108.505 33.355 -108.235 ;
        RECT 33.665 -108.320 33.835 -106.865 ;
        RECT 34.700 -106.910 34.915 -105.215 ;
        RECT 36.250 -106.190 36.465 -105.205 ;
        RECT 36.685 -106.120 37.380 -105.850 ;
        RECT 35.750 -106.420 36.465 -106.190 ;
        RECT 34.220 -107.140 34.915 -106.910 ;
        RECT 34.700 -107.365 34.915 -107.140 ;
        RECT 34.725 -108.320 34.895 -107.365 ;
        RECT 35.215 -108.285 35.385 -107.280 ;
        RECT 36.250 -107.375 36.465 -106.420 ;
        RECT 28.315 -108.685 33.355 -108.505 ;
        RECT 35.190 -108.705 35.405 -108.285 ;
        RECT 36.270 -108.320 36.440 -107.375 ;
        RECT 36.760 -108.275 36.930 -107.280 ;
        RECT 36.735 -108.705 36.950 -108.275 ;
        RECT 33.810 -108.875 36.970 -108.705 ;
        RECT 27.805 -109.140 36.970 -108.875 ;
        RECT 18.330 -109.990 19.010 -109.760 ;
        RECT 19.700 -110.040 26.070 -109.715 ;
        RECT 19.820 -111.410 20.550 -110.040 ;
        RECT 22.045 -111.410 22.775 -110.040 ;
        RECT 23.375 -111.410 24.105 -110.040 ;
        RECT 25.175 -111.410 25.905 -110.040 ;
        RECT 27.995 -111.410 28.980 -109.140 ;
        RECT 30.660 -111.410 31.645 -109.140 ;
        RECT 33.225 -109.185 36.970 -109.140 ;
        RECT 33.225 -111.410 34.210 -109.185 ;
        RECT 35.740 -111.410 36.725 -109.185 ;
        RECT 37.715 -111.410 39.020 -97.995 ;
        RECT 41.200 -98.250 77.530 -97.555 ;
        RECT 76.335 -100.570 77.510 -100.455 ;
        RECT 49.295 -101.795 77.510 -100.570 ;
        RECT 49.295 -101.805 76.890 -101.795 ;
        RECT 75.905 -102.650 77.240 -102.470 ;
        RECT 49.180 -103.825 77.240 -102.650 ;
        RECT 75.905 -103.960 77.240 -103.825 ;
        RECT 41.340 -105.620 42.430 -105.580 ;
        RECT 77.220 -105.620 77.985 -105.425 ;
        RECT 41.340 -105.995 77.985 -105.620 ;
        RECT 41.340 -106.025 42.430 -105.995 ;
        RECT 77.220 -106.180 77.985 -105.995 ;
        RECT 46.250 -106.725 46.500 -106.695 ;
        RECT 73.810 -106.725 74.300 -106.655 ;
        RECT 46.205 -107.340 74.300 -106.725 ;
        RECT 46.250 -107.360 46.500 -107.340 ;
        RECT 73.810 -107.475 74.300 -107.340 ;
        RECT 78.395 -108.750 79.035 -94.190 ;
        RECT 79.660 -108.305 80.320 -92.050 ;
        RECT 80.870 -105.425 81.315 -89.675 ;
        RECT 91.330 -95.745 94.055 -88.055 ;
        RECT 88.415 -98.275 418.280 -95.745 ;
        RECT 85.190 -101.470 86.280 -100.240 ;
        RECT 80.870 -106.180 81.355 -105.425 ;
        RECT 85.385 -105.755 86.095 -101.470 ;
        RECT 91.330 -105.595 94.055 -98.275 ;
        RECT 126.395 -100.770 128.045 -100.355 ;
        RECT 140.060 -100.580 141.475 -98.275 ;
        RECT 138.840 -100.720 142.165 -100.580 ;
        RECT 166.900 -100.655 168.685 -100.320 ;
        RECT 172.790 -100.655 174.575 -100.490 ;
        RECT 182.055 -100.635 183.470 -98.275 ;
        RECT 126.395 -101.665 132.290 -100.770 ;
        RECT 138.840 -101.010 144.015 -100.720 ;
        RECT 138.840 -101.415 139.270 -101.010 ;
        RECT 140.140 -101.195 140.315 -101.010 ;
        RECT 141.765 -101.025 144.015 -101.010 ;
        RECT 126.395 -101.825 128.045 -101.665 ;
        RECT 134.580 -101.845 139.270 -101.415 ;
        RECT 133.820 -103.295 134.470 -102.835 ;
        RECT 135.280 -103.125 135.450 -101.845 ;
        RECT 135.770 -103.125 135.940 -102.085 ;
        RECT 136.260 -103.125 136.430 -101.845 ;
        RECT 136.750 -102.955 136.920 -102.085 ;
        RECT 139.655 -102.735 139.825 -101.195 ;
        RECT 140.145 -102.735 140.315 -101.195 ;
        RECT 140.635 -102.735 140.805 -101.195 ;
        RECT 141.125 -102.735 141.295 -101.195 ;
        RECT 141.615 -102.735 141.785 -101.195 ;
        RECT 139.495 -102.950 139.850 -102.945 ;
        RECT 141.555 -102.950 141.925 -102.920 ;
        RECT 139.495 -102.955 141.925 -102.950 ;
        RECT 136.750 -103.125 141.925 -102.955 ;
        RECT 143.710 -103.060 144.015 -101.025 ;
        RECT 166.900 -101.600 174.575 -100.655 ;
        RECT 181.040 -100.775 184.365 -100.635 ;
        RECT 181.040 -101.065 186.215 -100.775 ;
        RECT 226.615 -100.830 228.030 -98.275 ;
        RECT 272.710 -100.660 274.125 -98.275 ;
        RECT 299.455 -100.500 301.335 -100.025 ;
        RECT 316.685 -100.330 318.220 -98.275 ;
        RECT 307.460 -100.500 308.710 -100.365 ;
        RECT 181.040 -101.470 181.470 -101.065 ;
        RECT 182.340 -101.250 182.515 -101.065 ;
        RECT 183.965 -101.080 186.215 -101.065 ;
        RECT 166.900 -101.655 168.685 -101.600 ;
        RECT 172.790 -101.825 174.575 -101.600 ;
        RECT 176.780 -101.900 181.470 -101.470 ;
        RECT 136.755 -103.145 141.925 -103.125 ;
        RECT 136.755 -103.155 139.500 -103.145 ;
        RECT 134.690 -103.295 135.055 -103.265 ;
        RECT 141.555 -103.275 141.925 -103.145 ;
        RECT 133.820 -103.500 135.055 -103.295 ;
        RECT 139.230 -103.435 139.905 -103.395 ;
        RECT 139.130 -103.445 139.905 -103.435 ;
        RECT 133.820 -103.585 134.470 -103.500 ;
        RECT 134.690 -103.565 135.055 -103.500 ;
        RECT 138.095 -103.625 139.905 -103.445 ;
        RECT 142.490 -103.490 146.415 -103.060 ;
        RECT 176.020 -103.350 176.670 -102.890 ;
        RECT 177.480 -103.180 177.650 -101.900 ;
        RECT 177.970 -103.180 178.140 -102.140 ;
        RECT 178.460 -103.180 178.630 -101.900 ;
        RECT 178.950 -103.010 179.120 -102.140 ;
        RECT 181.855 -102.790 182.025 -101.250 ;
        RECT 182.345 -102.790 182.515 -101.250 ;
        RECT 182.835 -102.790 183.005 -101.250 ;
        RECT 183.325 -102.790 183.495 -101.250 ;
        RECT 183.815 -102.790 183.985 -101.250 ;
        RECT 181.695 -103.005 182.050 -103.000 ;
        RECT 183.755 -103.005 184.125 -102.975 ;
        RECT 181.695 -103.010 184.125 -103.005 ;
        RECT 178.950 -103.180 184.125 -103.010 ;
        RECT 185.910 -103.115 186.215 -101.080 ;
        RECT 209.680 -101.100 211.005 -100.945 ;
        RECT 217.310 -101.100 218.795 -100.935 ;
        RECT 209.680 -101.935 218.795 -101.100 ;
        RECT 225.355 -100.970 228.680 -100.830 ;
        RECT 225.355 -101.260 230.530 -100.970 ;
        RECT 225.355 -101.665 225.785 -101.260 ;
        RECT 226.655 -101.445 226.830 -101.260 ;
        RECT 228.280 -101.275 230.530 -101.260 ;
        RECT 209.680 -102.270 211.005 -101.935 ;
        RECT 217.310 -102.045 218.795 -101.935 ;
        RECT 221.095 -102.095 225.785 -101.665 ;
        RECT 178.955 -103.200 184.125 -103.180 ;
        RECT 178.955 -103.210 181.700 -103.200 ;
        RECT 176.890 -103.350 177.255 -103.320 ;
        RECT 183.755 -103.330 184.125 -103.200 ;
        RECT 139.130 -103.635 139.905 -103.625 ;
        RECT 139.230 -103.665 139.905 -103.635 ;
        RECT 140.145 -103.550 142.240 -103.510 ;
        RECT 140.145 -103.700 142.295 -103.550 ;
        RECT 135.280 -104.775 135.450 -103.735 ;
        RECT 136.260 -104.775 136.430 -103.735 ;
        RECT 137.240 -104.775 137.410 -103.735 ;
        RECT 98.380 -105.405 101.520 -105.235 ;
        RECT 80.870 -107.845 81.315 -106.180 ;
        RECT 85.200 -106.700 86.095 -105.755 ;
        RECT 86.840 -106.125 95.690 -105.595 ;
        RECT 97.915 -106.075 98.085 -105.575 ;
        RECT 98.380 -105.660 98.590 -105.405 ;
        RECT 87.360 -106.855 87.600 -106.125 ;
        RECT 87.385 -107.710 87.555 -106.855 ;
        RECT 87.875 -107.625 88.045 -106.670 ;
        RECT 88.330 -106.870 88.570 -106.125 ;
        RECT 86.455 -107.845 87.180 -107.810 ;
        RECT 80.870 -108.050 87.180 -107.845 ;
        RECT 86.455 -108.090 87.180 -108.050 ;
        RECT 87.855 -107.880 88.065 -107.625 ;
        RECT 88.365 -107.710 88.535 -106.870 ;
        RECT 88.855 -107.625 89.025 -106.670 ;
        RECT 88.835 -107.880 89.045 -107.625 ;
        RECT 87.855 -108.090 91.785 -107.880 ;
        RECT 91.090 -108.180 91.785 -108.090 ;
        RECT 88.100 -108.305 88.825 -108.285 ;
        RECT 79.660 -108.510 88.825 -108.305 ;
        RECT 88.100 -108.565 88.825 -108.510 ;
        RECT 89.700 -108.725 90.425 -108.445 ;
        RECT 89.700 -108.750 90.000 -108.725 ;
        RECT 78.395 -108.955 90.000 -108.750 ;
        RECT 91.090 -109.090 91.300 -108.180 ;
        RECT 87.365 -109.320 89.610 -109.135 ;
        RECT 87.365 -109.575 87.570 -109.320 ;
        RECT 88.420 -109.540 88.630 -109.320 ;
        RECT -15.100 -112.050 -11.960 -111.880 ;
        RECT -66.100 -112.685 -65.325 -112.675 ;
        RECT -66.000 -112.725 -65.325 -112.685 ;
        RECT -68.475 -112.975 -65.730 -112.965 ;
        RECT -63.675 -112.975 -63.305 -112.845 ;
        RECT -68.475 -112.995 -63.305 -112.975 ;
        RECT -80.775 -113.705 -79.735 -113.695 ;
        RECT -128.320 -114.995 -125.195 -113.895 ;
        RECT -69.950 -114.275 -69.780 -112.995 ;
        RECT -69.460 -114.035 -69.290 -112.995 ;
        RECT -68.970 -114.275 -68.800 -112.995 ;
        RECT -68.480 -113.165 -63.305 -112.995 ;
        RECT -62.740 -113.060 -58.815 -112.630 ;
        RECT -10.275 -112.715 39.020 -111.410 ;
        RECT 87.385 -112.530 87.555 -109.575 ;
        RECT 88.445 -112.530 88.615 -109.540 ;
        RECT 88.935 -112.500 89.105 -109.490 ;
        RECT 89.400 -109.545 89.610 -109.320 ;
        RECT 90.460 -109.300 91.300 -109.090 ;
        RECT -68.480 -114.035 -68.310 -113.165 ;
        RECT -65.735 -113.170 -63.305 -113.165 ;
        RECT -65.735 -113.175 -65.380 -113.170 ;
        RECT -63.675 -113.200 -63.305 -113.170 ;
        RECT -70.650 -114.705 -65.960 -114.275 ;
        RECT -85.470 -114.995 -84.130 -114.760 ;
        RECT -128.320 -115.925 -84.130 -114.995 ;
        RECT -66.390 -115.110 -65.960 -114.705 ;
        RECT -65.575 -114.925 -65.405 -113.385 ;
        RECT -65.085 -114.925 -64.915 -113.385 ;
        RECT -64.595 -114.925 -64.425 -113.385 ;
        RECT -64.105 -114.925 -63.935 -113.385 ;
        RECT -63.615 -114.925 -63.445 -113.385 ;
        RECT -65.090 -115.110 -64.915 -114.925 ;
        RECT -61.520 -115.095 -61.215 -113.060 ;
        RECT -63.465 -115.110 -61.215 -115.095 ;
        RECT -66.390 -115.400 -61.215 -115.110 ;
        RECT -66.390 -115.540 -63.065 -115.400 ;
        RECT -128.320 -117.020 -125.195 -115.925 ;
        RECT -85.470 -116.085 -84.130 -115.925 ;
        RECT -67.970 -116.505 -64.830 -116.335 ;
        RECT -75.205 -116.620 -75.035 -116.600 ;
        RECT -75.235 -117.885 -75.005 -116.620 ;
        RECT -74.225 -117.560 -74.055 -116.600 ;
        RECT -73.245 -117.560 -73.075 -116.600 ;
        RECT -71.020 -116.620 -70.850 -116.600 ;
        RECT -72.125 -117.030 -71.840 -116.710 ;
        RECT -72.840 -117.275 -71.840 -117.030 ;
        RECT -74.255 -117.885 -74.025 -117.560 ;
        RECT -73.275 -117.885 -73.045 -117.560 ;
        RECT -75.235 -117.925 -73.045 -117.885 ;
        RECT -72.840 -117.925 -72.610 -117.275 ;
        RECT -72.125 -117.530 -71.840 -117.275 ;
        RECT -76.255 -118.110 -75.415 -117.960 ;
        RECT -76.290 -118.330 -75.415 -118.110 ;
        RECT -75.235 -118.115 -72.610 -117.925 ;
        RECT -71.050 -117.885 -70.820 -116.620 ;
        RECT -70.040 -117.560 -69.870 -116.600 ;
        RECT -69.060 -117.560 -68.890 -116.600 ;
        RECT -67.970 -116.730 -67.790 -116.505 ;
        RECT -70.070 -117.885 -69.840 -117.560 ;
        RECT -69.090 -117.885 -68.860 -117.560 ;
        RECT -71.050 -117.925 -68.860 -117.885 ;
        RECT -68.585 -117.805 -68.215 -116.965 ;
        RECT -67.965 -117.100 -67.795 -116.730 ;
        RECT -68.585 -117.925 -68.220 -117.805 ;
        RECT -72.070 -118.015 -71.230 -117.960 ;
        RECT -72.245 -118.020 -71.230 -118.015 ;
        RECT -76.290 -120.190 -76.050 -118.330 ;
        RECT -75.695 -119.295 -75.525 -118.500 ;
        RECT -75.235 -118.580 -75.005 -118.115 ;
        RECT -75.205 -119.040 -75.035 -118.580 ;
        RECT -74.715 -119.295 -74.545 -118.500 ;
        RECT -74.255 -118.580 -74.025 -118.115 ;
        RECT -73.275 -118.275 -72.610 -118.115 ;
        RECT -74.225 -119.040 -74.055 -118.580 ;
        RECT -73.735 -119.295 -73.565 -118.500 ;
        RECT -73.275 -118.580 -73.045 -118.275 ;
        RECT -72.430 -118.330 -71.230 -118.020 ;
        RECT -71.050 -118.115 -68.220 -117.925 ;
        RECT -73.245 -119.040 -73.075 -118.580 ;
        RECT -72.430 -119.050 -72.130 -118.330 ;
        RECT -71.510 -119.295 -71.340 -118.500 ;
        RECT -71.050 -118.580 -70.820 -118.115 ;
        RECT -71.020 -119.040 -70.850 -118.580 ;
        RECT -70.530 -119.295 -70.360 -118.500 ;
        RECT -70.070 -118.580 -69.840 -118.115 ;
        RECT -69.090 -118.275 -68.220 -118.115 ;
        RECT -67.995 -117.835 -67.760 -117.100 ;
        RECT -67.475 -117.135 -67.305 -116.675 ;
        RECT -66.990 -116.780 -66.780 -116.505 ;
        RECT -67.480 -117.395 -67.300 -117.135 ;
        RECT -66.985 -117.215 -66.815 -116.780 ;
        RECT -66.495 -117.125 -66.325 -116.675 ;
        RECT -66.020 -116.785 -65.810 -116.505 ;
        RECT -66.495 -117.215 -66.310 -117.125 ;
        RECT -66.005 -117.215 -65.835 -116.785 ;
        RECT -65.515 -117.125 -65.345 -116.675 ;
        RECT -65.040 -116.760 -64.830 -116.505 ;
        RECT -54.470 -116.505 -51.330 -116.335 ;
        RECT -61.705 -116.620 -61.535 -116.600 ;
        RECT -66.490 -117.395 -66.310 -117.215 ;
        RECT -65.520 -117.395 -65.340 -117.125 ;
        RECT -65.025 -117.215 -64.855 -116.760 ;
        RECT -64.535 -117.175 -64.365 -116.675 ;
        RECT -64.550 -117.395 -64.340 -117.175 ;
        RECT -67.480 -117.565 -64.340 -117.395 ;
        RECT -67.995 -118.205 -67.135 -117.835 ;
        RECT -65.215 -118.100 -64.340 -117.565 ;
        RECT -61.735 -117.885 -61.505 -116.620 ;
        RECT -60.725 -117.560 -60.555 -116.600 ;
        RECT -59.745 -117.560 -59.575 -116.600 ;
        RECT -57.520 -116.620 -57.350 -116.600 ;
        RECT -58.625 -116.970 -58.340 -116.710 ;
        RECT -59.365 -117.280 -58.340 -116.970 ;
        RECT -60.755 -117.885 -60.525 -117.560 ;
        RECT -59.775 -117.885 -59.545 -117.560 ;
        RECT -61.735 -117.925 -59.545 -117.885 ;
        RECT -59.365 -117.925 -59.055 -117.280 ;
        RECT -58.625 -117.530 -58.340 -117.280 ;
        RECT -62.755 -117.995 -61.915 -117.960 ;
        RECT -70.040 -119.040 -69.870 -118.580 ;
        RECT -69.550 -119.295 -69.380 -118.500 ;
        RECT -69.090 -118.580 -68.860 -118.275 ;
        RECT -69.060 -119.040 -68.890 -118.580 ;
        RECT -67.995 -118.880 -67.760 -118.205 ;
        RECT -65.215 -118.400 -63.885 -118.100 ;
        RECT -62.865 -118.295 -61.915 -117.995 ;
        RECT -62.755 -118.330 -61.915 -118.295 ;
        RECT -61.735 -118.115 -59.055 -117.925 ;
        RECT -57.550 -117.885 -57.320 -116.620 ;
        RECT -56.540 -117.560 -56.370 -116.600 ;
        RECT -55.560 -117.560 -55.390 -116.600 ;
        RECT -54.470 -116.730 -54.290 -116.505 ;
        RECT -56.570 -117.885 -56.340 -117.560 ;
        RECT -55.590 -117.885 -55.360 -117.560 ;
        RECT -57.550 -117.925 -55.360 -117.885 ;
        RECT -55.085 -117.805 -54.715 -116.965 ;
        RECT -54.465 -117.100 -54.295 -116.730 ;
        RECT -55.085 -117.925 -54.720 -117.805 ;
        RECT -58.570 -118.015 -57.730 -117.960 ;
        RECT -67.495 -118.570 -64.340 -118.400 ;
        RECT -67.495 -118.775 -67.290 -118.570 ;
        RECT -67.965 -119.230 -67.795 -118.880 ;
        RECT -75.740 -119.635 -68.885 -119.295 ;
        RECT -67.990 -119.520 -67.770 -119.230 ;
        RECT -67.475 -119.290 -67.305 -118.775 ;
        RECT -66.985 -119.175 -66.815 -118.750 ;
        RECT -66.505 -118.815 -66.300 -118.570 ;
        RECT -67.010 -119.520 -66.790 -119.175 ;
        RECT -66.495 -119.290 -66.325 -118.815 ;
        RECT -66.005 -119.175 -65.835 -118.750 ;
        RECT -65.535 -118.815 -65.330 -118.570 ;
        RECT -64.550 -118.605 -64.340 -118.570 ;
        RECT -66.030 -119.520 -65.810 -119.175 ;
        RECT -65.515 -119.290 -65.345 -118.815 ;
        RECT -65.025 -119.230 -64.855 -118.750 ;
        RECT -64.550 -118.820 -64.345 -118.605 ;
        RECT -65.045 -119.520 -64.825 -119.230 ;
        RECT -64.535 -119.290 -64.365 -118.820 ;
        RECT -62.195 -119.295 -62.025 -118.500 ;
        RECT -61.735 -118.580 -61.505 -118.115 ;
        RECT -61.705 -119.040 -61.535 -118.580 ;
        RECT -61.215 -119.295 -61.045 -118.500 ;
        RECT -60.755 -118.580 -60.525 -118.115 ;
        RECT -59.775 -118.275 -59.055 -118.115 ;
        RECT -60.725 -119.040 -60.555 -118.580 ;
        RECT -60.235 -119.295 -60.065 -118.500 ;
        RECT -59.775 -118.580 -59.545 -118.275 ;
        RECT -58.870 -118.330 -57.730 -118.015 ;
        RECT -57.550 -118.115 -54.720 -117.925 ;
        RECT -59.745 -119.040 -59.575 -118.580 ;
        RECT -58.870 -119.125 -58.570 -118.330 ;
        RECT -58.010 -119.295 -57.840 -118.500 ;
        RECT -57.550 -118.580 -57.320 -118.115 ;
        RECT -57.520 -119.040 -57.350 -118.580 ;
        RECT -57.030 -119.295 -56.860 -118.500 ;
        RECT -56.570 -118.580 -56.340 -118.115 ;
        RECT -55.590 -118.275 -54.720 -118.115 ;
        RECT -54.495 -117.835 -54.260 -117.100 ;
        RECT -53.975 -117.135 -53.805 -116.675 ;
        RECT -53.490 -116.780 -53.280 -116.505 ;
        RECT -53.980 -117.395 -53.800 -117.135 ;
        RECT -53.485 -117.215 -53.315 -116.780 ;
        RECT -52.995 -117.125 -52.825 -116.675 ;
        RECT -52.520 -116.785 -52.310 -116.505 ;
        RECT -52.995 -117.215 -52.810 -117.125 ;
        RECT -52.505 -117.215 -52.335 -116.785 ;
        RECT -52.015 -117.125 -51.845 -116.675 ;
        RECT -51.540 -116.760 -51.330 -116.505 ;
        RECT -43.210 -116.515 -42.010 -116.345 ;
        RECT -52.990 -117.395 -52.810 -117.215 ;
        RECT -52.020 -117.395 -51.840 -117.125 ;
        RECT -51.525 -117.215 -51.355 -116.760 ;
        RECT -51.035 -117.175 -50.865 -116.675 ;
        RECT -51.050 -117.395 -50.840 -117.175 ;
        RECT -53.980 -117.565 -50.840 -117.395 ;
        RECT -54.495 -118.205 -53.635 -117.835 ;
        RECT -51.715 -118.110 -50.840 -117.565 ;
        RECT -56.540 -119.040 -56.370 -118.580 ;
        RECT -56.050 -119.295 -55.880 -118.500 ;
        RECT -55.590 -118.580 -55.360 -118.275 ;
        RECT -55.560 -119.040 -55.390 -118.580 ;
        RECT -54.495 -118.880 -54.260 -118.205 ;
        RECT -51.715 -118.400 -50.465 -118.110 ;
        RECT -53.995 -118.410 -50.465 -118.400 ;
        RECT -53.995 -118.570 -50.840 -118.410 ;
        RECT -53.995 -118.775 -53.790 -118.570 ;
        RECT -54.465 -119.230 -54.295 -118.880 ;
        RECT -74.500 -119.835 -73.945 -119.635 ;
        RECT -74.555 -119.875 -73.870 -119.835 ;
        RECT -70.445 -119.875 -69.890 -119.635 ;
        RECT -67.990 -119.690 -64.825 -119.520 ;
        RECT -62.240 -119.305 -59.570 -119.295 ;
        RECT -58.055 -119.305 -55.385 -119.295 ;
        RECT -62.240 -119.635 -55.385 -119.305 ;
        RECT -54.490 -119.520 -54.270 -119.230 ;
        RECT -53.975 -119.290 -53.805 -118.775 ;
        RECT -53.485 -119.175 -53.315 -118.750 ;
        RECT -53.005 -118.815 -52.800 -118.570 ;
        RECT -53.510 -119.520 -53.290 -119.175 ;
        RECT -52.995 -119.290 -52.825 -118.815 ;
        RECT -52.505 -119.175 -52.335 -118.750 ;
        RECT -52.035 -118.815 -51.830 -118.570 ;
        RECT -51.050 -118.605 -50.840 -118.570 ;
        RECT -52.530 -119.520 -52.310 -119.175 ;
        RECT -52.015 -119.290 -51.845 -118.815 ;
        RECT -51.525 -119.230 -51.355 -118.750 ;
        RECT -51.050 -118.820 -50.845 -118.605 ;
        RECT -51.545 -119.520 -51.325 -119.230 ;
        RECT -51.035 -119.290 -50.865 -118.820 ;
        RECT -61.455 -119.865 -60.900 -119.635 ;
        RECT -60.540 -119.645 -57.940 -119.635 ;
        RECT -61.570 -119.875 -60.885 -119.865 ;
        RECT -57.065 -119.875 -56.510 -119.635 ;
        RECT -54.490 -119.690 -51.325 -119.520 ;
        RECT -44.240 -119.655 -44.070 -116.685 ;
        RECT -43.210 -116.735 -43.000 -116.515 ;
        RECT -48.380 -119.875 -47.720 -119.865 ;
        RECT -74.640 -120.070 -47.715 -119.875 ;
        RECT -74.555 -120.135 -73.870 -120.070 ;
        RECT -61.570 -120.165 -60.885 -120.070 ;
        RECT -48.380 -120.165 -47.720 -120.070 ;
        RECT -76.295 -120.875 -75.995 -120.190 ;
        RECT -63.745 -120.335 -63.060 -120.280 ;
        RECT -59.015 -120.335 -58.355 -120.285 ;
        RECT -74.640 -120.530 -45.990 -120.335 ;
        RECT -63.745 -120.580 -63.060 -120.530 ;
        RECT -59.015 -120.585 -58.355 -120.530 ;
        RECT -72.610 -120.765 -71.950 -120.725 ;
        RECT -49.995 -120.765 -49.335 -120.715 ;
        RECT -105.540 -121.490 -104.320 -121.300 ;
        RECT -111.090 -121.845 -108.775 -121.675 ;
        RECT -112.590 -124.980 -112.420 -122.025 ;
        RECT -112.610 -125.235 -112.405 -124.980 ;
        RECT -111.530 -125.015 -111.360 -122.025 ;
        RECT -111.090 -122.055 -110.825 -121.845 ;
        RECT -111.555 -125.235 -111.345 -125.015 ;
        RECT -111.040 -125.065 -110.870 -122.055 ;
        RECT -110.550 -125.010 -110.380 -122.025 ;
        RECT -110.045 -122.055 -109.765 -121.845 ;
        RECT -110.575 -125.235 -110.365 -125.010 ;
        RECT -109.985 -125.065 -109.815 -122.055 ;
        RECT -109.495 -124.975 -109.325 -122.025 ;
        RECT -109.055 -122.055 -108.775 -121.845 ;
        RECT -112.610 -125.420 -110.365 -125.235 ;
        RECT -109.515 -125.255 -109.305 -124.975 ;
        RECT -109.005 -125.065 -108.835 -122.055 ;
        RECT -106.560 -123.685 -106.390 -121.670 ;
        RECT -105.540 -121.810 -105.310 -121.490 ;
        RECT -106.565 -123.880 -106.385 -123.685 ;
        RECT -105.505 -123.710 -105.335 -121.810 ;
        RECT -105.015 -123.660 -104.845 -121.670 ;
        RECT -104.550 -121.810 -104.320 -121.490 ;
        RECT -101.015 -121.495 -99.795 -121.305 ;
        RECT -104.525 -123.480 -104.355 -121.810 ;
        RECT -105.050 -123.880 -104.825 -123.660 ;
        RECT -106.565 -124.060 -104.825 -123.880 ;
        RECT -104.540 -124.640 -104.290 -123.480 ;
        RECT -102.035 -123.690 -101.865 -121.675 ;
        RECT -101.015 -121.815 -100.785 -121.495 ;
        RECT -102.040 -123.885 -101.860 -123.690 ;
        RECT -100.980 -123.715 -100.810 -121.815 ;
        RECT -100.490 -123.665 -100.320 -121.675 ;
        RECT -100.025 -121.815 -99.795 -121.495 ;
        RECT -91.460 -121.685 -84.075 -121.120 ;
        RECT -100.000 -123.485 -99.830 -121.815 ;
        RECT -95.615 -123.160 -93.370 -123.070 ;
        RECT -91.460 -123.160 -91.155 -121.685 ;
        RECT -87.825 -122.275 -87.590 -121.685 ;
        RECT -98.175 -123.465 -91.155 -123.160 ;
        RECT -100.525 -123.885 -100.300 -123.665 ;
        RECT -102.040 -124.065 -100.300 -123.885 ;
        RECT -104.540 -124.705 -103.810 -124.640 ;
        RECT -104.820 -124.750 -103.810 -124.705 ;
        RECT -100.015 -124.645 -99.765 -123.485 ;
        RECT -100.015 -124.710 -99.155 -124.645 ;
        RECT -106.095 -124.930 -103.810 -124.750 ;
        RECT -100.295 -124.755 -99.155 -124.710 ;
        RECT -109.515 -125.465 -108.675 -125.255 ;
        RECT -108.885 -126.385 -108.675 -125.465 ;
        RECT -106.560 -125.925 -106.390 -125.130 ;
        RECT -106.095 -125.175 -105.870 -124.930 ;
        RECT -101.570 -124.935 -99.155 -124.755 ;
        RECT -108.930 -126.465 -108.245 -126.385 ;
        RECT -112.120 -126.675 -108.245 -126.465 ;
        RECT -112.590 -127.700 -112.420 -126.845 ;
        RECT -112.120 -126.930 -111.910 -126.675 ;
        RECT -112.615 -128.345 -112.375 -127.700 ;
        RECT -112.100 -127.885 -111.930 -126.930 ;
        RECT -111.610 -127.685 -111.440 -126.845 ;
        RECT -111.140 -126.930 -110.930 -126.675 ;
        RECT -106.580 -126.685 -106.360 -125.925 ;
        RECT -106.070 -126.170 -105.900 -125.175 ;
        RECT -105.580 -125.930 -105.410 -125.130 ;
        RECT -102.035 -125.930 -101.865 -125.135 ;
        RECT -101.570 -125.180 -101.345 -124.935 ;
        RECT -105.610 -126.685 -105.390 -125.930 ;
        RECT -107.225 -126.860 -104.240 -126.685 ;
        RECT -102.055 -126.690 -101.835 -125.930 ;
        RECT -101.545 -126.175 -101.375 -125.180 ;
        RECT -101.055 -125.935 -100.885 -125.135 ;
        RECT -98.175 -125.255 -97.870 -123.465 ;
        RECT -95.030 -123.635 -94.855 -123.465 ;
        RECT -95.515 -125.175 -95.345 -123.635 ;
        RECT -95.025 -125.175 -94.855 -123.635 ;
        RECT -94.535 -125.175 -94.365 -123.635 ;
        RECT -94.045 -125.175 -93.875 -123.635 ;
        RECT -93.555 -125.175 -93.385 -123.635 ;
        RECT -100.110 -125.560 -97.870 -125.255 ;
        RECT -95.675 -125.390 -95.320 -125.385 ;
        RECT -93.615 -125.390 -93.245 -125.360 ;
        RECT -95.675 -125.395 -93.245 -125.390 ;
        RECT -101.085 -126.690 -100.865 -125.935 ;
        RECT -100.110 -126.690 -99.805 -125.560 ;
        RECT -96.805 -125.585 -93.245 -125.395 ;
        RECT -91.460 -125.500 -91.155 -123.465 ;
        RECT -87.790 -123.745 -87.620 -122.275 ;
        RECT -87.300 -123.665 -87.130 -122.205 ;
        RECT -86.845 -122.280 -86.610 -121.685 ;
        RECT -88.335 -123.975 -87.560 -123.915 ;
        RECT -88.520 -124.145 -87.560 -123.975 ;
        RECT -88.335 -124.190 -87.560 -124.145 ;
        RECT -87.330 -124.015 -87.105 -123.665 ;
        RECT -86.810 -123.745 -86.640 -122.280 ;
        RECT -85.635 -122.330 -85.400 -121.685 ;
        RECT -85.600 -123.745 -85.430 -122.330 ;
        RECT -85.110 -123.700 -84.940 -122.205 ;
        RECT -76.290 -122.665 -76.050 -120.875 ;
        RECT -74.640 -120.960 -49.335 -120.765 ;
        RECT -72.610 -121.025 -71.950 -120.960 ;
        RECT -49.995 -121.015 -49.335 -120.960 ;
        RECT -46.185 -120.875 -45.990 -120.530 ;
        RECT -44.280 -120.875 -44.065 -119.655 ;
        RECT -43.180 -119.725 -43.010 -116.735 ;
        RECT -42.690 -119.625 -42.520 -116.685 ;
        RECT -42.220 -116.725 -42.010 -116.515 ;
        RECT -42.710 -119.895 -42.500 -119.625 ;
        RECT -42.200 -119.635 -42.030 -116.725 ;
        RECT -41.145 -119.605 -40.975 -116.685 ;
        RECT -10.275 -117.005 -8.785 -112.715 ;
        RECT -2.230 -117.005 -0.925 -112.715 ;
        RECT 1.955 -117.005 3.260 -112.715 ;
        RECT 7.155 -117.005 8.460 -112.715 ;
        RECT 14.445 -117.005 15.750 -112.715 ;
        RECT 20.515 -117.005 21.820 -112.715 ;
        RECT 30.245 -117.005 31.550 -112.715 ;
        RECT 37.715 -117.005 39.020 -112.715 ;
        RECT 88.885 -112.710 89.150 -112.500 ;
        RECT 89.425 -112.530 89.595 -109.545 ;
        RECT 89.990 -112.500 90.160 -109.490 ;
        RECT 90.460 -109.580 90.670 -109.300 ;
        RECT 89.930 -112.710 90.210 -112.500 ;
        RECT 90.480 -112.530 90.650 -109.580 ;
        RECT 90.970 -112.500 91.140 -109.490 ;
        RECT 90.920 -112.710 91.200 -112.500 ;
        RECT 88.885 -112.880 91.200 -112.710 ;
        RECT -28.600 -117.840 -25.460 -117.670 ;
        RECT -35.835 -117.955 -35.665 -117.935 ;
        RECT -35.865 -119.220 -35.635 -117.955 ;
        RECT -34.855 -118.895 -34.685 -117.935 ;
        RECT -33.875 -118.895 -33.705 -117.935 ;
        RECT -31.650 -117.955 -31.480 -117.935 ;
        RECT -32.755 -118.365 -32.470 -118.045 ;
        RECT -33.470 -118.610 -32.470 -118.365 ;
        RECT -34.885 -119.220 -34.655 -118.895 ;
        RECT -33.905 -119.220 -33.675 -118.895 ;
        RECT -35.865 -119.260 -33.675 -119.220 ;
        RECT -33.470 -119.260 -33.240 -118.610 ;
        RECT -32.755 -118.865 -32.470 -118.610 ;
        RECT -36.885 -119.445 -36.045 -119.295 ;
        RECT -43.205 -120.090 -42.500 -119.895 ;
        RECT -42.225 -119.900 -42.015 -119.635 ;
        RECT -41.165 -119.900 -40.955 -119.605 ;
        RECT -42.225 -120.080 -40.955 -119.900 ;
        RECT -36.920 -119.665 -36.045 -119.445 ;
        RECT -35.865 -119.450 -33.240 -119.260 ;
        RECT -31.680 -119.220 -31.450 -117.955 ;
        RECT -30.670 -118.895 -30.500 -117.935 ;
        RECT -29.690 -118.895 -29.520 -117.935 ;
        RECT -28.600 -118.065 -28.420 -117.840 ;
        RECT -30.700 -119.220 -30.470 -118.895 ;
        RECT -29.720 -119.220 -29.490 -118.895 ;
        RECT -31.680 -119.260 -29.490 -119.220 ;
        RECT -29.215 -119.140 -28.845 -118.300 ;
        RECT -28.595 -118.435 -28.425 -118.065 ;
        RECT -29.215 -119.260 -28.850 -119.140 ;
        RECT -32.700 -119.350 -31.860 -119.295 ;
        RECT -32.875 -119.355 -31.860 -119.350 ;
        RECT -43.205 -120.150 -42.990 -120.090 ;
        RECT -43.895 -120.425 -42.990 -120.150 ;
        RECT -43.205 -120.775 -42.990 -120.425 ;
        RECT -42.555 -120.310 -41.780 -120.260 ;
        RECT -39.990 -120.310 -39.330 -120.050 ;
        RECT -42.555 -120.490 -39.330 -120.310 ;
        RECT -42.555 -120.535 -41.780 -120.490 ;
        RECT -46.185 -121.075 -43.395 -120.875 ;
        RECT -43.205 -120.975 -41.435 -120.775 ;
        RECT -46.185 -121.090 -43.635 -121.075 ;
        RECT -75.700 -121.535 -73.030 -121.195 ;
        RECT -71.045 -121.310 -67.880 -121.140 ;
        RECT -75.695 -122.250 -75.525 -121.790 ;
        RECT -75.725 -122.555 -75.495 -122.250 ;
        RECT -75.205 -122.330 -75.035 -121.535 ;
        RECT -74.715 -122.250 -74.545 -121.790 ;
        RECT -75.875 -122.665 -75.495 -122.555 ;
        RECT -76.290 -122.715 -75.495 -122.665 ;
        RECT -74.745 -122.715 -74.515 -122.250 ;
        RECT -74.225 -122.330 -74.055 -121.535 ;
        RECT -73.735 -122.250 -73.565 -121.790 ;
        RECT -73.765 -122.715 -73.535 -122.250 ;
        RECT -73.245 -122.330 -73.075 -121.535 ;
        RECT -71.505 -122.010 -71.335 -121.540 ;
        RECT -71.045 -121.600 -70.825 -121.310 ;
        RECT -71.525 -122.225 -71.320 -122.010 ;
        RECT -71.015 -122.080 -70.845 -121.600 ;
        RECT -70.525 -122.015 -70.355 -121.540 ;
        RECT -70.060 -121.655 -69.840 -121.310 ;
        RECT -71.530 -122.260 -71.320 -122.225 ;
        RECT -70.540 -122.260 -70.335 -122.015 ;
        RECT -70.035 -122.080 -69.865 -121.655 ;
        RECT -69.545 -122.015 -69.375 -121.540 ;
        RECT -69.080 -121.655 -68.860 -121.310 ;
        RECT -69.570 -122.260 -69.365 -122.015 ;
        RECT -69.055 -122.080 -68.885 -121.655 ;
        RECT -68.565 -122.055 -68.395 -121.540 ;
        RECT -68.100 -121.600 -67.880 -121.310 ;
        RECT -66.985 -121.535 -59.530 -121.195 ;
        RECT -57.545 -121.310 -54.380 -121.140 ;
        RECT -68.075 -121.950 -67.905 -121.600 ;
        RECT -68.580 -122.260 -68.375 -122.055 ;
        RECT -71.530 -122.430 -68.375 -122.260 ;
        RECT -76.290 -122.850 -73.535 -122.715 ;
        RECT -76.285 -122.860 -73.535 -122.850 ;
        RECT -75.875 -122.905 -73.535 -122.860 ;
        RECT -73.355 -122.575 -72.515 -122.500 ;
        RECT -71.530 -122.575 -70.655 -122.430 ;
        RECT -73.355 -122.840 -70.655 -122.575 ;
        RECT -68.110 -122.625 -67.875 -121.950 ;
        RECT -66.980 -122.250 -66.810 -121.790 ;
        RECT -67.010 -122.555 -66.780 -122.250 ;
        RECT -66.490 -122.330 -66.320 -121.535 ;
        RECT -66.000 -122.250 -65.830 -121.790 ;
        RECT -73.355 -122.870 -72.515 -122.840 ;
        RECT -75.725 -122.945 -73.535 -122.905 ;
        RECT -75.725 -123.270 -75.495 -122.945 ;
        RECT -74.745 -123.270 -74.515 -122.945 ;
        RECT -85.130 -123.900 -84.910 -123.700 ;
        RECT -80.670 -123.900 -79.985 -123.550 ;
        RECT -85.130 -123.915 -79.985 -123.900 ;
        RECT -87.330 -124.215 -85.560 -124.015 ;
        RECT -85.370 -124.115 -79.985 -123.915 ;
        RECT -89.010 -124.500 -88.660 -124.490 ;
        RECT -86.985 -124.500 -86.210 -124.455 ;
        RECT -89.010 -124.680 -86.210 -124.500 ;
        RECT -96.805 -125.595 -95.670 -125.585 ;
        RECT -93.615 -125.715 -93.245 -125.585 ;
        RECT -98.535 -125.885 -97.950 -125.810 ;
        RECT -95.940 -125.875 -95.265 -125.835 ;
        RECT -96.040 -125.885 -95.265 -125.875 ;
        RECT -98.535 -126.065 -95.265 -125.885 ;
        RECT -92.680 -125.930 -89.605 -125.500 ;
        RECT -98.535 -126.425 -97.950 -126.065 ;
        RECT -96.040 -126.075 -95.265 -126.065 ;
        RECT -95.940 -126.105 -95.265 -126.075 ;
        RECT -95.025 -125.990 -92.930 -125.950 ;
        RECT -95.025 -126.140 -92.875 -125.990 ;
        RECT -102.700 -126.860 -99.715 -126.690 ;
        RECT -111.645 -128.345 -111.405 -127.685 ;
        RECT -111.120 -127.885 -110.950 -126.930 ;
        RECT -110.000 -127.135 -99.715 -126.860 ;
        RECT -110.000 -127.440 -100.795 -127.135 ;
        RECT -110.000 -128.345 -109.420 -127.440 ;
        RECT -95.025 -127.860 -94.855 -126.140 ;
        RECT -94.045 -127.860 -93.875 -126.140 ;
        RECT -93.180 -126.885 -92.875 -126.140 ;
        RECT -91.980 -126.710 -91.810 -125.930 ;
        RECT -91.490 -126.710 -91.320 -126.170 ;
        RECT -91.000 -126.710 -90.830 -125.930 ;
        RECT -90.510 -126.710 -90.340 -126.170 ;
        RECT -89.010 -126.655 -88.660 -124.680 ;
        RECT -86.985 -124.730 -86.210 -124.680 ;
        RECT -85.775 -124.565 -85.560 -124.215 ;
        RECT -85.775 -124.840 -84.870 -124.565 ;
        RECT -85.775 -124.900 -85.560 -124.840 ;
        RECT -87.810 -125.090 -86.540 -124.910 ;
        RECT -87.810 -125.385 -87.600 -125.090 ;
        RECT -86.750 -125.355 -86.540 -125.090 ;
        RECT -86.265 -125.095 -85.560 -124.900 ;
        RECT -92.570 -126.885 -92.205 -126.855 ;
        RECT -93.180 -126.950 -92.205 -126.885 ;
        RECT -93.070 -127.090 -92.205 -126.950 ;
        RECT -92.570 -127.155 -92.205 -127.090 ;
        RECT -90.020 -127.005 -88.630 -126.655 ;
        RECT -91.980 -127.865 -91.810 -127.325 ;
        RECT -91.000 -127.865 -90.830 -127.325 ;
        RECT -90.020 -127.865 -89.850 -127.005 ;
        RECT -87.790 -128.305 -87.620 -125.385 ;
        RECT -86.735 -128.265 -86.565 -125.355 ;
        RECT -86.265 -125.365 -86.055 -125.095 ;
        RECT -113.290 -128.430 -109.270 -128.345 ;
        RECT -113.290 -128.960 -108.850 -128.430 ;
        RECT -86.755 -128.475 -86.545 -128.265 ;
        RECT -86.245 -128.305 -86.075 -125.365 ;
        RECT -85.755 -128.255 -85.585 -125.265 ;
        RECT -84.700 -125.335 -84.485 -124.115 ;
        RECT -80.670 -124.380 -79.985 -124.115 ;
        RECT -75.695 -124.230 -75.525 -123.270 ;
        RECT -74.715 -124.230 -74.545 -123.270 ;
        RECT -73.765 -124.210 -73.535 -122.945 ;
        RECT -71.530 -123.265 -70.655 -122.840 ;
        RECT -68.735 -122.995 -67.875 -122.625 ;
        RECT -71.530 -123.435 -68.390 -123.265 ;
        RECT -71.530 -123.655 -71.320 -123.435 ;
        RECT -71.505 -124.155 -71.335 -123.655 ;
        RECT -71.015 -124.070 -70.845 -123.615 ;
        RECT -70.530 -123.705 -70.350 -123.435 ;
        RECT -69.560 -123.615 -69.380 -123.435 ;
        RECT -73.735 -124.230 -73.565 -124.210 ;
        RECT -71.040 -124.325 -70.830 -124.070 ;
        RECT -70.525 -124.155 -70.355 -123.705 ;
        RECT -70.035 -124.045 -69.865 -123.615 ;
        RECT -69.560 -123.705 -69.375 -123.615 ;
        RECT -70.060 -124.325 -69.850 -124.045 ;
        RECT -69.545 -124.155 -69.375 -123.705 ;
        RECT -69.055 -124.050 -68.885 -123.615 ;
        RECT -68.570 -123.695 -68.390 -123.435 ;
        RECT -69.090 -124.325 -68.880 -124.050 ;
        RECT -68.565 -124.155 -68.395 -123.695 ;
        RECT -68.110 -123.730 -67.875 -122.995 ;
        RECT -67.650 -122.715 -66.780 -122.555 ;
        RECT -66.030 -122.715 -65.800 -122.250 ;
        RECT -65.510 -122.330 -65.340 -121.535 ;
        RECT -65.020 -122.250 -64.850 -121.790 ;
        RECT -65.050 -122.715 -64.820 -122.250 ;
        RECT -64.530 -122.330 -64.360 -121.535 ;
        RECT -67.650 -122.905 -64.820 -122.715 ;
        RECT -64.640 -122.525 -63.800 -122.500 ;
        RECT -63.500 -122.525 -63.200 -122.160 ;
        RECT -64.640 -122.815 -63.200 -122.525 ;
        RECT -62.925 -122.610 -62.625 -122.035 ;
        RECT -62.195 -122.250 -62.025 -121.790 ;
        RECT -62.225 -122.555 -61.995 -122.250 ;
        RECT -61.705 -122.330 -61.535 -121.535 ;
        RECT -61.215 -122.250 -61.045 -121.790 ;
        RECT -62.375 -122.610 -61.995 -122.555 ;
        RECT -64.640 -122.870 -63.800 -122.815 ;
        RECT -63.500 -122.820 -63.200 -122.815 ;
        RECT -62.950 -122.715 -61.995 -122.610 ;
        RECT -61.245 -122.715 -61.015 -122.250 ;
        RECT -60.725 -122.330 -60.555 -121.535 ;
        RECT -60.235 -122.250 -60.065 -121.790 ;
        RECT -60.265 -122.715 -60.035 -122.250 ;
        RECT -59.745 -122.330 -59.575 -121.535 ;
        RECT -58.020 -122.010 -57.790 -121.400 ;
        RECT -57.545 -121.600 -57.325 -121.310 ;
        RECT -58.025 -122.060 -57.790 -122.010 ;
        RECT -58.025 -122.225 -57.820 -122.060 ;
        RECT -57.515 -122.080 -57.345 -121.600 ;
        RECT -57.025 -122.015 -56.855 -121.540 ;
        RECT -56.560 -121.655 -56.340 -121.310 ;
        RECT -58.030 -122.260 -57.820 -122.225 ;
        RECT -57.040 -122.260 -56.835 -122.015 ;
        RECT -56.535 -122.080 -56.365 -121.655 ;
        RECT -56.045 -122.015 -55.875 -121.540 ;
        RECT -55.580 -121.655 -55.360 -121.310 ;
        RECT -56.070 -122.260 -55.865 -122.015 ;
        RECT -55.555 -122.080 -55.385 -121.655 ;
        RECT -55.065 -122.055 -54.895 -121.540 ;
        RECT -54.600 -121.600 -54.380 -121.310 ;
        RECT -53.485 -121.535 -46.405 -121.195 ;
        RECT -54.575 -121.950 -54.405 -121.600 ;
        RECT -55.080 -122.260 -54.875 -122.055 ;
        RECT -58.030 -122.430 -54.875 -122.260 ;
        RECT -62.950 -122.835 -60.035 -122.715 ;
        RECT -67.650 -123.025 -67.285 -122.905 ;
        RECT -68.075 -124.100 -67.905 -123.730 ;
        RECT -67.655 -123.865 -67.285 -123.025 ;
        RECT -67.010 -122.945 -64.820 -122.905 ;
        RECT -67.010 -123.270 -66.780 -122.945 ;
        RECT -66.030 -123.270 -65.800 -122.945 ;
        RECT -68.080 -124.325 -67.900 -124.100 ;
        RECT -66.980 -124.230 -66.810 -123.270 ;
        RECT -66.000 -124.230 -65.830 -123.270 ;
        RECT -65.050 -124.210 -64.820 -122.945 ;
        RECT -64.030 -123.505 -63.745 -123.300 ;
        RECT -62.950 -123.505 -62.725 -122.835 ;
        RECT -62.375 -122.905 -60.035 -122.835 ;
        RECT -59.855 -122.540 -59.015 -122.500 ;
        RECT -58.030 -122.540 -57.155 -122.430 ;
        RECT -59.855 -122.825 -57.155 -122.540 ;
        RECT -54.610 -122.625 -54.375 -121.950 ;
        RECT -53.480 -122.250 -53.310 -121.790 ;
        RECT -53.510 -122.555 -53.280 -122.250 ;
        RECT -52.990 -122.330 -52.820 -121.535 ;
        RECT -52.500 -122.250 -52.330 -121.790 ;
        RECT -59.855 -122.870 -59.015 -122.825 ;
        RECT -62.225 -122.945 -60.035 -122.905 ;
        RECT -62.225 -123.270 -61.995 -122.945 ;
        RECT -61.245 -123.270 -61.015 -122.945 ;
        RECT -64.030 -123.730 -62.725 -123.505 ;
        RECT -64.030 -124.120 -63.745 -123.730 ;
        RECT -65.020 -124.230 -64.850 -124.210 ;
        RECT -62.195 -124.230 -62.025 -123.270 ;
        RECT -61.215 -124.230 -61.045 -123.270 ;
        RECT -60.265 -124.210 -60.035 -122.945 ;
        RECT -58.030 -123.265 -57.155 -122.825 ;
        RECT -55.235 -122.995 -54.375 -122.625 ;
        RECT -58.030 -123.435 -54.890 -123.265 ;
        RECT -58.030 -123.655 -57.820 -123.435 ;
        RECT -58.005 -124.155 -57.835 -123.655 ;
        RECT -57.515 -124.070 -57.345 -123.615 ;
        RECT -57.030 -123.705 -56.850 -123.435 ;
        RECT -56.060 -123.615 -55.880 -123.435 ;
        RECT -60.235 -124.230 -60.065 -124.210 ;
        RECT -71.040 -124.495 -67.900 -124.325 ;
        RECT -57.540 -124.325 -57.330 -124.070 ;
        RECT -57.025 -124.155 -56.855 -123.705 ;
        RECT -56.535 -124.045 -56.365 -123.615 ;
        RECT -56.060 -123.705 -55.875 -123.615 ;
        RECT -56.560 -124.325 -56.350 -124.045 ;
        RECT -56.045 -124.155 -55.875 -123.705 ;
        RECT -55.555 -124.050 -55.385 -123.615 ;
        RECT -55.070 -123.695 -54.890 -123.435 ;
        RECT -55.590 -124.325 -55.380 -124.050 ;
        RECT -55.065 -124.155 -54.895 -123.695 ;
        RECT -54.610 -123.730 -54.375 -122.995 ;
        RECT -54.150 -122.715 -53.280 -122.555 ;
        RECT -52.530 -122.715 -52.300 -122.250 ;
        RECT -52.010 -122.330 -51.840 -121.535 ;
        RECT -51.520 -122.250 -51.350 -121.790 ;
        RECT -51.550 -122.715 -51.320 -122.250 ;
        RECT -51.030 -122.330 -50.860 -121.535 ;
        RECT -54.150 -122.905 -51.320 -122.715 ;
        RECT -51.140 -122.525 -50.300 -122.500 ;
        RECT -51.140 -122.585 -50.125 -122.525 ;
        RECT -49.840 -122.585 -49.540 -122.155 ;
        RECT -49.070 -122.250 -48.900 -121.790 ;
        RECT -49.100 -122.555 -48.870 -122.250 ;
        RECT -48.580 -122.330 -48.410 -121.535 ;
        RECT -48.090 -122.250 -47.920 -121.790 ;
        RECT -49.250 -122.585 -48.870 -122.555 ;
        RECT -51.140 -122.715 -48.870 -122.585 ;
        RECT -48.120 -122.715 -47.890 -122.250 ;
        RECT -47.600 -122.330 -47.430 -121.535 ;
        RECT -47.110 -122.250 -46.940 -121.790 ;
        RECT -47.140 -122.715 -46.910 -122.250 ;
        RECT -46.620 -122.330 -46.450 -121.535 ;
        RECT -46.185 -122.500 -45.990 -121.090 ;
        RECT -43.855 -121.290 -43.635 -121.090 ;
        RECT -51.140 -122.795 -46.910 -122.715 ;
        RECT -51.140 -122.815 -50.125 -122.795 ;
        RECT -49.840 -122.815 -49.540 -122.795 ;
        RECT -51.140 -122.870 -50.300 -122.815 ;
        RECT -49.250 -122.905 -46.910 -122.795 ;
        RECT -46.730 -122.870 -45.890 -122.500 ;
        RECT -43.825 -122.785 -43.655 -121.290 ;
        RECT -43.335 -122.660 -43.165 -121.245 ;
        RECT -54.150 -123.025 -53.785 -122.905 ;
        RECT -54.575 -124.100 -54.405 -123.730 ;
        RECT -54.155 -123.865 -53.785 -123.025 ;
        RECT -53.510 -122.945 -51.320 -122.905 ;
        RECT -53.510 -123.270 -53.280 -122.945 ;
        RECT -52.530 -123.270 -52.300 -122.945 ;
        RECT -54.580 -124.325 -54.400 -124.100 ;
        RECT -53.480 -124.230 -53.310 -123.270 ;
        RECT -52.500 -124.230 -52.330 -123.270 ;
        RECT -51.550 -124.210 -51.320 -122.945 ;
        RECT -49.100 -122.945 -46.910 -122.905 ;
        RECT -49.100 -123.270 -48.870 -122.945 ;
        RECT -48.120 -123.270 -47.890 -122.945 ;
        RECT -50.530 -124.120 -50.245 -123.300 ;
        RECT -51.520 -124.230 -51.350 -124.210 ;
        RECT -49.070 -124.230 -48.900 -123.270 ;
        RECT -48.090 -124.230 -47.920 -123.270 ;
        RECT -47.140 -124.210 -46.910 -122.945 ;
        RECT -43.365 -123.310 -43.130 -122.660 ;
        RECT -42.125 -122.710 -41.955 -121.245 ;
        RECT -41.660 -121.325 -41.435 -120.975 ;
        RECT -41.205 -120.845 -40.430 -120.800 ;
        RECT -38.615 -120.845 -37.905 -120.760 ;
        RECT -41.205 -121.015 -37.905 -120.845 ;
        RECT -41.205 -121.075 -40.430 -121.015 ;
        RECT -38.615 -121.080 -37.905 -121.015 ;
        RECT -42.155 -123.310 -41.920 -122.710 ;
        RECT -41.635 -122.785 -41.465 -121.325 ;
        RECT -41.145 -122.715 -40.975 -121.245 ;
        RECT -36.920 -121.525 -36.680 -119.665 ;
        RECT -36.325 -120.630 -36.155 -119.835 ;
        RECT -35.865 -119.915 -35.635 -119.450 ;
        RECT -35.835 -120.375 -35.665 -119.915 ;
        RECT -35.345 -120.630 -35.175 -119.835 ;
        RECT -34.885 -119.915 -34.655 -119.450 ;
        RECT -33.905 -119.610 -33.240 -119.450 ;
        RECT -34.855 -120.375 -34.685 -119.915 ;
        RECT -34.365 -120.630 -34.195 -119.835 ;
        RECT -33.905 -119.915 -33.675 -119.610 ;
        RECT -33.060 -119.665 -31.860 -119.355 ;
        RECT -31.680 -119.450 -28.850 -119.260 ;
        RECT -33.875 -120.375 -33.705 -119.915 ;
        RECT -33.060 -120.385 -32.760 -119.665 ;
        RECT -32.140 -120.630 -31.970 -119.835 ;
        RECT -31.680 -119.915 -31.450 -119.450 ;
        RECT -31.650 -120.375 -31.480 -119.915 ;
        RECT -31.160 -120.630 -30.990 -119.835 ;
        RECT -30.700 -119.915 -30.470 -119.450 ;
        RECT -29.720 -119.610 -28.850 -119.450 ;
        RECT -28.625 -119.170 -28.390 -118.435 ;
        RECT -28.105 -118.470 -27.935 -118.010 ;
        RECT -27.620 -118.115 -27.410 -117.840 ;
        RECT -28.110 -118.730 -27.930 -118.470 ;
        RECT -27.615 -118.550 -27.445 -118.115 ;
        RECT -27.125 -118.460 -26.955 -118.010 ;
        RECT -26.650 -118.120 -26.440 -117.840 ;
        RECT -27.125 -118.550 -26.940 -118.460 ;
        RECT -26.635 -118.550 -26.465 -118.120 ;
        RECT -26.145 -118.460 -25.975 -118.010 ;
        RECT -25.670 -118.095 -25.460 -117.840 ;
        RECT -15.100 -117.840 -11.960 -117.670 ;
        RECT -22.335 -117.955 -22.165 -117.935 ;
        RECT -27.120 -118.730 -26.940 -118.550 ;
        RECT -26.150 -118.730 -25.970 -118.460 ;
        RECT -25.655 -118.550 -25.485 -118.095 ;
        RECT -25.165 -118.510 -24.995 -118.010 ;
        RECT -25.180 -118.730 -24.970 -118.510 ;
        RECT -28.110 -118.900 -24.970 -118.730 ;
        RECT -28.625 -119.540 -27.765 -119.170 ;
        RECT -25.845 -119.435 -24.970 -118.900 ;
        RECT -22.365 -119.220 -22.135 -117.955 ;
        RECT -21.355 -118.895 -21.185 -117.935 ;
        RECT -20.375 -118.895 -20.205 -117.935 ;
        RECT -18.150 -117.955 -17.980 -117.935 ;
        RECT -19.255 -118.305 -18.970 -118.045 ;
        RECT -19.995 -118.615 -18.970 -118.305 ;
        RECT -21.385 -119.220 -21.155 -118.895 ;
        RECT -20.405 -119.220 -20.175 -118.895 ;
        RECT -22.365 -119.260 -20.175 -119.220 ;
        RECT -19.995 -119.260 -19.685 -118.615 ;
        RECT -19.255 -118.865 -18.970 -118.615 ;
        RECT -23.385 -119.330 -22.545 -119.295 ;
        RECT -30.670 -120.375 -30.500 -119.915 ;
        RECT -30.180 -120.630 -30.010 -119.835 ;
        RECT -29.720 -119.915 -29.490 -119.610 ;
        RECT -29.690 -120.375 -29.520 -119.915 ;
        RECT -28.625 -120.215 -28.390 -119.540 ;
        RECT -25.845 -119.735 -24.515 -119.435 ;
        RECT -23.495 -119.630 -22.545 -119.330 ;
        RECT -23.385 -119.665 -22.545 -119.630 ;
        RECT -22.365 -119.450 -19.685 -119.260 ;
        RECT -18.180 -119.220 -17.950 -117.955 ;
        RECT -17.170 -118.895 -17.000 -117.935 ;
        RECT -16.190 -118.895 -16.020 -117.935 ;
        RECT -15.100 -118.065 -14.920 -117.840 ;
        RECT -17.200 -119.220 -16.970 -118.895 ;
        RECT -16.220 -119.220 -15.990 -118.895 ;
        RECT -18.180 -119.260 -15.990 -119.220 ;
        RECT -15.715 -119.140 -15.345 -118.300 ;
        RECT -15.095 -118.435 -14.925 -118.065 ;
        RECT -15.715 -119.260 -15.350 -119.140 ;
        RECT -19.200 -119.350 -18.360 -119.295 ;
        RECT -28.125 -119.905 -24.970 -119.735 ;
        RECT -28.125 -120.110 -27.920 -119.905 ;
        RECT -28.595 -120.565 -28.425 -120.215 ;
        RECT -36.370 -120.970 -29.515 -120.630 ;
        RECT -28.620 -120.855 -28.400 -120.565 ;
        RECT -28.105 -120.625 -27.935 -120.110 ;
        RECT -27.615 -120.510 -27.445 -120.085 ;
        RECT -27.135 -120.150 -26.930 -119.905 ;
        RECT -27.640 -120.855 -27.420 -120.510 ;
        RECT -27.125 -120.625 -26.955 -120.150 ;
        RECT -26.635 -120.510 -26.465 -120.085 ;
        RECT -26.165 -120.150 -25.960 -119.905 ;
        RECT -25.180 -119.940 -24.970 -119.905 ;
        RECT -26.660 -120.855 -26.440 -120.510 ;
        RECT -26.145 -120.625 -25.975 -120.150 ;
        RECT -25.655 -120.565 -25.485 -120.085 ;
        RECT -25.180 -120.155 -24.975 -119.940 ;
        RECT -25.675 -120.855 -25.455 -120.565 ;
        RECT -25.165 -120.625 -24.995 -120.155 ;
        RECT -22.825 -120.630 -22.655 -119.835 ;
        RECT -22.365 -119.915 -22.135 -119.450 ;
        RECT -22.335 -120.375 -22.165 -119.915 ;
        RECT -21.845 -120.630 -21.675 -119.835 ;
        RECT -21.385 -119.915 -21.155 -119.450 ;
        RECT -20.405 -119.610 -19.685 -119.450 ;
        RECT -21.355 -120.375 -21.185 -119.915 ;
        RECT -20.865 -120.630 -20.695 -119.835 ;
        RECT -20.405 -119.915 -20.175 -119.610 ;
        RECT -19.500 -119.665 -18.360 -119.350 ;
        RECT -18.180 -119.450 -15.350 -119.260 ;
        RECT -20.375 -120.375 -20.205 -119.915 ;
        RECT -19.500 -120.460 -19.200 -119.665 ;
        RECT -18.640 -120.630 -18.470 -119.835 ;
        RECT -18.180 -119.915 -17.950 -119.450 ;
        RECT -18.150 -120.375 -17.980 -119.915 ;
        RECT -17.660 -120.630 -17.490 -119.835 ;
        RECT -17.200 -119.915 -16.970 -119.450 ;
        RECT -16.220 -119.610 -15.350 -119.450 ;
        RECT -15.125 -119.170 -14.890 -118.435 ;
        RECT -14.605 -118.470 -14.435 -118.010 ;
        RECT -14.120 -118.115 -13.910 -117.840 ;
        RECT -14.610 -118.730 -14.430 -118.470 ;
        RECT -14.115 -118.550 -13.945 -118.115 ;
        RECT -13.625 -118.460 -13.455 -118.010 ;
        RECT -13.150 -118.120 -12.940 -117.840 ;
        RECT -13.625 -118.550 -13.440 -118.460 ;
        RECT -13.135 -118.550 -12.965 -118.120 ;
        RECT -12.645 -118.460 -12.475 -118.010 ;
        RECT -12.170 -118.095 -11.960 -117.840 ;
        RECT -13.620 -118.730 -13.440 -118.550 ;
        RECT -12.650 -118.730 -12.470 -118.460 ;
        RECT -12.155 -118.550 -11.985 -118.095 ;
        RECT -11.665 -118.510 -11.495 -118.010 ;
        RECT -10.275 -118.310 39.020 -117.005 ;
        RECT 67.750 -116.370 70.320 -115.555 ;
        RECT 76.550 -116.370 77.655 -116.230 ;
        RECT 67.750 -117.020 77.655 -116.370 ;
        RECT 67.750 -117.680 70.320 -117.020 ;
        RECT -11.680 -118.730 -11.470 -118.510 ;
        RECT -14.610 -118.900 -11.470 -118.730 ;
        RECT -15.125 -119.540 -14.265 -119.170 ;
        RECT -12.345 -119.445 -11.470 -118.900 ;
        RECT -17.170 -120.375 -17.000 -119.915 ;
        RECT -16.680 -120.630 -16.510 -119.835 ;
        RECT -16.220 -119.915 -15.990 -119.610 ;
        RECT -16.190 -120.375 -16.020 -119.915 ;
        RECT -15.125 -120.215 -14.890 -119.540 ;
        RECT -12.345 -119.735 -11.095 -119.445 ;
        RECT -14.625 -119.745 -11.095 -119.735 ;
        RECT -14.625 -119.905 -11.470 -119.745 ;
        RECT -14.625 -120.110 -14.420 -119.905 ;
        RECT -15.095 -120.565 -14.925 -120.215 ;
        RECT -35.130 -121.170 -34.575 -120.970 ;
        RECT -35.185 -121.210 -34.500 -121.170 ;
        RECT -31.075 -121.210 -30.520 -120.970 ;
        RECT -28.620 -121.025 -25.455 -120.855 ;
        RECT -22.870 -120.640 -20.200 -120.630 ;
        RECT -18.685 -120.640 -16.015 -120.630 ;
        RECT -22.870 -120.970 -16.015 -120.640 ;
        RECT -15.120 -120.855 -14.900 -120.565 ;
        RECT -14.605 -120.625 -14.435 -120.110 ;
        RECT -14.115 -120.510 -13.945 -120.085 ;
        RECT -13.635 -120.150 -13.430 -119.905 ;
        RECT -14.140 -120.855 -13.920 -120.510 ;
        RECT -13.625 -120.625 -13.455 -120.150 ;
        RECT -13.135 -120.510 -12.965 -120.085 ;
        RECT -12.665 -120.150 -12.460 -119.905 ;
        RECT -11.680 -119.940 -11.470 -119.905 ;
        RECT -13.160 -120.855 -12.940 -120.510 ;
        RECT -12.645 -120.625 -12.475 -120.150 ;
        RECT -12.155 -120.565 -11.985 -120.085 ;
        RECT -11.680 -120.155 -11.475 -119.940 ;
        RECT -12.175 -120.855 -11.955 -120.565 ;
        RECT -11.665 -120.625 -11.495 -120.155 ;
        RECT -22.085 -121.200 -21.530 -120.970 ;
        RECT -21.170 -120.980 -18.570 -120.970 ;
        RECT -22.200 -121.210 -21.515 -121.200 ;
        RECT -17.695 -121.210 -17.140 -120.970 ;
        RECT -15.120 -121.025 -11.955 -120.855 ;
        RECT -10.275 -121.200 -8.785 -118.310 ;
        RECT -5.045 -119.635 -4.395 -118.310 ;
        RECT -3.515 -119.635 -2.865 -118.310 ;
        RECT -1.930 -119.635 -1.280 -118.310 ;
        RECT 0.300 -119.635 0.950 -118.310 ;
        RECT -5.110 -119.960 1.260 -119.635 ;
        RECT -10.275 -121.210 -8.350 -121.200 ;
        RECT -35.270 -121.405 -8.345 -121.210 ;
        RECT -35.185 -121.470 -34.500 -121.405 ;
        RECT -22.200 -121.500 -21.515 -121.405 ;
        RECT -9.010 -121.500 -8.350 -121.405 ;
        RECT -36.925 -122.210 -36.625 -121.525 ;
        RECT -24.375 -121.670 -23.690 -121.615 ;
        RECT -19.645 -121.670 -18.985 -121.620 ;
        RECT -35.270 -121.865 -6.620 -121.670 ;
        RECT -24.375 -121.915 -23.690 -121.865 ;
        RECT -19.645 -121.920 -18.985 -121.865 ;
        RECT -33.240 -122.100 -32.580 -122.060 ;
        RECT -10.625 -122.100 -9.965 -122.050 ;
        RECT -41.175 -123.310 -40.940 -122.715 ;
        RECT -38.620 -123.310 -38.095 -123.280 ;
        RECT -44.265 -123.720 -38.095 -123.310 ;
        RECT -38.620 -123.755 -38.095 -123.720 ;
        RECT -36.920 -124.000 -36.680 -122.210 ;
        RECT -35.270 -122.295 -9.965 -122.100 ;
        RECT -33.240 -122.360 -32.580 -122.295 ;
        RECT -10.625 -122.350 -9.965 -122.295 ;
        RECT -36.330 -122.870 -33.660 -122.530 ;
        RECT -31.675 -122.645 -28.510 -122.475 ;
        RECT -36.325 -123.585 -36.155 -123.125 ;
        RECT -36.355 -123.890 -36.125 -123.585 ;
        RECT -35.835 -123.665 -35.665 -122.870 ;
        RECT -35.345 -123.585 -35.175 -123.125 ;
        RECT -36.505 -124.000 -36.125 -123.890 ;
        RECT -36.920 -124.050 -36.125 -124.000 ;
        RECT -35.375 -124.050 -35.145 -123.585 ;
        RECT -34.855 -123.665 -34.685 -122.870 ;
        RECT -34.365 -123.585 -34.195 -123.125 ;
        RECT -34.395 -124.050 -34.165 -123.585 ;
        RECT -33.875 -123.665 -33.705 -122.870 ;
        RECT -32.135 -123.345 -31.965 -122.875 ;
        RECT -31.675 -122.935 -31.455 -122.645 ;
        RECT -32.155 -123.560 -31.950 -123.345 ;
        RECT -31.645 -123.415 -31.475 -122.935 ;
        RECT -31.155 -123.350 -30.985 -122.875 ;
        RECT -30.690 -122.990 -30.470 -122.645 ;
        RECT -32.160 -123.595 -31.950 -123.560 ;
        RECT -31.170 -123.595 -30.965 -123.350 ;
        RECT -30.665 -123.415 -30.495 -122.990 ;
        RECT -30.175 -123.350 -30.005 -122.875 ;
        RECT -29.710 -122.990 -29.490 -122.645 ;
        RECT -30.200 -123.595 -29.995 -123.350 ;
        RECT -29.685 -123.415 -29.515 -122.990 ;
        RECT -29.195 -123.390 -29.025 -122.875 ;
        RECT -28.730 -122.935 -28.510 -122.645 ;
        RECT -27.615 -122.870 -20.160 -122.530 ;
        RECT -18.175 -122.645 -15.010 -122.475 ;
        RECT -28.705 -123.285 -28.535 -122.935 ;
        RECT -29.210 -123.595 -29.005 -123.390 ;
        RECT -32.160 -123.765 -29.005 -123.595 ;
        RECT -36.920 -124.185 -34.165 -124.050 ;
        RECT -36.915 -124.195 -34.165 -124.185 ;
        RECT -47.110 -124.230 -46.940 -124.210 ;
        RECT -36.505 -124.240 -34.165 -124.195 ;
        RECT -33.985 -123.910 -33.145 -123.835 ;
        RECT -32.160 -123.910 -31.285 -123.765 ;
        RECT -33.985 -124.175 -31.285 -123.910 ;
        RECT -28.740 -123.960 -28.505 -123.285 ;
        RECT -27.610 -123.585 -27.440 -123.125 ;
        RECT -27.640 -123.890 -27.410 -123.585 ;
        RECT -27.120 -123.665 -26.950 -122.870 ;
        RECT -26.630 -123.585 -26.460 -123.125 ;
        RECT -33.985 -124.205 -33.145 -124.175 ;
        RECT -57.540 -124.495 -54.400 -124.325 ;
        RECT -36.355 -124.280 -34.165 -124.240 ;
        RECT -36.355 -124.605 -36.125 -124.280 ;
        RECT -35.375 -124.605 -35.145 -124.280 ;
        RECT -83.570 -124.990 -83.045 -124.630 ;
        RECT -85.765 -128.475 -85.555 -128.255 ;
        RECT -84.695 -128.305 -84.525 -125.335 ;
        RECT -86.755 -128.645 -85.555 -128.475 ;
        RECT -113.290 -129.095 -109.270 -128.960 ;
        RECT -114.355 -131.310 -109.440 -131.155 ;
        RECT -114.355 -131.635 -107.965 -131.310 ;
        RECT -114.355 -131.730 -109.440 -131.635 ;
        RECT -114.275 -137.155 -114.105 -132.575 ;
        RECT -113.785 -133.615 -113.615 -131.730 ;
        RECT -111.720 -132.085 -109.515 -131.915 ;
        RECT -112.210 -134.435 -112.040 -132.575 ;
        RECT -111.720 -134.115 -111.550 -132.085 ;
        RECT -110.670 -132.100 -109.515 -132.085 ;
        RECT -111.230 -134.435 -111.060 -132.575 ;
        RECT -110.670 -132.630 -110.495 -132.100 ;
        RECT -110.665 -134.115 -110.495 -132.630 ;
        RECT -110.175 -134.115 -110.005 -132.575 ;
        RECT -109.690 -132.620 -109.515 -132.100 ;
        RECT -109.685 -134.115 -109.515 -132.620 ;
        RECT -110.180 -134.430 -110.005 -134.115 ;
        RECT -109.115 -134.430 -108.945 -132.580 ;
        RECT -108.625 -134.120 -108.455 -131.635 ;
        RECT -94.895 -132.505 -94.725 -131.465 ;
        RECT -93.915 -132.505 -93.745 -131.465 ;
        RECT -92.935 -132.505 -92.765 -131.465 ;
        RECT -90.030 -132.540 -89.860 -130.820 ;
        RECT -89.050 -132.540 -88.880 -130.820 ;
        RECT -86.985 -131.355 -86.815 -130.815 ;
        RECT -86.005 -131.355 -85.835 -130.815 ;
        RECT -87.575 -131.590 -87.210 -131.525 ;
        RECT -88.075 -131.730 -87.210 -131.590 ;
        RECT -88.185 -131.795 -87.210 -131.730 ;
        RECT -88.185 -132.540 -87.880 -131.795 ;
        RECT -87.575 -131.825 -87.210 -131.795 ;
        RECT -85.025 -131.675 -84.855 -130.815 ;
        RECT -83.515 -131.675 -83.165 -124.990 ;
        RECT -36.325 -125.565 -36.155 -124.605 ;
        RECT -35.345 -125.565 -35.175 -124.605 ;
        RECT -34.395 -125.545 -34.165 -124.280 ;
        RECT -32.160 -124.600 -31.285 -124.175 ;
        RECT -29.365 -124.330 -28.505 -123.960 ;
        RECT -32.160 -124.770 -29.020 -124.600 ;
        RECT -32.160 -124.990 -31.950 -124.770 ;
        RECT -32.135 -125.490 -31.965 -124.990 ;
        RECT -31.645 -125.405 -31.475 -124.950 ;
        RECT -31.160 -125.040 -30.980 -124.770 ;
        RECT -30.190 -124.950 -30.010 -124.770 ;
        RECT -34.365 -125.565 -34.195 -125.545 ;
        RECT -31.670 -125.660 -31.460 -125.405 ;
        RECT -31.155 -125.490 -30.985 -125.040 ;
        RECT -30.665 -125.380 -30.495 -124.950 ;
        RECT -30.190 -125.040 -30.005 -124.950 ;
        RECT -30.690 -125.660 -30.480 -125.380 ;
        RECT -30.175 -125.490 -30.005 -125.040 ;
        RECT -29.685 -125.385 -29.515 -124.950 ;
        RECT -29.200 -125.030 -29.020 -124.770 ;
        RECT -29.720 -125.660 -29.510 -125.385 ;
        RECT -29.195 -125.490 -29.025 -125.030 ;
        RECT -28.740 -125.065 -28.505 -124.330 ;
        RECT -28.280 -124.050 -27.410 -123.890 ;
        RECT -26.660 -124.050 -26.430 -123.585 ;
        RECT -26.140 -123.665 -25.970 -122.870 ;
        RECT -25.650 -123.585 -25.480 -123.125 ;
        RECT -25.680 -124.050 -25.450 -123.585 ;
        RECT -25.160 -123.665 -24.990 -122.870 ;
        RECT -28.280 -124.240 -25.450 -124.050 ;
        RECT -25.270 -123.860 -24.430 -123.835 ;
        RECT -24.130 -123.860 -23.830 -123.495 ;
        RECT -25.270 -124.150 -23.830 -123.860 ;
        RECT -23.555 -123.945 -23.255 -123.370 ;
        RECT -22.825 -123.585 -22.655 -123.125 ;
        RECT -22.855 -123.890 -22.625 -123.585 ;
        RECT -22.335 -123.665 -22.165 -122.870 ;
        RECT -21.845 -123.585 -21.675 -123.125 ;
        RECT -23.005 -123.945 -22.625 -123.890 ;
        RECT -25.270 -124.205 -24.430 -124.150 ;
        RECT -24.130 -124.155 -23.830 -124.150 ;
        RECT -23.580 -124.050 -22.625 -123.945 ;
        RECT -21.875 -124.050 -21.645 -123.585 ;
        RECT -21.355 -123.665 -21.185 -122.870 ;
        RECT -20.865 -123.585 -20.695 -123.125 ;
        RECT -20.895 -124.050 -20.665 -123.585 ;
        RECT -20.375 -123.665 -20.205 -122.870 ;
        RECT -18.650 -123.345 -18.420 -122.735 ;
        RECT -18.175 -122.935 -17.955 -122.645 ;
        RECT -18.655 -123.395 -18.420 -123.345 ;
        RECT -18.655 -123.560 -18.450 -123.395 ;
        RECT -18.145 -123.415 -17.975 -122.935 ;
        RECT -17.655 -123.350 -17.485 -122.875 ;
        RECT -17.190 -122.990 -16.970 -122.645 ;
        RECT -18.660 -123.595 -18.450 -123.560 ;
        RECT -17.670 -123.595 -17.465 -123.350 ;
        RECT -17.165 -123.415 -16.995 -122.990 ;
        RECT -16.675 -123.350 -16.505 -122.875 ;
        RECT -16.210 -122.990 -15.990 -122.645 ;
        RECT -16.700 -123.595 -16.495 -123.350 ;
        RECT -16.185 -123.415 -16.015 -122.990 ;
        RECT -15.695 -123.390 -15.525 -122.875 ;
        RECT -15.230 -122.935 -15.010 -122.645 ;
        RECT -14.115 -122.870 -7.035 -122.530 ;
        RECT -15.205 -123.285 -15.035 -122.935 ;
        RECT -15.710 -123.595 -15.505 -123.390 ;
        RECT -18.660 -123.765 -15.505 -123.595 ;
        RECT -23.580 -124.170 -20.665 -124.050 ;
        RECT -28.280 -124.360 -27.915 -124.240 ;
        RECT -28.705 -125.435 -28.535 -125.065 ;
        RECT -28.285 -125.200 -27.915 -124.360 ;
        RECT -27.640 -124.280 -25.450 -124.240 ;
        RECT -27.640 -124.605 -27.410 -124.280 ;
        RECT -26.660 -124.605 -26.430 -124.280 ;
        RECT -28.710 -125.660 -28.530 -125.435 ;
        RECT -27.610 -125.565 -27.440 -124.605 ;
        RECT -26.630 -125.565 -26.460 -124.605 ;
        RECT -25.680 -125.545 -25.450 -124.280 ;
        RECT -24.660 -124.840 -24.375 -124.635 ;
        RECT -23.580 -124.840 -23.355 -124.170 ;
        RECT -23.005 -124.240 -20.665 -124.170 ;
        RECT -20.485 -123.875 -19.645 -123.835 ;
        RECT -18.660 -123.875 -17.785 -123.765 ;
        RECT -20.485 -124.160 -17.785 -123.875 ;
        RECT -15.240 -123.960 -15.005 -123.285 ;
        RECT -14.110 -123.585 -13.940 -123.125 ;
        RECT -14.140 -123.890 -13.910 -123.585 ;
        RECT -13.620 -123.665 -13.450 -122.870 ;
        RECT -13.130 -123.585 -12.960 -123.125 ;
        RECT -20.485 -124.205 -19.645 -124.160 ;
        RECT -22.855 -124.280 -20.665 -124.240 ;
        RECT -22.855 -124.605 -22.625 -124.280 ;
        RECT -21.875 -124.605 -21.645 -124.280 ;
        RECT -24.660 -125.065 -23.355 -124.840 ;
        RECT -24.660 -125.455 -24.375 -125.065 ;
        RECT -25.650 -125.565 -25.480 -125.545 ;
        RECT -22.825 -125.565 -22.655 -124.605 ;
        RECT -21.845 -125.565 -21.675 -124.605 ;
        RECT -20.895 -125.545 -20.665 -124.280 ;
        RECT -18.660 -124.600 -17.785 -124.160 ;
        RECT -15.865 -124.330 -15.005 -123.960 ;
        RECT -18.660 -124.770 -15.520 -124.600 ;
        RECT -18.660 -124.990 -18.450 -124.770 ;
        RECT -18.635 -125.490 -18.465 -124.990 ;
        RECT -18.145 -125.405 -17.975 -124.950 ;
        RECT -17.660 -125.040 -17.480 -124.770 ;
        RECT -16.690 -124.950 -16.510 -124.770 ;
        RECT -20.865 -125.565 -20.695 -125.545 ;
        RECT -31.670 -125.830 -28.530 -125.660 ;
        RECT -18.170 -125.660 -17.960 -125.405 ;
        RECT -17.655 -125.490 -17.485 -125.040 ;
        RECT -17.165 -125.380 -16.995 -124.950 ;
        RECT -16.690 -125.040 -16.505 -124.950 ;
        RECT -17.190 -125.660 -16.980 -125.380 ;
        RECT -16.675 -125.490 -16.505 -125.040 ;
        RECT -16.185 -125.385 -16.015 -124.950 ;
        RECT -15.700 -125.030 -15.520 -124.770 ;
        RECT -16.220 -125.660 -16.010 -125.385 ;
        RECT -15.695 -125.490 -15.525 -125.030 ;
        RECT -15.240 -125.065 -15.005 -124.330 ;
        RECT -14.780 -124.050 -13.910 -123.890 ;
        RECT -13.160 -124.050 -12.930 -123.585 ;
        RECT -12.640 -123.665 -12.470 -122.870 ;
        RECT -12.150 -123.585 -11.980 -123.125 ;
        RECT -12.180 -124.050 -11.950 -123.585 ;
        RECT -11.660 -123.665 -11.490 -122.870 ;
        RECT -14.780 -124.240 -11.950 -124.050 ;
        RECT -11.770 -123.860 -10.930 -123.835 ;
        RECT -11.770 -123.920 -10.755 -123.860 ;
        RECT -10.470 -123.920 -10.170 -123.490 ;
        RECT -9.700 -123.585 -9.530 -123.125 ;
        RECT -9.730 -123.890 -9.500 -123.585 ;
        RECT -9.210 -123.665 -9.040 -122.870 ;
        RECT -8.720 -123.585 -8.550 -123.125 ;
        RECT -9.880 -123.920 -9.500 -123.890 ;
        RECT -11.770 -124.050 -9.500 -123.920 ;
        RECT -8.750 -124.050 -8.520 -123.585 ;
        RECT -8.230 -123.665 -8.060 -122.870 ;
        RECT -7.740 -123.585 -7.570 -123.125 ;
        RECT -7.770 -124.050 -7.540 -123.585 ;
        RECT -7.250 -123.665 -7.080 -122.870 ;
        RECT -6.815 -123.835 -6.620 -121.865 ;
        RECT -5.050 -123.165 -4.880 -120.900 ;
        RECT -4.560 -121.940 -4.390 -119.960 ;
        RECT -2.495 -120.410 -0.290 -120.240 ;
        RECT -2.985 -122.760 -2.815 -120.900 ;
        RECT -2.495 -122.440 -2.325 -120.410 ;
        RECT -1.445 -120.425 -0.290 -120.410 ;
        RECT -2.005 -122.760 -1.835 -120.900 ;
        RECT -1.445 -120.955 -1.270 -120.425 ;
        RECT -1.440 -122.440 -1.270 -120.955 ;
        RECT -0.950 -122.440 -0.780 -120.900 ;
        RECT -0.465 -120.945 -0.290 -120.425 ;
        RECT -0.460 -122.440 -0.290 -120.945 ;
        RECT -0.955 -122.755 -0.780 -122.440 ;
        RECT 0.110 -122.755 0.280 -120.905 ;
        RECT 0.600 -122.445 0.770 -119.960 ;
        RECT 4.920 -120.710 5.675 -118.310 ;
        RECT 6.805 -120.620 7.425 -118.310 ;
        RECT 8.455 -120.620 9.075 -118.310 ;
        RECT 10.490 -120.520 11.170 -120.290 ;
        RECT 6.805 -120.710 9.380 -120.620 ;
        RECT -0.955 -122.760 0.280 -122.755 ;
        RECT 1.090 -122.760 1.260 -120.905 ;
        RECT -2.985 -122.930 -1.820 -122.760 ;
        RECT -0.955 -122.930 1.260 -122.760 ;
        RECT 4.920 -120.925 9.380 -120.710 ;
        RECT 4.920 -121.015 7.170 -120.925 ;
        RECT -5.805 -123.430 -4.880 -123.165 ;
        RECT -11.770 -124.130 -7.540 -124.050 ;
        RECT -11.770 -124.150 -10.755 -124.130 ;
        RECT -10.470 -124.150 -10.170 -124.130 ;
        RECT -11.770 -124.205 -10.930 -124.150 ;
        RECT -9.880 -124.240 -7.540 -124.130 ;
        RECT -7.360 -124.205 -6.520 -123.835 ;
        RECT -14.780 -124.360 -14.415 -124.240 ;
        RECT -15.205 -125.435 -15.035 -125.065 ;
        RECT -14.785 -125.200 -14.415 -124.360 ;
        RECT -14.140 -124.280 -11.950 -124.240 ;
        RECT -14.140 -124.605 -13.910 -124.280 ;
        RECT -13.160 -124.605 -12.930 -124.280 ;
        RECT -15.210 -125.660 -15.030 -125.435 ;
        RECT -14.110 -125.565 -13.940 -124.605 ;
        RECT -13.130 -125.565 -12.960 -124.605 ;
        RECT -12.180 -125.545 -11.950 -124.280 ;
        RECT -9.730 -124.280 -7.540 -124.240 ;
        RECT -9.730 -124.605 -9.500 -124.280 ;
        RECT -8.750 -124.605 -8.520 -124.280 ;
        RECT -11.160 -125.455 -10.875 -124.635 ;
        RECT -12.150 -125.565 -11.980 -125.545 ;
        RECT -9.700 -125.565 -9.530 -124.605 ;
        RECT -8.720 -125.565 -8.550 -124.605 ;
        RECT -7.770 -125.545 -7.540 -124.280 ;
        RECT -7.740 -125.565 -7.570 -125.545 ;
        RECT -18.170 -125.830 -15.030 -125.660 ;
        RECT -6.815 -126.950 -6.620 -124.205 ;
        RECT -5.050 -125.480 -4.880 -123.430 ;
        RECT -4.705 -123.200 -4.030 -123.165 ;
        RECT -2.005 -123.200 -1.820 -122.930 ;
        RECT 4.920 -123.050 5.225 -121.015 ;
        RECT 8.620 -121.185 8.795 -120.925 ;
        RECT 7.150 -122.725 7.320 -121.185 ;
        RECT 7.640 -122.725 7.810 -121.185 ;
        RECT 8.130 -122.725 8.300 -121.185 ;
        RECT 8.620 -122.725 8.790 -121.185 ;
        RECT 9.110 -122.725 9.280 -121.185 ;
        RECT 7.010 -122.940 7.380 -122.910 ;
        RECT 9.085 -122.940 9.440 -122.935 ;
        RECT 7.010 -122.945 9.440 -122.940 ;
        RECT -4.705 -123.385 -1.820 -123.200 ;
        RECT -4.705 -123.435 -4.030 -123.385 ;
        RECT -2.005 -124.075 -1.820 -123.385 ;
        RECT -1.650 -123.210 -0.975 -123.175 ;
        RECT -1.650 -123.380 3.130 -123.210 ;
        RECT -1.650 -123.445 -0.975 -123.380 ;
        RECT -0.710 -123.600 -0.035 -123.565 ;
        RECT 2.105 -123.600 2.785 -123.565 ;
        RECT -0.710 -123.790 2.785 -123.600 ;
        RECT -0.710 -123.835 -0.035 -123.790 ;
        RECT 2.105 -123.795 2.785 -123.790 ;
        RECT -2.005 -124.260 0.770 -124.075 ;
        RECT 0.970 -124.245 1.930 -123.975 ;
        RECT 2.960 -124.205 3.130 -123.380 ;
        RECT 3.370 -123.480 6.445 -123.050 ;
        RECT 7.010 -123.135 10.345 -122.945 ;
        RECT 7.010 -123.265 7.380 -123.135 ;
        RECT 9.435 -123.145 10.345 -123.135 ;
        RECT 9.030 -123.415 9.705 -123.385 ;
        RECT 9.030 -123.435 9.855 -123.415 ;
        RECT -1.360 -125.480 -1.190 -124.260 ;
        RECT -0.380 -125.480 -0.210 -124.260 ;
        RECT 0.600 -125.480 0.770 -124.260 ;
        RECT 1.700 -124.665 1.930 -124.245 ;
        RECT 2.930 -124.555 3.785 -124.205 ;
        RECT 4.105 -124.260 4.275 -123.720 ;
        RECT 4.595 -124.260 4.765 -123.480 ;
        RECT 5.085 -124.260 5.255 -123.720 ;
        RECT 5.575 -124.260 5.745 -123.480 ;
        RECT 6.695 -123.540 8.790 -123.500 ;
        RECT 6.640 -123.690 8.790 -123.540 ;
        RECT 9.030 -123.615 9.965 -123.435 ;
        RECT 9.030 -123.655 9.920 -123.615 ;
        RECT 3.615 -125.415 3.785 -124.555 ;
        RECT 5.970 -124.435 6.335 -124.405 ;
        RECT 6.640 -124.435 6.945 -123.690 ;
        RECT 5.970 -124.500 6.945 -124.435 ;
        RECT 5.970 -124.640 6.835 -124.500 ;
        RECT 5.970 -124.705 6.335 -124.640 ;
        RECT 4.595 -125.415 4.765 -124.875 ;
        RECT 5.575 -125.415 5.745 -124.875 ;
        RECT 7.640 -125.410 7.810 -123.690 ;
        RECT 8.620 -125.410 8.790 -123.690 ;
        RECT -6.815 -127.205 -6.130 -126.950 ;
        RECT 9.740 -127.405 9.920 -123.655 ;
        RECT -37.980 -127.680 -37.300 -127.450 ;
        RECT 9.145 -127.635 9.920 -127.405 ;
        RECT -110.180 -134.435 -108.945 -134.430 ;
        RECT -108.135 -134.435 -107.965 -132.580 ;
        RECT -90.945 -132.605 -90.270 -132.575 ;
        RECT -91.045 -132.615 -90.270 -132.605 ;
        RECT -96.355 -132.740 -95.705 -132.655 ;
        RECT -95.485 -132.740 -95.120 -132.675 ;
        RECT -99.030 -132.770 -98.740 -132.765 ;
        RECT -96.355 -132.770 -95.120 -132.740 ;
        RECT -99.030 -132.945 -95.120 -132.770 ;
        RECT -92.080 -132.795 -90.270 -132.615 ;
        RECT -90.030 -132.690 -87.880 -132.540 ;
        RECT -90.030 -132.730 -87.935 -132.690 ;
        RECT -86.985 -132.750 -86.815 -131.970 ;
        RECT -86.495 -132.510 -86.325 -131.970 ;
        RECT -86.005 -132.750 -85.835 -131.970 ;
        RECT -85.515 -132.510 -85.345 -131.970 ;
        RECT -85.025 -132.025 -83.165 -131.675 ;
        RECT -91.045 -132.805 -90.270 -132.795 ;
        RECT -90.945 -132.845 -90.270 -132.805 ;
        RECT -99.030 -133.110 -95.705 -132.945 ;
        RECT -95.485 -132.975 -95.120 -132.945 ;
        RECT -99.030 -133.450 -98.740 -133.110 ;
        RECT -96.355 -133.405 -95.705 -133.110 ;
        RECT -93.420 -133.095 -90.675 -133.085 ;
        RECT -88.620 -133.095 -88.250 -132.965 ;
        RECT -93.420 -133.115 -88.250 -133.095 ;
        RECT -112.210 -134.605 -111.045 -134.435 ;
        RECT -110.180 -134.605 -107.965 -134.435 ;
        RECT -113.930 -134.875 -113.255 -134.840 ;
        RECT -111.230 -134.875 -111.045 -134.605 ;
        RECT -113.930 -135.060 -111.045 -134.875 ;
        RECT -113.930 -135.110 -113.255 -135.060 ;
        RECT -111.230 -135.750 -111.045 -135.060 ;
        RECT -110.875 -134.885 -110.200 -134.850 ;
        RECT -107.730 -134.885 -107.440 -134.370 ;
        RECT -94.895 -134.395 -94.725 -133.115 ;
        RECT -94.405 -134.155 -94.235 -133.115 ;
        RECT -93.915 -134.395 -93.745 -133.115 ;
        RECT -93.425 -133.285 -88.250 -133.115 ;
        RECT -87.685 -133.180 -83.760 -132.750 ;
        RECT -93.425 -134.155 -93.255 -133.285 ;
        RECT -90.680 -133.290 -88.250 -133.285 ;
        RECT -90.680 -133.295 -90.325 -133.290 ;
        RECT -88.620 -133.320 -88.250 -133.290 ;
        RECT -110.875 -135.055 -107.440 -134.885 ;
        RECT -110.875 -135.120 -110.200 -135.055 ;
        RECT -109.935 -135.275 -109.260 -135.240 ;
        RECT -104.080 -135.275 -103.790 -134.780 ;
        RECT -95.595 -134.825 -90.905 -134.395 ;
        RECT -109.935 -135.465 -103.790 -135.275 ;
        RECT -109.935 -135.510 -109.260 -135.465 ;
        RECT -108.255 -135.695 -107.580 -135.650 ;
        RECT -99.455 -135.695 -99.165 -135.210 ;
        RECT -91.335 -135.230 -90.905 -134.825 ;
        RECT -90.520 -135.045 -90.350 -133.505 ;
        RECT -90.030 -135.045 -89.860 -133.505 ;
        RECT -89.540 -135.045 -89.370 -133.505 ;
        RECT -89.050 -135.045 -88.880 -133.505 ;
        RECT -88.560 -135.045 -88.390 -133.505 ;
        RECT -90.035 -135.230 -89.860 -135.045 ;
        RECT -86.465 -135.215 -86.160 -133.180 ;
        RECT -88.410 -135.230 -86.160 -135.215 ;
        RECT -91.335 -135.520 -86.160 -135.230 ;
        RECT -37.780 -135.335 -37.610 -127.680 ;
        RECT -25.580 -128.045 -24.900 -127.815 ;
        RECT 10.145 -127.825 10.345 -123.145 ;
        RECT 10.820 -124.195 11.170 -120.520 ;
        RECT 12.945 -120.700 13.700 -118.310 ;
        RECT 15.155 -120.610 15.910 -118.310 ;
        RECT 16.620 -120.610 17.375 -118.310 ;
        RECT 19.820 -119.680 20.550 -118.310 ;
        RECT 22.045 -119.680 22.775 -118.310 ;
        RECT 23.375 -119.680 24.105 -118.310 ;
        RECT 25.175 -119.680 25.905 -118.310 ;
        RECT 18.330 -119.960 19.010 -119.730 ;
        RECT 15.155 -120.700 17.405 -120.610 ;
        RECT 12.945 -120.915 17.405 -120.700 ;
        RECT 12.945 -121.005 15.195 -120.915 ;
        RECT 12.945 -123.040 13.250 -121.005 ;
        RECT 16.645 -121.175 16.820 -120.915 ;
        RECT 15.175 -122.715 15.345 -121.175 ;
        RECT 15.665 -122.715 15.835 -121.175 ;
        RECT 16.155 -122.715 16.325 -121.175 ;
        RECT 16.645 -122.715 16.815 -121.175 ;
        RECT 17.135 -122.715 17.305 -121.175 ;
        RECT 18.680 -122.235 19.005 -119.960 ;
        RECT 19.700 -120.005 26.070 -119.680 ;
        RECT 19.760 -122.235 19.930 -120.945 ;
        RECT 20.250 -121.985 20.420 -120.005 ;
        RECT 22.315 -120.455 24.520 -120.285 ;
        RECT 18.680 -122.525 19.930 -122.235 ;
        RECT 15.035 -122.930 15.405 -122.900 ;
        RECT 17.110 -122.930 17.465 -122.925 ;
        RECT 15.035 -122.935 17.465 -122.930 ;
        RECT 11.395 -123.470 14.470 -123.040 ;
        RECT 15.035 -123.125 18.485 -122.935 ;
        RECT 15.035 -123.255 15.405 -123.125 ;
        RECT 17.460 -123.135 18.485 -123.125 ;
        RECT 17.055 -123.415 17.730 -123.375 ;
        RECT 17.055 -123.425 17.990 -123.415 ;
        RECT 10.820 -124.545 11.810 -124.195 ;
        RECT 12.130 -124.250 12.300 -123.710 ;
        RECT 12.620 -124.250 12.790 -123.470 ;
        RECT 13.110 -124.250 13.280 -123.710 ;
        RECT 13.600 -124.250 13.770 -123.470 ;
        RECT 14.720 -123.530 16.815 -123.490 ;
        RECT 14.665 -123.680 16.815 -123.530 ;
        RECT 17.055 -123.615 18.090 -123.425 ;
        RECT 17.055 -123.645 17.730 -123.615 ;
        RECT 11.640 -125.405 11.810 -124.545 ;
        RECT 13.995 -124.425 14.360 -124.395 ;
        RECT 14.665 -124.425 14.970 -123.680 ;
        RECT 13.995 -124.490 14.970 -124.425 ;
        RECT 13.995 -124.630 14.860 -124.490 ;
        RECT 13.995 -124.695 14.360 -124.630 ;
        RECT 12.620 -125.405 12.790 -124.865 ;
        RECT 13.600 -125.405 13.770 -124.865 ;
        RECT 15.665 -125.400 15.835 -123.680 ;
        RECT 16.645 -125.400 16.815 -123.680 ;
        RECT -25.580 -129.310 -25.380 -128.045 ;
        RECT 9.665 -128.055 10.345 -127.825 ;
        RECT -25.595 -129.990 -25.365 -129.310 ;
        RECT 17.910 -130.250 18.090 -123.615 ;
        RECT 10.485 -130.430 18.090 -130.250 ;
        RECT 10.485 -130.990 10.665 -130.430 ;
        RECT 18.285 -130.600 18.485 -123.135 ;
        RECT 19.760 -125.525 19.930 -122.525 ;
        RECT 21.825 -122.805 21.995 -120.945 ;
        RECT 22.315 -122.485 22.485 -120.455 ;
        RECT 23.365 -120.470 24.520 -120.455 ;
        RECT 22.805 -122.805 22.975 -120.945 ;
        RECT 23.365 -121.000 23.540 -120.470 ;
        RECT 23.370 -122.485 23.540 -121.000 ;
        RECT 23.860 -122.485 24.030 -120.945 ;
        RECT 24.345 -120.990 24.520 -120.470 ;
        RECT 24.350 -122.485 24.520 -120.990 ;
        RECT 23.855 -122.800 24.030 -122.485 ;
        RECT 24.920 -122.800 25.090 -120.950 ;
        RECT 25.410 -122.490 25.580 -120.005 ;
        RECT 27.995 -120.580 28.980 -118.310 ;
        RECT 30.660 -120.580 31.645 -118.310 ;
        RECT 33.225 -120.535 34.210 -118.310 ;
        RECT 35.740 -120.535 36.725 -118.310 ;
        RECT 37.715 -120.445 39.020 -118.310 ;
        RECT 45.440 -117.995 45.760 -117.880 ;
        RECT 72.265 -117.995 72.680 -117.020 ;
        RECT 76.550 -117.130 77.655 -117.020 ;
        RECT 45.440 -118.410 72.680 -117.995 ;
        RECT 45.440 -118.470 45.760 -118.410 ;
        RECT 91.965 -118.800 92.710 -106.125 ;
        RECT 93.040 -107.560 93.700 -106.885 ;
        RECT 93.040 -109.235 93.570 -107.560 ;
        RECT 94.770 -108.775 95.690 -106.125 ;
        RECT 97.890 -106.295 98.100 -106.075 ;
        RECT 98.405 -106.115 98.575 -105.660 ;
        RECT 98.895 -106.025 99.065 -105.575 ;
        RECT 99.360 -105.685 99.570 -105.405 ;
        RECT 98.890 -106.295 99.070 -106.025 ;
        RECT 99.385 -106.115 99.555 -105.685 ;
        RECT 99.875 -106.025 100.045 -105.575 ;
        RECT 100.330 -105.680 100.540 -105.405 ;
        RECT 99.860 -106.115 100.045 -106.025 ;
        RECT 100.365 -106.115 100.535 -105.680 ;
        RECT 100.855 -106.035 101.025 -105.575 ;
        RECT 101.340 -105.630 101.520 -105.405 ;
        RECT 111.880 -105.405 115.020 -105.235 ;
        RECT 101.345 -106.000 101.515 -105.630 ;
        RECT 99.860 -106.295 100.040 -106.115 ;
        RECT 100.850 -106.295 101.030 -106.035 ;
        RECT 97.890 -106.465 101.030 -106.295 ;
        RECT 97.890 -107.010 98.765 -106.465 ;
        RECT 101.310 -106.735 101.545 -106.000 ;
        RECT 101.765 -106.705 102.135 -105.865 ;
        RECT 102.440 -106.460 102.610 -105.500 ;
        RECT 103.420 -106.460 103.590 -105.500 ;
        RECT 104.400 -105.520 104.570 -105.500 ;
        RECT 97.515 -107.300 98.765 -107.010 ;
        RECT 100.685 -107.105 101.545 -106.735 ;
        RECT 97.515 -107.310 101.045 -107.300 ;
        RECT 97.890 -107.470 101.045 -107.310 ;
        RECT 97.890 -107.505 98.100 -107.470 ;
        RECT 97.895 -107.720 98.100 -107.505 ;
        RECT 97.915 -108.190 98.085 -107.720 ;
        RECT 98.405 -108.130 98.575 -107.650 ;
        RECT 98.880 -107.715 99.085 -107.470 ;
        RECT 98.375 -108.420 98.595 -108.130 ;
        RECT 98.895 -108.190 99.065 -107.715 ;
        RECT 99.385 -108.075 99.555 -107.650 ;
        RECT 99.850 -107.715 100.055 -107.470 ;
        RECT 99.360 -108.420 99.580 -108.075 ;
        RECT 99.875 -108.190 100.045 -107.715 ;
        RECT 100.365 -108.075 100.535 -107.650 ;
        RECT 100.840 -107.675 101.045 -107.470 ;
        RECT 100.340 -108.420 100.560 -108.075 ;
        RECT 100.855 -108.190 101.025 -107.675 ;
        RECT 101.310 -107.780 101.545 -107.105 ;
        RECT 101.770 -106.825 102.135 -106.705 ;
        RECT 102.410 -106.785 102.640 -106.460 ;
        RECT 103.390 -106.785 103.620 -106.460 ;
        RECT 104.370 -106.785 104.600 -105.520 ;
        RECT 105.390 -105.870 105.675 -105.610 ;
        RECT 105.390 -106.180 106.415 -105.870 ;
        RECT 105.390 -106.430 105.675 -106.180 ;
        RECT 102.410 -106.825 104.600 -106.785 ;
        RECT 101.770 -107.015 104.600 -106.825 ;
        RECT 106.105 -106.825 106.415 -106.180 ;
        RECT 106.625 -106.460 106.795 -105.500 ;
        RECT 107.605 -106.460 107.775 -105.500 ;
        RECT 108.585 -105.520 108.755 -105.500 ;
        RECT 106.595 -106.785 106.825 -106.460 ;
        RECT 107.575 -106.785 107.805 -106.460 ;
        RECT 108.555 -106.785 108.785 -105.520 ;
        RECT 111.415 -106.075 111.585 -105.575 ;
        RECT 111.880 -105.660 112.090 -105.405 ;
        RECT 106.595 -106.825 108.785 -106.785 ;
        RECT 101.770 -107.175 102.640 -107.015 ;
        RECT 102.410 -107.480 102.640 -107.175 ;
        RECT 101.345 -108.130 101.515 -107.780 ;
        RECT 102.440 -107.940 102.610 -107.480 ;
        RECT 101.320 -108.420 101.540 -108.130 ;
        RECT 102.930 -108.195 103.100 -107.400 ;
        RECT 103.390 -107.480 103.620 -107.015 ;
        RECT 103.420 -107.940 103.590 -107.480 ;
        RECT 103.910 -108.195 104.080 -107.400 ;
        RECT 104.370 -107.480 104.600 -107.015 ;
        RECT 104.780 -106.915 105.620 -106.860 ;
        RECT 104.780 -107.230 105.920 -106.915 ;
        RECT 106.105 -107.015 108.785 -106.825 ;
        RECT 111.390 -106.295 111.600 -106.075 ;
        RECT 111.905 -106.115 112.075 -105.660 ;
        RECT 112.395 -106.025 112.565 -105.575 ;
        RECT 112.860 -105.685 113.070 -105.405 ;
        RECT 112.390 -106.295 112.570 -106.025 ;
        RECT 112.885 -106.115 113.055 -105.685 ;
        RECT 113.375 -106.025 113.545 -105.575 ;
        RECT 113.830 -105.680 114.040 -105.405 ;
        RECT 113.360 -106.115 113.545 -106.025 ;
        RECT 113.865 -106.115 114.035 -105.680 ;
        RECT 114.355 -106.035 114.525 -105.575 ;
        RECT 114.840 -105.630 115.020 -105.405 ;
        RECT 140.145 -105.420 140.315 -103.700 ;
        RECT 141.125 -105.420 141.295 -103.700 ;
        RECT 141.990 -104.445 142.295 -103.700 ;
        RECT 143.190 -104.270 143.360 -103.490 ;
        RECT 143.680 -104.270 143.850 -103.730 ;
        RECT 144.170 -104.270 144.340 -103.490 ;
        RECT 176.020 -103.555 177.255 -103.350 ;
        RECT 181.430 -103.490 182.105 -103.450 ;
        RECT 181.330 -103.500 182.105 -103.490 ;
        RECT 176.020 -103.640 176.670 -103.555 ;
        RECT 176.890 -103.620 177.255 -103.555 ;
        RECT 180.295 -103.680 182.105 -103.500 ;
        RECT 184.690 -103.545 188.615 -103.115 ;
        RECT 220.335 -103.545 220.985 -103.085 ;
        RECT 221.795 -103.375 221.965 -102.095 ;
        RECT 222.285 -103.375 222.455 -102.335 ;
        RECT 222.775 -103.375 222.945 -102.095 ;
        RECT 223.265 -103.205 223.435 -102.335 ;
        RECT 226.170 -102.985 226.340 -101.445 ;
        RECT 226.660 -102.985 226.830 -101.445 ;
        RECT 227.150 -102.985 227.320 -101.445 ;
        RECT 227.640 -102.985 227.810 -101.445 ;
        RECT 228.130 -102.985 228.300 -101.445 ;
        RECT 226.010 -103.200 226.365 -103.195 ;
        RECT 228.070 -103.200 228.440 -103.170 ;
        RECT 226.010 -103.205 228.440 -103.200 ;
        RECT 223.265 -103.375 228.440 -103.205 ;
        RECT 230.225 -103.310 230.530 -101.275 ;
        RECT 254.000 -101.115 255.130 -101.070 ;
        RECT 262.265 -101.115 263.495 -100.715 ;
        RECT 254.000 -101.780 263.495 -101.115 ;
        RECT 271.345 -100.800 274.670 -100.660 ;
        RECT 271.345 -101.090 276.520 -100.800 ;
        RECT 271.345 -101.495 271.775 -101.090 ;
        RECT 272.645 -101.275 272.820 -101.090 ;
        RECT 274.270 -101.105 276.520 -101.090 ;
        RECT 254.000 -102.240 255.130 -101.780 ;
        RECT 262.265 -101.815 263.495 -101.780 ;
        RECT 267.085 -101.925 271.775 -101.495 ;
        RECT 223.270 -103.395 228.440 -103.375 ;
        RECT 223.270 -103.405 226.015 -103.395 ;
        RECT 221.205 -103.545 221.570 -103.515 ;
        RECT 228.070 -103.525 228.440 -103.395 ;
        RECT 181.330 -103.690 182.105 -103.680 ;
        RECT 181.430 -103.720 182.105 -103.690 ;
        RECT 182.345 -103.605 184.440 -103.565 ;
        RECT 144.660 -104.270 144.830 -103.730 ;
        RECT 182.345 -103.755 184.495 -103.605 ;
        RECT 142.600 -104.445 142.965 -104.415 ;
        RECT 141.990 -104.510 142.965 -104.445 ;
        RECT 142.100 -104.650 142.965 -104.510 ;
        RECT 142.600 -104.715 142.965 -104.650 ;
        RECT 145.150 -104.565 147.010 -104.215 ;
        RECT 143.190 -105.425 143.360 -104.885 ;
        RECT 144.170 -105.425 144.340 -104.885 ;
        RECT 145.150 -105.425 145.320 -104.565 ;
        RECT 114.845 -106.000 115.015 -105.630 ;
        RECT 113.360 -106.295 113.540 -106.115 ;
        RECT 114.350 -106.295 114.530 -106.035 ;
        RECT 111.390 -106.465 114.530 -106.295 ;
        RECT 106.105 -107.175 106.825 -107.015 ;
        RECT 104.400 -107.940 104.570 -107.480 ;
        RECT 104.890 -108.195 105.060 -107.400 ;
        RECT 105.620 -108.025 105.920 -107.230 ;
        RECT 106.595 -107.480 106.825 -107.175 ;
        RECT 106.625 -107.940 106.795 -107.480 ;
        RECT 107.115 -108.195 107.285 -107.400 ;
        RECT 107.575 -107.480 107.805 -107.015 ;
        RECT 107.605 -107.940 107.775 -107.480 ;
        RECT 108.095 -108.195 108.265 -107.400 ;
        RECT 108.555 -107.480 108.785 -107.015 ;
        RECT 108.965 -106.895 109.805 -106.860 ;
        RECT 108.965 -107.195 109.915 -106.895 ;
        RECT 111.390 -107.000 112.265 -106.465 ;
        RECT 114.810 -106.735 115.045 -106.000 ;
        RECT 115.265 -106.705 115.635 -105.865 ;
        RECT 115.940 -106.460 116.110 -105.500 ;
        RECT 116.920 -106.460 117.090 -105.500 ;
        RECT 117.900 -105.520 118.070 -105.500 ;
        RECT 108.965 -107.230 109.805 -107.195 ;
        RECT 110.935 -107.300 112.265 -107.000 ;
        RECT 114.185 -107.105 115.045 -106.735 ;
        RECT 108.585 -107.940 108.755 -107.480 ;
        RECT 109.075 -108.195 109.245 -107.400 ;
        RECT 111.390 -107.470 114.545 -107.300 ;
        RECT 111.390 -107.505 111.600 -107.470 ;
        RECT 111.395 -107.720 111.600 -107.505 ;
        RECT 111.415 -108.190 111.585 -107.720 ;
        RECT 111.905 -108.130 112.075 -107.650 ;
        RECT 112.380 -107.715 112.585 -107.470 ;
        RECT 98.375 -108.590 101.540 -108.420 ;
        RECT 102.435 -108.205 105.105 -108.195 ;
        RECT 106.620 -108.205 109.290 -108.195 ;
        RECT 102.435 -108.535 109.290 -108.205 ;
        RECT 111.875 -108.420 112.095 -108.130 ;
        RECT 112.395 -108.190 112.565 -107.715 ;
        RECT 112.885 -108.075 113.055 -107.650 ;
        RECT 113.350 -107.715 113.555 -107.470 ;
        RECT 112.860 -108.420 113.080 -108.075 ;
        RECT 113.375 -108.190 113.545 -107.715 ;
        RECT 113.865 -108.075 114.035 -107.650 ;
        RECT 114.340 -107.675 114.545 -107.470 ;
        RECT 113.840 -108.420 114.060 -108.075 ;
        RECT 114.355 -108.190 114.525 -107.675 ;
        RECT 114.810 -107.780 115.045 -107.105 ;
        RECT 115.270 -106.825 115.635 -106.705 ;
        RECT 115.910 -106.785 116.140 -106.460 ;
        RECT 116.890 -106.785 117.120 -106.460 ;
        RECT 117.870 -106.785 118.100 -105.520 ;
        RECT 118.890 -105.930 119.175 -105.610 ;
        RECT 118.890 -106.175 119.890 -105.930 ;
        RECT 118.890 -106.430 119.175 -106.175 ;
        RECT 115.910 -106.825 118.100 -106.785 ;
        RECT 115.270 -107.015 118.100 -106.825 ;
        RECT 119.660 -106.825 119.890 -106.175 ;
        RECT 120.125 -106.460 120.295 -105.500 ;
        RECT 121.105 -106.460 121.275 -105.500 ;
        RECT 122.085 -105.520 122.255 -105.500 ;
        RECT 120.095 -106.785 120.325 -106.460 ;
        RECT 121.075 -106.785 121.305 -106.460 ;
        RECT 122.055 -106.785 122.285 -105.520 ;
        RECT 120.095 -106.825 122.285 -106.785 ;
        RECT 115.270 -107.175 116.140 -107.015 ;
        RECT 115.910 -107.480 116.140 -107.175 ;
        RECT 114.845 -108.130 115.015 -107.780 ;
        RECT 115.940 -107.940 116.110 -107.480 ;
        RECT 114.820 -108.420 115.040 -108.130 ;
        RECT 116.430 -108.195 116.600 -107.400 ;
        RECT 116.890 -107.480 117.120 -107.015 ;
        RECT 116.920 -107.940 117.090 -107.480 ;
        RECT 117.410 -108.195 117.580 -107.400 ;
        RECT 117.870 -107.480 118.100 -107.015 ;
        RECT 118.280 -106.915 119.120 -106.860 ;
        RECT 118.280 -106.920 119.295 -106.915 ;
        RECT 118.280 -107.230 119.480 -106.920 ;
        RECT 119.660 -107.015 122.285 -106.825 ;
        RECT 119.660 -107.175 120.325 -107.015 ;
        RECT 117.900 -107.940 118.070 -107.480 ;
        RECT 118.390 -108.195 118.560 -107.400 ;
        RECT 119.180 -107.950 119.480 -107.230 ;
        RECT 120.095 -107.480 120.325 -107.175 ;
        RECT 120.125 -107.940 120.295 -107.480 ;
        RECT 120.615 -108.195 120.785 -107.400 ;
        RECT 121.075 -107.480 121.305 -107.015 ;
        RECT 121.105 -107.940 121.275 -107.480 ;
        RECT 121.595 -108.195 121.765 -107.400 ;
        RECT 122.055 -107.480 122.285 -107.015 ;
        RECT 122.465 -107.010 123.305 -106.860 ;
        RECT 122.465 -107.230 123.340 -107.010 ;
        RECT 122.085 -107.940 122.255 -107.480 ;
        RECT 122.575 -108.195 122.745 -107.400 ;
        RECT 103.560 -108.775 104.115 -108.535 ;
        RECT 104.990 -108.545 107.590 -108.535 ;
        RECT 107.950 -108.765 108.505 -108.535 ;
        RECT 111.875 -108.590 115.040 -108.420 ;
        RECT 115.935 -108.535 122.790 -108.195 ;
        RECT 107.935 -108.775 108.620 -108.765 ;
        RECT 116.940 -108.775 117.495 -108.535 ;
        RECT 120.995 -108.735 121.550 -108.535 ;
        RECT 120.920 -108.775 121.605 -108.735 ;
        RECT 94.765 -108.970 121.690 -108.775 ;
        RECT 94.770 -109.065 95.430 -108.970 ;
        RECT 107.935 -109.065 108.620 -108.970 ;
        RECT 120.920 -109.035 121.605 -108.970 ;
        RECT 123.100 -109.090 123.340 -107.230 ;
        RECT 143.420 -107.765 144.620 -107.595 ;
        RECT 105.405 -109.235 106.065 -109.185 ;
        RECT 110.110 -109.235 110.795 -109.180 ;
        RECT 93.040 -109.430 121.690 -109.235 ;
        RECT 93.040 -111.400 93.235 -109.430 ;
        RECT 105.405 -109.485 106.065 -109.430 ;
        RECT 110.110 -109.480 110.795 -109.430 ;
        RECT 96.385 -109.665 97.045 -109.615 ;
        RECT 119.000 -109.665 119.660 -109.625 ;
        RECT 96.385 -109.860 121.690 -109.665 ;
        RECT 123.045 -109.775 123.345 -109.090 ;
        RECT 130.990 -109.620 132.285 -109.405 ;
        RECT 96.385 -109.915 97.045 -109.860 ;
        RECT 119.000 -109.925 119.660 -109.860 ;
        RECT 93.455 -110.435 100.535 -110.095 ;
        RECT 101.430 -110.210 104.595 -110.040 ;
        RECT 93.500 -111.230 93.670 -110.435 ;
        RECT 93.990 -111.150 94.160 -110.690 ;
        RECT 92.940 -111.770 93.780 -111.400 ;
        RECT 93.960 -111.615 94.190 -111.150 ;
        RECT 94.480 -111.230 94.650 -110.435 ;
        RECT 94.970 -111.150 95.140 -110.690 ;
        RECT 94.940 -111.615 95.170 -111.150 ;
        RECT 95.460 -111.230 95.630 -110.435 ;
        RECT 95.950 -111.150 96.120 -110.690 ;
        RECT 95.920 -111.455 96.150 -111.150 ;
        RECT 95.920 -111.485 96.300 -111.455 ;
        RECT 96.590 -111.485 96.890 -111.055 ;
        RECT 97.910 -111.230 98.080 -110.435 ;
        RECT 98.400 -111.150 98.570 -110.690 ;
        RECT 97.350 -111.425 98.190 -111.400 ;
        RECT 97.175 -111.485 98.190 -111.425 ;
        RECT 95.920 -111.615 98.190 -111.485 ;
        RECT 93.960 -111.695 98.190 -111.615 ;
        RECT 93.960 -111.805 96.300 -111.695 ;
        RECT 96.590 -111.715 96.890 -111.695 ;
        RECT 97.175 -111.715 98.190 -111.695 ;
        RECT 97.350 -111.770 98.190 -111.715 ;
        RECT 98.370 -111.615 98.600 -111.150 ;
        RECT 98.890 -111.230 99.060 -110.435 ;
        RECT 99.380 -111.150 99.550 -110.690 ;
        RECT 99.350 -111.615 99.580 -111.150 ;
        RECT 99.870 -111.230 100.040 -110.435 ;
        RECT 101.430 -110.500 101.650 -110.210 ;
        RECT 100.360 -111.150 100.530 -110.690 ;
        RECT 101.455 -110.850 101.625 -110.500 ;
        RECT 100.330 -111.455 100.560 -111.150 ;
        RECT 100.330 -111.615 101.200 -111.455 ;
        RECT 98.370 -111.805 101.200 -111.615 ;
        RECT 93.960 -111.845 96.150 -111.805 ;
        RECT 93.960 -113.110 94.190 -111.845 ;
        RECT 94.940 -112.170 95.170 -111.845 ;
        RECT 95.920 -112.170 96.150 -111.845 ;
        RECT 98.370 -111.845 100.560 -111.805 ;
        RECT 93.990 -113.130 94.160 -113.110 ;
        RECT 94.970 -113.130 95.140 -112.170 ;
        RECT 95.950 -113.130 96.120 -112.170 ;
        RECT 97.295 -113.020 97.580 -112.200 ;
        RECT 98.370 -113.110 98.600 -111.845 ;
        RECT 99.350 -112.170 99.580 -111.845 ;
        RECT 100.330 -112.170 100.560 -111.845 ;
        RECT 100.835 -111.925 101.200 -111.805 ;
        RECT 101.425 -111.525 101.660 -110.850 ;
        RECT 101.945 -110.955 102.115 -110.440 ;
        RECT 102.410 -110.555 102.630 -110.210 ;
        RECT 101.925 -111.160 102.130 -110.955 ;
        RECT 102.435 -110.980 102.605 -110.555 ;
        RECT 102.925 -110.915 103.095 -110.440 ;
        RECT 103.390 -110.555 103.610 -110.210 ;
        RECT 102.915 -111.160 103.120 -110.915 ;
        RECT 103.415 -110.980 103.585 -110.555 ;
        RECT 103.905 -110.915 104.075 -110.440 ;
        RECT 104.375 -110.500 104.595 -110.210 ;
        RECT 103.885 -111.160 104.090 -110.915 ;
        RECT 104.395 -110.980 104.565 -110.500 ;
        RECT 104.840 -110.910 105.070 -110.300 ;
        RECT 106.580 -110.435 114.035 -110.095 ;
        RECT 114.930 -110.210 118.095 -110.040 ;
        RECT 104.840 -110.960 105.075 -110.910 ;
        RECT 104.870 -111.125 105.075 -110.960 ;
        RECT 104.870 -111.160 105.080 -111.125 ;
        RECT 101.925 -111.330 105.080 -111.160 ;
        RECT 106.625 -111.230 106.795 -110.435 ;
        RECT 107.115 -111.150 107.285 -110.690 ;
        RECT 104.205 -111.440 105.080 -111.330 ;
        RECT 106.065 -111.440 106.905 -111.400 ;
        RECT 101.425 -111.895 102.285 -111.525 ;
        RECT 104.205 -111.725 106.905 -111.440 ;
        RECT 98.400 -113.130 98.570 -113.110 ;
        RECT 99.380 -113.130 99.550 -112.170 ;
        RECT 100.360 -113.130 100.530 -112.170 ;
        RECT 100.835 -112.765 101.205 -111.925 ;
        RECT 101.425 -112.630 101.660 -111.895 ;
        RECT 104.205 -112.165 105.080 -111.725 ;
        RECT 106.065 -111.770 106.905 -111.725 ;
        RECT 107.085 -111.615 107.315 -111.150 ;
        RECT 107.605 -111.230 107.775 -110.435 ;
        RECT 108.095 -111.150 108.265 -110.690 ;
        RECT 108.065 -111.615 108.295 -111.150 ;
        RECT 108.585 -111.230 108.755 -110.435 ;
        RECT 109.075 -111.150 109.245 -110.690 ;
        RECT 109.045 -111.455 109.275 -111.150 ;
        RECT 109.045 -111.510 109.425 -111.455 ;
        RECT 109.675 -111.510 109.975 -110.935 ;
        RECT 110.250 -111.425 110.550 -111.060 ;
        RECT 111.410 -111.230 111.580 -110.435 ;
        RECT 111.900 -111.150 112.070 -110.690 ;
        RECT 110.850 -111.425 111.690 -111.400 ;
        RECT 109.045 -111.615 110.000 -111.510 ;
        RECT 107.085 -111.735 110.000 -111.615 ;
        RECT 110.250 -111.715 111.690 -111.425 ;
        RECT 110.250 -111.720 110.550 -111.715 ;
        RECT 101.940 -112.335 105.080 -112.165 ;
        RECT 101.940 -112.595 102.120 -112.335 ;
        RECT 102.930 -112.515 103.110 -112.335 ;
        RECT 101.455 -113.000 101.625 -112.630 ;
        RECT 101.450 -113.225 101.630 -113.000 ;
        RECT 101.945 -113.055 102.115 -112.595 ;
        RECT 102.435 -112.950 102.605 -112.515 ;
        RECT 102.925 -112.605 103.110 -112.515 ;
        RECT 102.430 -113.225 102.640 -112.950 ;
        RECT 102.925 -113.055 103.095 -112.605 ;
        RECT 103.415 -112.945 103.585 -112.515 ;
        RECT 103.900 -112.605 104.080 -112.335 ;
        RECT 103.400 -113.225 103.610 -112.945 ;
        RECT 103.905 -113.055 104.075 -112.605 ;
        RECT 104.395 -112.970 104.565 -112.515 ;
        RECT 104.870 -112.555 105.080 -112.335 ;
        RECT 107.085 -111.805 109.425 -111.735 ;
        RECT 107.085 -111.845 109.275 -111.805 ;
        RECT 104.380 -113.225 104.590 -112.970 ;
        RECT 104.885 -113.055 105.055 -112.555 ;
        RECT 107.085 -113.110 107.315 -111.845 ;
        RECT 108.065 -112.170 108.295 -111.845 ;
        RECT 109.045 -112.170 109.275 -111.845 ;
        RECT 107.115 -113.130 107.285 -113.110 ;
        RECT 108.095 -113.130 108.265 -112.170 ;
        RECT 109.075 -113.130 109.245 -112.170 ;
        RECT 109.775 -112.405 110.000 -111.735 ;
        RECT 110.850 -111.770 111.690 -111.715 ;
        RECT 111.870 -111.615 112.100 -111.150 ;
        RECT 112.390 -111.230 112.560 -110.435 ;
        RECT 112.880 -111.150 113.050 -110.690 ;
        RECT 112.850 -111.615 113.080 -111.150 ;
        RECT 113.370 -111.230 113.540 -110.435 ;
        RECT 114.930 -110.500 115.150 -110.210 ;
        RECT 113.860 -111.150 114.030 -110.690 ;
        RECT 114.955 -110.850 115.125 -110.500 ;
        RECT 113.830 -111.455 114.060 -111.150 ;
        RECT 113.830 -111.615 114.700 -111.455 ;
        RECT 111.870 -111.805 114.700 -111.615 ;
        RECT 111.870 -111.845 114.060 -111.805 ;
        RECT 110.795 -112.405 111.080 -112.200 ;
        RECT 109.775 -112.630 111.080 -112.405 ;
        RECT 110.795 -113.020 111.080 -112.630 ;
        RECT 111.870 -113.110 112.100 -111.845 ;
        RECT 112.850 -112.170 113.080 -111.845 ;
        RECT 113.830 -112.170 114.060 -111.845 ;
        RECT 114.335 -111.925 114.700 -111.805 ;
        RECT 114.925 -111.525 115.160 -110.850 ;
        RECT 115.445 -110.955 115.615 -110.440 ;
        RECT 115.910 -110.555 116.130 -110.210 ;
        RECT 115.425 -111.160 115.630 -110.955 ;
        RECT 115.935 -110.980 116.105 -110.555 ;
        RECT 116.425 -110.915 116.595 -110.440 ;
        RECT 116.890 -110.555 117.110 -110.210 ;
        RECT 116.415 -111.160 116.620 -110.915 ;
        RECT 116.915 -110.980 117.085 -110.555 ;
        RECT 117.405 -110.915 117.575 -110.440 ;
        RECT 117.875 -110.500 118.095 -110.210 ;
        RECT 120.080 -110.435 122.750 -110.095 ;
        RECT 117.385 -111.160 117.590 -110.915 ;
        RECT 117.895 -110.980 118.065 -110.500 ;
        RECT 118.385 -110.910 118.555 -110.440 ;
        RECT 118.370 -111.125 118.575 -110.910 ;
        RECT 118.370 -111.160 118.580 -111.125 ;
        RECT 115.425 -111.330 118.580 -111.160 ;
        RECT 120.125 -111.230 120.295 -110.435 ;
        RECT 120.615 -111.150 120.785 -110.690 ;
        RECT 117.705 -111.475 118.580 -111.330 ;
        RECT 119.565 -111.475 120.405 -111.400 ;
        RECT 114.925 -111.895 115.785 -111.525 ;
        RECT 117.705 -111.740 120.405 -111.475 ;
        RECT 111.900 -113.130 112.070 -113.110 ;
        RECT 112.880 -113.130 113.050 -112.170 ;
        RECT 113.860 -113.130 114.030 -112.170 ;
        RECT 114.335 -112.765 114.705 -111.925 ;
        RECT 114.925 -112.630 115.160 -111.895 ;
        RECT 117.705 -112.165 118.580 -111.740 ;
        RECT 119.565 -111.770 120.405 -111.740 ;
        RECT 120.585 -111.615 120.815 -111.150 ;
        RECT 121.105 -111.230 121.275 -110.435 ;
        RECT 121.595 -111.150 121.765 -110.690 ;
        RECT 121.565 -111.615 121.795 -111.150 ;
        RECT 122.085 -111.230 122.255 -110.435 ;
        RECT 122.575 -111.150 122.745 -110.690 ;
        RECT 122.545 -111.455 122.775 -111.150 ;
        RECT 122.545 -111.565 122.925 -111.455 ;
        RECT 123.100 -111.565 123.340 -109.775 ;
        RECT 126.660 -110.175 132.285 -109.620 ;
        RECT 135.150 -110.100 135.320 -108.380 ;
        RECT 136.130 -110.100 136.300 -108.380 ;
        RECT 138.195 -108.915 138.365 -108.375 ;
        RECT 139.175 -108.915 139.345 -108.375 ;
        RECT 137.605 -109.150 137.970 -109.085 ;
        RECT 137.105 -109.290 137.970 -109.150 ;
        RECT 136.995 -109.355 137.970 -109.290 ;
        RECT 136.995 -110.100 137.300 -109.355 ;
        RECT 137.605 -109.385 137.970 -109.355 ;
        RECT 140.155 -109.235 140.325 -108.375 ;
        RECT 134.235 -110.165 134.910 -110.135 ;
        RECT 134.135 -110.175 134.910 -110.165 ;
        RECT 126.660 -110.355 134.910 -110.175 ;
        RECT 135.150 -110.250 137.300 -110.100 ;
        RECT 135.150 -110.290 137.245 -110.250 ;
        RECT 138.195 -110.310 138.365 -109.530 ;
        RECT 138.685 -110.070 138.855 -109.530 ;
        RECT 139.175 -110.310 139.345 -109.530 ;
        RECT 139.665 -110.070 139.835 -109.530 ;
        RECT 140.155 -109.585 141.545 -109.235 ;
        RECT 126.660 -110.645 132.285 -110.355 ;
        RECT 134.135 -110.365 134.910 -110.355 ;
        RECT 134.235 -110.405 134.910 -110.365 ;
        RECT 130.990 -110.720 132.285 -110.645 ;
        RECT 133.370 -110.655 134.505 -110.645 ;
        RECT 136.560 -110.655 136.930 -110.525 ;
        RECT 133.370 -110.845 136.930 -110.655 ;
        RECT 137.495 -110.740 140.570 -110.310 ;
        RECT 122.545 -111.615 123.340 -111.565 ;
        RECT 120.585 -111.750 123.340 -111.615 ;
        RECT 120.585 -111.760 123.335 -111.750 ;
        RECT 115.440 -112.335 118.580 -112.165 ;
        RECT 115.440 -112.595 115.620 -112.335 ;
        RECT 116.430 -112.515 116.610 -112.335 ;
        RECT 114.955 -113.000 115.125 -112.630 ;
        RECT 101.450 -113.395 104.590 -113.225 ;
        RECT 114.950 -113.225 115.130 -113.000 ;
        RECT 115.445 -113.055 115.615 -112.595 ;
        RECT 115.935 -112.950 116.105 -112.515 ;
        RECT 116.425 -112.605 116.610 -112.515 ;
        RECT 115.930 -113.225 116.140 -112.950 ;
        RECT 116.425 -113.055 116.595 -112.605 ;
        RECT 116.915 -112.945 117.085 -112.515 ;
        RECT 117.400 -112.605 117.580 -112.335 ;
        RECT 116.900 -113.225 117.110 -112.945 ;
        RECT 117.405 -113.055 117.575 -112.605 ;
        RECT 117.895 -112.970 118.065 -112.515 ;
        RECT 118.370 -112.555 118.580 -112.335 ;
        RECT 120.585 -111.805 122.925 -111.760 ;
        RECT 120.585 -111.845 122.775 -111.805 ;
        RECT 117.880 -113.225 118.090 -112.970 ;
        RECT 118.385 -113.055 118.555 -112.555 ;
        RECT 120.585 -113.110 120.815 -111.845 ;
        RECT 121.565 -112.170 121.795 -111.845 ;
        RECT 122.545 -112.170 122.775 -111.845 ;
        RECT 120.615 -113.130 120.785 -113.110 ;
        RECT 121.595 -113.130 121.765 -112.170 ;
        RECT 122.575 -113.130 122.745 -112.170 ;
        RECT 114.950 -113.395 118.090 -113.225 ;
        RECT 103.615 -114.900 104.415 -114.240 ;
        RECT 103.650 -115.815 104.325 -114.900 ;
        RECT 108.405 -115.510 123.025 -115.025 ;
        RECT 103.600 -116.475 104.400 -115.815 ;
        RECT 106.215 -118.070 106.385 -115.850 ;
        RECT 107.195 -118.070 107.365 -115.850 ;
        RECT 106.215 -118.075 107.365 -118.070 ;
        RECT 103.085 -118.140 103.745 -118.090 ;
        RECT 105.300 -118.135 105.975 -118.105 ;
        RECT 105.200 -118.140 105.975 -118.135 ;
        RECT 103.085 -118.320 105.975 -118.140 ;
        RECT 106.215 -118.260 107.435 -118.075 ;
        RECT 103.085 -118.390 103.745 -118.320 ;
        RECT 105.200 -118.335 105.975 -118.320 ;
        RECT 105.300 -118.375 105.975 -118.335 ;
        RECT 107.265 -118.435 107.435 -118.260 ;
        RECT 107.915 -118.435 108.215 -118.135 ;
        RECT 95.940 -118.800 103.920 -118.585 ;
        RECT 86.695 -118.910 103.920 -118.800 ;
        RECT 104.850 -118.600 105.645 -118.595 ;
        RECT 104.850 -118.625 105.650 -118.600 ;
        RECT 106.390 -118.625 107.065 -118.595 ;
        RECT 104.850 -118.820 107.065 -118.625 ;
        RECT 104.850 -118.825 105.920 -118.820 ;
        RECT 104.850 -118.890 105.650 -118.825 ;
        RECT 106.390 -118.865 107.065 -118.820 ;
        RECT 107.265 -118.740 108.215 -118.435 ;
        RECT 104.850 -118.895 105.645 -118.890 ;
        RECT 86.695 -119.245 96.840 -118.910 ;
        RECT 43.835 -119.515 44.130 -119.480 ;
        RECT 43.835 -119.930 63.715 -119.515 ;
        RECT 43.835 -119.955 44.130 -119.930 ;
        RECT 33.225 -120.580 36.970 -120.535 ;
        RECT 27.805 -120.845 36.970 -120.580 ;
        RECT 23.855 -122.805 25.090 -122.800 ;
        RECT 25.900 -122.805 26.070 -120.950 ;
        RECT 27.805 -121.460 28.000 -120.845 ;
        RECT 33.810 -121.015 36.970 -120.845 ;
        RECT 28.315 -121.215 33.355 -121.035 ;
        RECT 27.825 -122.405 27.995 -121.460 ;
        RECT 21.825 -122.975 22.990 -122.805 ;
        RECT 23.855 -122.975 26.070 -122.805 ;
        RECT 27.815 -122.820 28.000 -122.405 ;
        RECT 28.315 -122.440 28.485 -121.215 ;
        RECT 29.895 -122.410 30.065 -121.400 ;
        RECT 30.385 -122.395 30.555 -121.400 ;
        RECT 31.705 -122.395 31.875 -121.400 ;
        RECT 29.880 -122.515 30.065 -122.410 ;
        RECT 29.285 -122.700 30.065 -122.515 ;
        RECT 30.375 -122.590 31.875 -122.395 ;
        RECT 29.285 -122.820 29.470 -122.700 ;
        RECT 20.105 -123.245 20.780 -123.210 ;
        RECT 22.805 -123.245 22.990 -122.975 ;
        RECT 27.815 -123.005 29.470 -122.820 ;
        RECT 32.195 -122.855 32.365 -121.400 ;
        RECT 33.175 -121.485 33.355 -121.215 ;
        RECT 33.175 -122.440 33.345 -121.485 ;
        RECT 33.665 -122.855 33.835 -121.400 ;
        RECT 34.725 -122.355 34.895 -121.400 ;
        RECT 35.190 -121.435 35.405 -121.015 ;
        RECT 34.700 -122.580 34.915 -122.355 ;
        RECT 35.215 -122.440 35.385 -121.435 ;
        RECT 36.270 -122.345 36.440 -121.400 ;
        RECT 36.735 -121.445 36.950 -121.015 ;
        RECT 34.220 -122.810 34.915 -122.580 ;
        RECT 31.030 -123.025 33.835 -122.855 ;
        RECT 20.105 -123.430 22.990 -123.245 ;
        RECT 20.105 -123.480 20.780 -123.430 ;
        RECT 22.805 -124.120 22.990 -123.430 ;
        RECT 23.160 -123.255 23.835 -123.220 ;
        RECT 23.160 -123.425 27.255 -123.255 ;
        RECT 31.030 -123.335 31.200 -123.025 ;
        RECT 23.160 -123.490 23.835 -123.425 ;
        RECT 24.100 -123.645 24.775 -123.610 ;
        RECT 24.100 -123.835 26.905 -123.645 ;
        RECT 24.100 -123.880 24.775 -123.835 ;
        RECT 25.775 -124.065 26.455 -124.020 ;
        RECT 22.805 -124.305 25.580 -124.120 ;
        RECT 25.775 -124.250 26.550 -124.065 ;
        RECT 25.780 -124.290 26.455 -124.250 ;
        RECT 23.450 -125.525 23.620 -124.305 ;
        RECT 24.430 -125.525 24.600 -124.305 ;
        RECT 25.410 -125.525 25.580 -124.305 ;
        RECT -11.595 -131.170 10.665 -130.990 ;
        RECT 10.975 -130.770 18.485 -130.600 ;
        RECT 26.735 -130.680 26.905 -123.835 ;
        RECT -11.595 -131.410 -11.350 -131.170 ;
        RECT 0.455 -131.390 1.135 -131.345 ;
        RECT 10.975 -131.390 11.145 -130.770 ;
        RECT 25.205 -130.850 26.905 -130.680 ;
        RECT 11.370 -131.045 12.050 -131.030 ;
        RECT 25.205 -131.045 25.375 -130.850 ;
        RECT 11.370 -131.215 25.375 -131.045 ;
        RECT 25.895 -131.140 26.575 -131.110 ;
        RECT 27.085 -131.140 27.255 -123.425 ;
        RECT 27.820 -123.680 28.515 -123.410 ;
        RECT 30.470 -123.505 31.200 -123.335 ;
        RECT 30.470 -124.080 30.640 -123.505 ;
        RECT 31.565 -123.530 32.260 -123.260 ;
        RECT 27.570 -124.250 30.640 -124.080 ;
        RECT 30.945 -123.885 33.345 -123.715 ;
        RECT 27.825 -125.990 27.995 -124.430 ;
        RECT 28.315 -125.470 28.485 -124.250 ;
        RECT 28.805 -125.990 28.975 -124.430 ;
        RECT 29.405 -125.645 29.575 -124.430 ;
        RECT 29.895 -125.470 30.065 -124.250 ;
        RECT 30.385 -125.645 30.555 -124.430 ;
        RECT 30.945 -125.645 31.115 -123.885 ;
        RECT 29.405 -125.815 31.115 -125.645 ;
        RECT 31.295 -124.255 32.365 -124.085 ;
        RECT 31.295 -125.990 31.465 -124.255 ;
        RECT 32.195 -125.470 32.365 -124.255 ;
        RECT 33.175 -125.470 33.345 -123.885 ;
        RECT 33.610 -123.900 34.305 -123.630 ;
        RECT 34.700 -124.505 34.915 -122.810 ;
        RECT 36.250 -123.300 36.465 -122.345 ;
        RECT 36.760 -122.440 36.930 -121.445 ;
        RECT 37.715 -121.750 43.490 -120.445 ;
        RECT 60.400 -120.875 61.825 -120.585 ;
        RECT 63.300 -120.875 63.715 -119.930 ;
        RECT 87.340 -120.005 87.560 -119.245 ;
        RECT 87.360 -120.800 87.530 -120.005 ;
        RECT 87.850 -120.755 88.020 -119.760 ;
        RECT 88.310 -120.000 88.530 -119.245 ;
        RECT 60.400 -121.015 85.200 -120.875 ;
        RECT 86.890 -121.015 87.620 -120.975 ;
        RECT 60.400 -121.195 87.620 -121.015 ;
        RECT 87.825 -121.000 88.050 -120.755 ;
        RECT 88.340 -120.800 88.510 -120.000 ;
        RECT 92.070 -120.005 92.290 -119.245 ;
        RECT 92.090 -120.800 92.260 -120.005 ;
        RECT 92.580 -120.755 92.750 -119.760 ;
        RECT 93.040 -120.000 93.260 -119.245 ;
        RECT 87.825 -121.005 89.795 -121.000 ;
        RECT 87.825 -121.180 90.040 -121.005 ;
        RECT 91.620 -121.015 92.350 -120.975 ;
        RECT 60.400 -121.345 85.200 -121.195 ;
        RECT 86.890 -121.275 87.620 -121.195 ;
        RECT 89.100 -121.225 90.040 -121.180 ;
        RECT 91.325 -121.195 92.350 -121.015 ;
        RECT 92.555 -121.000 92.780 -120.755 ;
        RECT 93.070 -120.800 93.240 -120.000 ;
        RECT 92.555 -121.180 95.905 -121.000 ;
        RECT 89.380 -121.305 90.040 -121.225 ;
        RECT 91.620 -121.275 92.350 -121.195 ;
        RECT 93.830 -121.225 95.905 -121.180 ;
        RECT 60.400 -121.680 61.825 -121.345 ;
        RECT 88.005 -121.460 88.720 -121.375 ;
        RECT 85.715 -121.640 88.720 -121.460 ;
        RECT 35.750 -123.530 36.465 -123.300 ;
        RECT 34.725 -125.470 34.895 -124.505 ;
        RECT 36.250 -124.515 36.465 -123.530 ;
        RECT 36.685 -123.870 37.380 -123.600 ;
        RECT 36.270 -125.470 36.440 -124.515 ;
        RECT 27.825 -126.160 31.465 -125.990 ;
        RECT 11.370 -131.260 12.050 -131.215 ;
        RECT 25.895 -131.310 27.255 -131.140 ;
        RECT 25.895 -131.340 26.575 -131.310 ;
        RECT -12.030 -131.640 -11.350 -131.410 ;
        RECT 0.290 -131.560 11.145 -131.390 ;
        RECT 0.455 -131.575 1.135 -131.560 ;
        RECT 37.715 -131.725 39.020 -121.750 ;
        RECT 42.185 -125.720 43.490 -121.750 ;
        RECT 85.715 -121.905 85.895 -121.640 ;
        RECT 88.005 -121.675 88.720 -121.640 ;
        RECT 65.310 -122.715 85.895 -121.905 ;
        RECT 87.355 -122.050 89.095 -121.870 ;
        RECT 87.355 -122.245 87.535 -122.050 ;
        RECT 44.600 -123.530 44.945 -123.440 ;
        RECT 70.665 -123.530 71.220 -122.715 ;
        RECT 44.600 -124.085 71.220 -123.530 ;
        RECT 44.600 -124.135 44.945 -124.085 ;
        RECT 87.360 -124.260 87.530 -122.245 ;
        RECT 88.415 -124.120 88.585 -122.220 ;
        RECT 88.870 -122.270 89.095 -122.050 ;
        RECT 88.380 -124.440 88.610 -124.120 ;
        RECT 88.905 -124.260 89.075 -122.270 ;
        RECT 89.380 -122.450 89.630 -121.305 ;
        RECT 92.735 -121.460 93.450 -121.375 ;
        RECT 91.320 -121.640 93.450 -121.460 ;
        RECT 92.735 -121.675 93.450 -121.640 ;
        RECT 92.085 -122.050 93.825 -121.870 ;
        RECT 92.085 -122.245 92.265 -122.050 ;
        RECT 89.395 -124.120 89.565 -122.450 ;
        RECT 89.370 -124.440 89.600 -124.120 ;
        RECT 92.090 -124.260 92.260 -122.245 ;
        RECT 93.145 -124.120 93.315 -122.220 ;
        RECT 93.600 -122.270 93.825 -122.050 ;
        RECT 88.380 -124.630 89.600 -124.440 ;
        RECT 93.110 -124.440 93.340 -124.120 ;
        RECT 93.635 -124.260 93.805 -122.270 ;
        RECT 94.110 -122.450 94.360 -121.225 ;
        RECT 94.125 -124.120 94.295 -122.450 ;
        RECT 94.560 -122.550 94.860 -121.720 ;
        RECT 95.735 -122.160 95.905 -121.225 ;
        RECT 96.180 -121.710 96.350 -119.855 ;
        RECT 96.670 -121.395 96.840 -119.245 ;
        RECT 97.730 -119.360 99.935 -119.190 ;
        RECT 97.730 -119.375 98.885 -119.360 ;
        RECT 97.160 -121.705 97.330 -119.855 ;
        RECT 97.730 -119.895 97.905 -119.375 ;
        RECT 97.730 -121.390 97.900 -119.895 ;
        RECT 98.220 -121.390 98.390 -119.850 ;
        RECT 98.710 -119.905 98.885 -119.375 ;
        RECT 98.710 -121.390 98.880 -119.905 ;
        RECT 98.220 -121.705 98.395 -121.390 ;
        RECT 97.160 -121.710 98.395 -121.705 ;
        RECT 99.275 -121.710 99.445 -119.850 ;
        RECT 99.765 -121.390 99.935 -119.360 ;
        RECT 100.255 -121.710 100.425 -119.850 ;
        RECT 101.830 -120.890 102.000 -118.910 ;
        RECT 102.340 -118.990 103.920 -118.910 ;
        RECT 102.340 -119.165 103.915 -118.990 ;
        RECT 96.180 -121.880 98.395 -121.710 ;
        RECT 99.260 -121.880 100.425 -121.710 ;
        RECT 102.320 -121.815 102.490 -119.850 ;
        RECT 103.510 -120.695 103.915 -119.165 ;
        RECT 105.725 -120.680 105.895 -119.120 ;
        RECT 106.215 -120.260 106.385 -119.120 ;
        RECT 106.775 -120.260 106.945 -119.120 ;
        RECT 107.265 -120.160 107.435 -118.740 ;
        RECT 107.915 -118.805 108.215 -118.740 ;
        RECT 106.215 -120.435 106.945 -120.260 ;
        RECT 105.560 -120.695 107.955 -120.680 ;
        RECT 108.405 -120.695 108.755 -115.510 ;
        RECT 103.510 -121.485 108.755 -120.695 ;
        RECT 105.430 -121.700 108.755 -121.485 ;
        RECT 109.040 -119.905 109.390 -116.235 ;
        RECT 109.875 -119.615 110.045 -115.510 ;
        RECT 110.365 -119.895 110.535 -116.075 ;
        RECT 111.875 -119.615 112.045 -115.510 ;
        RECT 111.525 -119.895 112.195 -119.830 ;
        RECT 109.040 -120.175 110.185 -119.905 ;
        RECT 110.365 -120.065 112.195 -119.895 ;
        RECT 98.415 -122.160 99.090 -122.125 ;
        RECT 95.710 -122.330 99.090 -122.160 ;
        RECT 98.415 -122.395 99.090 -122.330 ;
        RECT 99.260 -122.150 99.445 -121.880 ;
        RECT 102.320 -121.995 103.705 -121.815 ;
        RECT 101.470 -122.150 102.145 -122.115 ;
        RECT 99.260 -122.335 102.145 -122.150 ;
        RECT 97.475 -122.550 98.150 -122.515 ;
        RECT 94.560 -122.740 98.150 -122.550 ;
        RECT 97.475 -122.785 98.150 -122.740 ;
        RECT 95.795 -122.970 96.470 -122.925 ;
        RECT 95.135 -123.145 96.470 -122.970 ;
        RECT 99.260 -123.025 99.445 -122.335 ;
        RECT 101.470 -122.385 102.145 -122.335 ;
        RECT 95.135 -123.630 95.435 -123.145 ;
        RECT 95.700 -123.155 96.470 -123.145 ;
        RECT 95.795 -123.195 96.470 -123.155 ;
        RECT 96.670 -123.210 99.445 -123.025 ;
        RECT 94.100 -124.440 94.330 -124.120 ;
        RECT 96.670 -124.430 96.840 -123.210 ;
        RECT 97.650 -124.430 97.820 -123.210 ;
        RECT 98.630 -124.430 98.800 -123.210 ;
        RECT 102.320 -124.430 102.490 -121.995 ;
        RECT 103.050 -122.115 103.705 -121.995 ;
        RECT 105.475 -122.495 105.645 -121.700 ;
        RECT 105.965 -122.415 106.135 -121.955 ;
        RECT 104.915 -123.035 105.755 -122.665 ;
        RECT 105.935 -122.880 106.165 -122.415 ;
        RECT 106.455 -122.495 106.625 -121.700 ;
        RECT 106.945 -122.415 107.115 -121.955 ;
        RECT 106.915 -122.880 107.145 -122.415 ;
        RECT 107.435 -122.495 107.605 -121.700 ;
        RECT 107.925 -122.415 108.095 -121.955 ;
        RECT 107.895 -122.720 108.125 -122.415 ;
        RECT 109.040 -122.720 109.390 -120.175 ;
        RECT 107.895 -122.880 109.390 -122.720 ;
        RECT 105.935 -123.070 109.390 -122.880 ;
        RECT 105.935 -123.110 108.125 -123.070 ;
        RECT 105.935 -124.375 106.165 -123.110 ;
        RECT 106.915 -123.435 107.145 -123.110 ;
        RECT 107.895 -123.435 108.125 -123.110 ;
        RECT 105.965 -124.395 106.135 -124.375 ;
        RECT 106.945 -124.395 107.115 -123.435 ;
        RECT 107.925 -124.395 108.095 -123.435 ;
        RECT 110.365 -124.040 110.535 -120.065 ;
        RECT 111.525 -120.100 112.195 -120.065 ;
        RECT 112.365 -119.845 112.535 -116.075 ;
        RECT 112.905 -119.845 113.495 -119.785 ;
        RECT 112.365 -120.015 113.495 -119.845 ;
        RECT 112.365 -124.040 112.535 -120.015 ;
        RECT 112.905 -120.075 113.495 -120.015 ;
        RECT 114.260 -119.895 114.610 -118.990 ;
        RECT 114.875 -119.615 115.045 -115.510 ;
        RECT 114.260 -120.165 115.130 -119.895 ;
        RECT 115.365 -119.945 115.535 -116.075 ;
        RECT 116.875 -119.615 117.045 -115.510 ;
        RECT 116.525 -119.945 117.195 -119.905 ;
        RECT 115.365 -120.140 117.195 -119.945 ;
        RECT 115.365 -124.040 115.535 -120.140 ;
        RECT 116.525 -120.175 117.195 -120.140 ;
        RECT 117.365 -119.980 117.535 -116.075 ;
        RECT 118.290 -119.980 118.880 -119.920 ;
        RECT 117.365 -120.150 118.880 -119.980 ;
        RECT 117.365 -124.040 117.535 -120.150 ;
        RECT 118.290 -120.210 118.880 -120.150 ;
        RECT 119.215 -119.930 119.565 -118.995 ;
        RECT 119.875 -119.615 120.045 -115.510 ;
        RECT 119.215 -120.200 120.130 -119.930 ;
        RECT 120.365 -119.950 120.535 -116.075 ;
        RECT 121.875 -119.615 122.045 -115.510 ;
        RECT 122.365 -119.900 122.535 -116.075 ;
        RECT 133.425 -116.205 133.805 -110.845 ;
        RECT 134.500 -110.850 136.930 -110.845 ;
        RECT 134.500 -110.855 134.855 -110.850 ;
        RECT 136.560 -110.880 136.930 -110.850 ;
        RECT 134.660 -112.605 134.830 -111.065 ;
        RECT 135.150 -112.605 135.320 -111.065 ;
        RECT 135.640 -112.605 135.810 -111.065 ;
        RECT 136.130 -112.605 136.300 -111.065 ;
        RECT 136.620 -112.605 136.790 -111.065 ;
        RECT 135.145 -112.865 135.320 -112.605 ;
        RECT 138.715 -112.775 139.020 -110.740 ;
        RECT 141.165 -111.560 141.515 -109.585 ;
        RECT 142.385 -110.855 142.555 -107.935 ;
        RECT 143.420 -107.975 143.630 -107.765 ;
        RECT 142.365 -111.150 142.575 -110.855 ;
        RECT 143.440 -110.885 143.610 -107.975 ;
        RECT 143.930 -110.875 144.100 -107.935 ;
        RECT 144.410 -107.985 144.620 -107.765 ;
        RECT 143.425 -111.150 143.635 -110.885 ;
        RECT 142.365 -111.330 143.635 -111.150 ;
        RECT 143.910 -111.145 144.120 -110.875 ;
        RECT 144.420 -110.975 144.590 -107.985 ;
        RECT 145.480 -110.905 145.650 -107.935 ;
        RECT 143.910 -111.340 144.615 -111.145 ;
        RECT 144.400 -111.400 144.615 -111.340 ;
        RECT 143.190 -111.560 143.965 -111.510 ;
        RECT 141.165 -111.740 143.965 -111.560 ;
        RECT 141.165 -111.750 141.515 -111.740 ;
        RECT 143.190 -111.785 143.965 -111.740 ;
        RECT 144.400 -111.675 145.305 -111.400 ;
        RECT 144.400 -112.025 144.615 -111.675 ;
        RECT 141.840 -112.095 142.615 -112.050 ;
        RECT 141.655 -112.265 142.615 -112.095 ;
        RECT 141.840 -112.325 142.615 -112.265 ;
        RECT 142.845 -112.225 144.615 -112.025 ;
        RECT 145.475 -112.125 145.690 -110.905 ;
        RECT 146.660 -111.250 147.010 -104.565 ;
        RECT 177.480 -104.830 177.650 -103.790 ;
        RECT 178.460 -104.830 178.630 -103.790 ;
        RECT 179.440 -104.830 179.610 -103.790 ;
        RECT 182.345 -105.475 182.515 -103.755 ;
        RECT 183.325 -105.475 183.495 -103.755 ;
        RECT 184.190 -104.500 184.495 -103.755 ;
        RECT 185.390 -104.325 185.560 -103.545 ;
        RECT 185.880 -104.325 186.050 -103.785 ;
        RECT 186.370 -104.325 186.540 -103.545 ;
        RECT 220.335 -103.750 221.570 -103.545 ;
        RECT 225.745 -103.685 226.420 -103.645 ;
        RECT 225.645 -103.695 226.420 -103.685 ;
        RECT 186.860 -104.325 187.030 -103.785 ;
        RECT 220.335 -103.835 220.985 -103.750 ;
        RECT 221.205 -103.815 221.570 -103.750 ;
        RECT 224.610 -103.875 226.420 -103.695 ;
        RECT 229.005 -103.740 232.930 -103.310 ;
        RECT 266.325 -103.375 266.975 -102.915 ;
        RECT 267.785 -103.205 267.955 -101.925 ;
        RECT 268.275 -103.205 268.445 -102.165 ;
        RECT 268.765 -103.205 268.935 -101.925 ;
        RECT 269.255 -103.035 269.425 -102.165 ;
        RECT 272.160 -102.815 272.330 -101.275 ;
        RECT 272.650 -102.815 272.820 -101.275 ;
        RECT 273.140 -102.815 273.310 -101.275 ;
        RECT 273.630 -102.815 273.800 -101.275 ;
        RECT 274.120 -102.815 274.290 -101.275 ;
        RECT 272.000 -103.030 272.355 -103.025 ;
        RECT 274.060 -103.030 274.430 -103.000 ;
        RECT 272.000 -103.035 274.430 -103.030 ;
        RECT 269.255 -103.205 274.430 -103.035 ;
        RECT 276.215 -103.140 276.520 -101.105 ;
        RECT 299.455 -101.255 308.710 -100.500 ;
        RECT 315.115 -100.470 318.440 -100.330 ;
        RECT 315.115 -100.760 320.290 -100.470 ;
        RECT 315.115 -101.165 315.545 -100.760 ;
        RECT 316.415 -100.945 316.590 -100.760 ;
        RECT 318.040 -100.775 320.290 -100.760 ;
        RECT 299.455 -101.595 301.335 -101.255 ;
        RECT 307.460 -101.510 308.710 -101.255 ;
        RECT 310.855 -101.595 315.545 -101.165 ;
        RECT 310.095 -103.045 310.745 -102.585 ;
        RECT 311.555 -102.875 311.725 -101.595 ;
        RECT 312.045 -102.875 312.215 -101.835 ;
        RECT 312.535 -102.875 312.705 -101.595 ;
        RECT 313.025 -102.705 313.195 -101.835 ;
        RECT 315.930 -102.485 316.100 -100.945 ;
        RECT 316.420 -102.485 316.590 -100.945 ;
        RECT 316.910 -102.485 317.080 -100.945 ;
        RECT 317.400 -102.485 317.570 -100.945 ;
        RECT 317.890 -102.485 318.060 -100.945 ;
        RECT 315.770 -102.700 316.125 -102.695 ;
        RECT 317.830 -102.700 318.200 -102.670 ;
        RECT 315.770 -102.705 318.200 -102.700 ;
        RECT 313.025 -102.875 318.200 -102.705 ;
        RECT 319.985 -102.810 320.290 -100.775 ;
        RECT 343.335 -100.530 345.025 -100.050 ;
        RECT 362.215 -100.245 363.915 -98.275 ;
        RECT 389.485 -100.225 390.835 -99.620 ;
        RECT 399.550 -100.225 401.025 -100.015 ;
        RECT 408.895 -100.055 409.950 -98.275 ;
        RECT 353.275 -100.530 354.615 -100.325 ;
        RECT 343.335 -101.185 354.615 -100.530 ;
        RECT 360.880 -100.385 364.205 -100.245 ;
        RECT 360.880 -100.675 366.055 -100.385 ;
        RECT 360.880 -101.080 361.310 -100.675 ;
        RECT 362.180 -100.860 362.355 -100.675 ;
        RECT 363.805 -100.690 366.055 -100.675 ;
        RECT 343.335 -101.505 345.025 -101.185 ;
        RECT 353.275 -101.525 354.615 -101.185 ;
        RECT 356.620 -101.510 361.310 -101.080 ;
        RECT 313.030 -102.895 318.200 -102.875 ;
        RECT 313.030 -102.905 315.775 -102.895 ;
        RECT 310.965 -103.045 311.330 -103.015 ;
        RECT 317.830 -103.025 318.200 -102.895 ;
        RECT 269.260 -103.225 274.430 -103.205 ;
        RECT 269.260 -103.235 272.005 -103.225 ;
        RECT 267.195 -103.375 267.560 -103.345 ;
        RECT 274.060 -103.355 274.430 -103.225 ;
        RECT 266.325 -103.580 267.560 -103.375 ;
        RECT 271.735 -103.515 272.410 -103.475 ;
        RECT 271.635 -103.525 272.410 -103.515 ;
        RECT 266.325 -103.665 266.975 -103.580 ;
        RECT 267.195 -103.645 267.560 -103.580 ;
        RECT 270.600 -103.705 272.410 -103.525 ;
        RECT 274.995 -103.570 278.920 -103.140 ;
        RECT 310.095 -103.250 311.330 -103.045 ;
        RECT 315.505 -103.185 316.180 -103.145 ;
        RECT 315.405 -103.195 316.180 -103.185 ;
        RECT 310.095 -103.335 310.745 -103.250 ;
        RECT 310.965 -103.315 311.330 -103.250 ;
        RECT 314.370 -103.375 316.180 -103.195 ;
        RECT 318.765 -103.240 322.690 -102.810 ;
        RECT 355.860 -102.960 356.510 -102.500 ;
        RECT 357.320 -102.790 357.490 -101.510 ;
        RECT 357.810 -102.790 357.980 -101.750 ;
        RECT 358.300 -102.790 358.470 -101.510 ;
        RECT 358.790 -102.620 358.960 -101.750 ;
        RECT 361.695 -102.400 361.865 -100.860 ;
        RECT 362.185 -102.400 362.355 -100.860 ;
        RECT 362.675 -102.400 362.845 -100.860 ;
        RECT 363.165 -102.400 363.335 -100.860 ;
        RECT 363.655 -102.400 363.825 -100.860 ;
        RECT 361.535 -102.615 361.890 -102.610 ;
        RECT 363.595 -102.615 363.965 -102.585 ;
        RECT 361.535 -102.620 363.965 -102.615 ;
        RECT 358.790 -102.790 363.965 -102.620 ;
        RECT 365.750 -102.725 366.055 -100.690 ;
        RECT 389.485 -100.920 401.025 -100.225 ;
        RECT 407.700 -100.195 411.025 -100.055 ;
        RECT 407.700 -100.485 412.875 -100.195 ;
        RECT 407.700 -100.890 408.130 -100.485 ;
        RECT 409.000 -100.670 409.175 -100.485 ;
        RECT 410.625 -100.500 412.875 -100.485 ;
        RECT 389.485 -101.045 390.835 -100.920 ;
        RECT 399.550 -101.380 401.025 -100.920 ;
        RECT 403.440 -101.320 408.130 -100.890 ;
        RECT 358.795 -102.810 363.965 -102.790 ;
        RECT 358.795 -102.820 361.540 -102.810 ;
        RECT 356.730 -102.960 357.095 -102.930 ;
        RECT 363.595 -102.940 363.965 -102.810 ;
        RECT 355.860 -103.165 357.095 -102.960 ;
        RECT 361.270 -103.100 361.945 -103.060 ;
        RECT 361.170 -103.110 361.945 -103.100 ;
        RECT 315.405 -103.385 316.180 -103.375 ;
        RECT 315.505 -103.415 316.180 -103.385 ;
        RECT 316.420 -103.300 318.515 -103.260 ;
        RECT 316.420 -103.450 318.570 -103.300 ;
        RECT 271.635 -103.715 272.410 -103.705 ;
        RECT 225.645 -103.885 226.420 -103.875 ;
        RECT 225.745 -103.915 226.420 -103.885 ;
        RECT 226.660 -103.800 228.755 -103.760 ;
        RECT 226.660 -103.950 228.810 -103.800 ;
        RECT 184.800 -104.500 185.165 -104.470 ;
        RECT 184.190 -104.565 185.165 -104.500 ;
        RECT 184.300 -104.705 185.165 -104.565 ;
        RECT 184.800 -104.770 185.165 -104.705 ;
        RECT 187.350 -104.620 189.210 -104.270 ;
        RECT 185.390 -105.480 185.560 -104.940 ;
        RECT 186.370 -105.480 186.540 -104.940 ;
        RECT 187.350 -105.480 187.520 -104.620 ;
        RECT 153.240 -107.045 154.845 -106.875 ;
        RECT 152.345 -109.725 152.515 -107.225 ;
        RECT 152.340 -109.955 152.515 -109.725 ;
        RECT 153.240 -109.955 153.440 -107.045 ;
        RECT 153.685 -107.245 153.860 -107.045 ;
        RECT 153.690 -109.765 153.860 -107.245 ;
        RECT 154.180 -109.730 154.350 -107.225 ;
        RECT 154.670 -107.240 154.845 -107.045 ;
        RECT 152.340 -110.155 153.440 -109.955 ;
        RECT 154.165 -110.330 154.355 -109.730 ;
        RECT 154.670 -109.765 154.840 -107.240 ;
        RECT 155.320 -110.145 155.490 -107.225 ;
        RECT 156.950 -109.795 157.120 -107.225 ;
        RECT 158.090 -108.675 158.260 -107.225 ;
        RECT 185.620 -107.820 186.820 -107.650 ;
        RECT 158.085 -109.140 158.270 -108.675 ;
        RECT 158.085 -109.325 158.770 -109.140 ;
        RECT 156.950 -109.965 157.745 -109.795 ;
        RECT 156.065 -110.145 156.755 -110.090 ;
        RECT 152.345 -110.520 154.355 -110.330 ;
        RECT 154.690 -110.315 156.755 -110.145 ;
        RECT 151.160 -110.575 151.850 -110.525 ;
        RECT 149.210 -110.745 151.850 -110.575 ;
        RECT 146.605 -111.610 147.130 -111.250 ;
        RECT 149.210 -112.125 149.425 -110.745 ;
        RECT 151.160 -110.795 151.850 -110.745 ;
        RECT 151.440 -111.250 152.130 -111.205 ;
        RECT 150.390 -111.420 152.130 -111.250 ;
        RECT 150.390 -112.055 150.750 -111.420 ;
        RECT 151.440 -111.475 152.130 -111.420 ;
        RECT 150.390 -112.100 150.810 -112.055 ;
        RECT 136.770 -112.865 139.020 -112.775 ;
        RECT 134.560 -113.080 139.020 -112.865 ;
        RECT 134.560 -113.170 136.805 -113.080 ;
        RECT 138.715 -114.555 139.020 -113.080 ;
        RECT 142.385 -113.965 142.555 -112.495 ;
        RECT 142.845 -112.575 143.070 -112.225 ;
        RECT 144.805 -112.325 149.425 -112.125 ;
        RECT 145.045 -112.340 149.425 -112.325 ;
        RECT 142.350 -114.555 142.585 -113.965 ;
        RECT 142.875 -114.035 143.045 -112.575 ;
        RECT 143.365 -113.960 143.535 -112.495 ;
        RECT 144.575 -113.910 144.745 -112.495 ;
        RECT 145.045 -112.540 145.265 -112.340 ;
        RECT 150.415 -112.450 150.810 -112.100 ;
        RECT 143.330 -114.555 143.565 -113.960 ;
        RECT 144.540 -114.555 144.775 -113.910 ;
        RECT 145.065 -114.035 145.235 -112.540 ;
        RECT 151.855 -113.660 152.025 -112.205 ;
        RECT 151.845 -114.215 152.030 -113.660 ;
        RECT 152.345 -113.745 152.515 -110.520 ;
        RECT 153.490 -110.870 153.680 -110.520 ;
        RECT 154.690 -110.710 154.860 -110.315 ;
        RECT 156.065 -110.360 156.755 -110.315 ;
        RECT 153.440 -111.560 153.710 -110.870 ;
        RECT 154.205 -110.880 154.860 -110.710 ;
        RECT 155.190 -110.795 155.880 -110.525 ;
        RECT 157.115 -110.870 157.385 -110.180 ;
        RECT 157.575 -110.185 157.745 -109.965 ;
        RECT 157.575 -110.455 158.405 -110.185 ;
        RECT 154.205 -113.745 154.375 -110.880 ;
        RECT 157.575 -111.030 157.745 -110.455 ;
        RECT 158.005 -111.030 158.275 -110.945 ;
        RECT 154.695 -111.225 155.490 -111.050 ;
        RECT 157.575 -111.055 158.275 -111.030 ;
        RECT 157.435 -111.200 158.275 -111.055 ;
        RECT 154.695 -113.745 154.865 -111.225 ;
        RECT 155.320 -113.745 155.490 -111.225 ;
        RECT 155.810 -113.660 155.980 -111.205 ;
        RECT 156.460 -113.655 156.630 -111.205 ;
        RECT 149.160 -114.235 152.215 -114.215 ;
        RECT 155.805 -114.235 155.990 -113.660 ;
        RECT 156.445 -114.235 156.630 -113.655 ;
        RECT 156.950 -113.745 157.120 -111.205 ;
        RECT 157.435 -111.225 157.745 -111.200 ;
        RECT 157.440 -113.745 157.610 -111.225 ;
        RECT 158.005 -111.240 158.275 -111.200 ;
        RECT 158.580 -111.790 158.770 -109.325 ;
        RECT 170.995 -110.230 174.235 -109.960 ;
        RECT 177.350 -110.155 177.520 -108.435 ;
        RECT 178.330 -110.155 178.500 -108.435 ;
        RECT 180.395 -108.970 180.565 -108.430 ;
        RECT 181.375 -108.970 181.545 -108.430 ;
        RECT 179.805 -109.205 180.170 -109.140 ;
        RECT 179.305 -109.345 180.170 -109.205 ;
        RECT 179.195 -109.410 180.170 -109.345 ;
        RECT 179.195 -110.155 179.500 -109.410 ;
        RECT 179.805 -109.440 180.170 -109.410 ;
        RECT 182.355 -109.290 182.525 -108.430 ;
        RECT 176.435 -110.220 177.110 -110.190 ;
        RECT 176.335 -110.230 177.110 -110.220 ;
        RECT 170.995 -110.410 177.110 -110.230 ;
        RECT 177.350 -110.305 179.500 -110.155 ;
        RECT 177.350 -110.345 179.445 -110.305 ;
        RECT 180.395 -110.365 180.565 -109.585 ;
        RECT 180.885 -110.125 181.055 -109.585 ;
        RECT 181.375 -110.365 181.545 -109.585 ;
        RECT 181.865 -110.125 182.035 -109.585 ;
        RECT 182.355 -109.640 183.745 -109.290 ;
        RECT 170.995 -110.690 174.235 -110.410 ;
        RECT 176.335 -110.420 177.110 -110.410 ;
        RECT 176.435 -110.460 177.110 -110.420 ;
        RECT 158.580 -111.980 160.040 -111.790 ;
        RECT 158.090 -113.650 158.260 -112.205 ;
        RECT 158.580 -112.230 158.770 -111.980 ;
        RECT 158.080 -114.235 158.265 -113.650 ;
        RECT 158.580 -113.745 158.750 -112.230 ;
        RECT 149.160 -114.555 158.830 -114.235 ;
        RECT 138.715 -114.780 158.830 -114.555 ;
        RECT 138.715 -115.120 149.725 -114.780 ;
        RECT 151.465 -115.040 158.830 -114.780 ;
        RECT 129.445 -116.485 133.805 -116.205 ;
        RECT 159.850 -116.455 160.040 -111.980 ;
        RECT 129.445 -116.865 149.975 -116.485 ;
        RECT 129.445 -116.935 133.805 -116.865 ;
        RECT 122.770 -119.900 123.360 -119.860 ;
        RECT 121.490 -119.950 122.160 -119.915 ;
        RECT 120.365 -120.145 122.160 -119.950 ;
        RECT 120.365 -124.040 120.535 -120.145 ;
        RECT 121.490 -120.185 122.160 -120.145 ;
        RECT 122.365 -120.070 123.375 -119.900 ;
        RECT 122.365 -124.040 122.535 -120.070 ;
        RECT 122.770 -120.150 123.360 -120.070 ;
        RECT 93.110 -124.630 94.330 -124.440 ;
        RECT 42.185 -127.025 47.035 -125.720 ;
        RECT 42.145 -127.590 43.100 -127.560 ;
        RECT 42.145 -128.005 44.960 -127.590 ;
        RECT 42.145 -128.095 43.100 -128.005 ;
        RECT -31.240 -131.835 -28.080 -131.790 ;
        RECT -18.740 -131.835 -15.580 -131.790 ;
        RECT -6.240 -131.835 -3.080 -131.790 ;
        RECT 6.260 -131.835 9.420 -131.790 ;
        RECT 18.760 -131.835 21.920 -131.790 ;
        RECT 33.680 -131.835 39.020 -131.725 ;
        RECT -37.245 -131.840 -28.080 -131.835 ;
        RECT -24.745 -131.840 39.020 -131.835 ;
        RECT -37.245 -132.100 39.020 -131.840 ;
        RECT -37.245 -132.715 -37.050 -132.100 ;
        RECT -31.240 -132.270 -24.550 -132.100 ;
        RECT -18.740 -132.270 -15.580 -132.100 ;
        RECT -36.735 -132.470 -31.695 -132.290 ;
        RECT -37.225 -133.660 -37.055 -132.715 ;
        RECT -37.235 -134.075 -37.050 -133.660 ;
        RECT -36.735 -133.695 -36.565 -132.470 ;
        RECT -35.155 -133.665 -34.985 -132.655 ;
        RECT -34.665 -133.650 -34.495 -132.655 ;
        RECT -33.345 -133.650 -33.175 -132.655 ;
        RECT -35.170 -133.770 -34.985 -133.665 ;
        RECT -35.765 -133.955 -34.985 -133.770 ;
        RECT -34.675 -133.845 -33.175 -133.650 ;
        RECT -35.765 -134.075 -35.580 -133.955 ;
        RECT -37.235 -134.260 -35.580 -134.075 ;
        RECT -32.855 -134.110 -32.685 -132.655 ;
        RECT -31.875 -132.740 -31.695 -132.470 ;
        RECT -31.875 -133.695 -31.705 -132.740 ;
        RECT -31.385 -134.110 -31.215 -132.655 ;
        RECT -30.325 -133.610 -30.155 -132.655 ;
        RECT -29.860 -132.690 -29.645 -132.270 ;
        RECT -28.685 -132.275 -24.550 -132.270 ;
        RECT -30.350 -133.835 -30.135 -133.610 ;
        RECT -29.835 -133.695 -29.665 -132.690 ;
        RECT -28.780 -133.600 -28.610 -132.655 ;
        RECT -28.315 -132.700 -28.100 -132.275 ;
        RECT -30.830 -134.065 -30.135 -133.835 ;
        RECT -34.020 -134.280 -31.215 -134.110 ;
        RECT -34.020 -134.590 -33.850 -134.280 ;
        RECT -37.230 -134.935 -36.535 -134.665 ;
        RECT -34.580 -134.760 -33.850 -134.590 ;
        RECT -34.580 -135.335 -34.410 -134.760 ;
        RECT -33.485 -134.785 -32.790 -134.515 ;
        RECT -37.780 -135.505 -34.410 -135.335 ;
        RECT -34.105 -135.140 -31.705 -134.970 ;
        RECT -91.335 -135.660 -88.010 -135.520 ;
        RECT -111.230 -135.935 -108.455 -135.750 ;
        RECT -108.255 -135.870 -99.165 -135.695 ;
        RECT -108.255 -135.880 -107.485 -135.870 ;
        RECT -108.255 -135.920 -107.580 -135.880 ;
        RECT -99.455 -135.895 -99.165 -135.870 ;
        RECT -110.585 -137.155 -110.415 -135.935 ;
        RECT -109.605 -137.155 -109.435 -135.935 ;
        RECT -108.625 -137.155 -108.455 -135.935 ;
        RECT -45.730 -136.475 -44.730 -136.355 ;
        RECT -97.635 -137.155 -44.730 -136.475 ;
        RECT -45.730 -137.210 -44.730 -137.155 ;
        RECT -37.225 -137.245 -37.055 -135.685 ;
        RECT -36.735 -136.725 -36.565 -135.505 ;
        RECT -36.245 -137.245 -36.075 -135.685 ;
        RECT -35.645 -136.900 -35.475 -135.685 ;
        RECT -35.155 -136.725 -34.985 -135.505 ;
        RECT -34.665 -136.900 -34.495 -135.685 ;
        RECT -34.105 -136.900 -33.935 -135.140 ;
        RECT -35.645 -137.070 -33.935 -136.900 ;
        RECT -33.755 -135.510 -32.685 -135.340 ;
        RECT -33.755 -137.245 -33.585 -135.510 ;
        RECT -32.855 -136.725 -32.685 -135.510 ;
        RECT -31.875 -136.725 -31.705 -135.140 ;
        RECT -31.440 -135.155 -30.745 -134.885 ;
        RECT -30.350 -135.760 -30.135 -134.065 ;
        RECT -28.800 -134.555 -28.585 -133.600 ;
        RECT -28.290 -133.695 -28.120 -132.700 ;
        RECT -24.745 -132.715 -24.550 -132.275 ;
        RECT -24.235 -132.470 -19.195 -132.290 ;
        RECT -25.595 -133.520 -25.365 -132.840 ;
        RECT -29.300 -134.785 -28.585 -134.555 ;
        RECT -30.325 -136.725 -30.155 -135.760 ;
        RECT -28.800 -135.770 -28.585 -134.785 ;
        RECT -28.365 -135.125 -27.670 -134.855 ;
        RECT -25.565 -135.335 -25.395 -133.520 ;
        RECT -24.725 -133.660 -24.555 -132.715 ;
        RECT -24.735 -134.075 -24.550 -133.660 ;
        RECT -24.235 -133.695 -24.065 -132.470 ;
        RECT -22.655 -133.665 -22.485 -132.655 ;
        RECT -22.165 -133.650 -21.995 -132.655 ;
        RECT -20.845 -133.650 -20.675 -132.655 ;
        RECT -22.670 -133.770 -22.485 -133.665 ;
        RECT -23.265 -133.955 -22.485 -133.770 ;
        RECT -22.175 -133.845 -20.675 -133.650 ;
        RECT -23.265 -134.075 -23.080 -133.955 ;
        RECT -24.735 -134.260 -23.080 -134.075 ;
        RECT -20.355 -134.110 -20.185 -132.655 ;
        RECT -19.375 -132.740 -19.195 -132.470 ;
        RECT -19.375 -133.695 -19.205 -132.740 ;
        RECT -18.885 -134.110 -18.715 -132.655 ;
        RECT -17.825 -133.610 -17.655 -132.655 ;
        RECT -17.360 -132.690 -17.145 -132.270 ;
        RECT -17.850 -133.835 -17.635 -133.610 ;
        RECT -17.335 -133.695 -17.165 -132.690 ;
        RECT -16.280 -133.600 -16.110 -132.655 ;
        RECT -15.815 -132.700 -15.600 -132.270 ;
        RECT -18.330 -134.065 -17.635 -133.835 ;
        RECT -21.520 -134.280 -18.715 -134.110 ;
        RECT -21.520 -134.590 -21.350 -134.280 ;
        RECT -24.730 -134.935 -24.035 -134.665 ;
        RECT -22.080 -134.760 -21.350 -134.590 ;
        RECT -22.080 -135.335 -21.910 -134.760 ;
        RECT -20.985 -134.785 -20.290 -134.515 ;
        RECT -25.565 -135.505 -21.910 -135.335 ;
        RECT -21.605 -135.140 -19.205 -134.970 ;
        RECT -28.780 -136.725 -28.610 -135.770 ;
        RECT -37.225 -137.415 -33.585 -137.245 ;
        RECT -24.725 -137.245 -24.555 -135.685 ;
        RECT -24.235 -136.725 -24.065 -135.505 ;
        RECT -23.745 -137.245 -23.575 -135.685 ;
        RECT -23.145 -136.900 -22.975 -135.685 ;
        RECT -22.655 -136.725 -22.485 -135.505 ;
        RECT -22.165 -136.900 -21.995 -135.685 ;
        RECT -21.605 -136.900 -21.435 -135.140 ;
        RECT -23.145 -137.070 -21.435 -136.900 ;
        RECT -21.255 -135.510 -20.185 -135.340 ;
        RECT -21.255 -137.245 -21.085 -135.510 ;
        RECT -20.355 -136.725 -20.185 -135.510 ;
        RECT -19.375 -136.725 -19.205 -135.140 ;
        RECT -18.940 -135.155 -18.245 -134.885 ;
        RECT -17.850 -135.760 -17.635 -134.065 ;
        RECT -16.300 -134.555 -16.085 -133.600 ;
        RECT -15.790 -133.695 -15.620 -132.700 ;
        RECT -12.245 -132.715 -12.050 -132.100 ;
        RECT -6.240 -132.270 -3.080 -132.100 ;
        RECT -11.735 -132.470 -6.695 -132.290 ;
        RECT -12.855 -133.500 -12.625 -132.820 ;
        RECT -16.800 -134.785 -16.085 -134.555 ;
        RECT -17.825 -136.725 -17.655 -135.760 ;
        RECT -16.300 -135.770 -16.085 -134.785 ;
        RECT -15.865 -135.125 -15.170 -134.855 ;
        RECT -12.825 -135.335 -12.655 -133.500 ;
        RECT -12.225 -133.660 -12.055 -132.715 ;
        RECT -12.235 -134.075 -12.050 -133.660 ;
        RECT -11.735 -133.695 -11.565 -132.470 ;
        RECT -10.155 -133.665 -9.985 -132.655 ;
        RECT -9.665 -133.650 -9.495 -132.655 ;
        RECT -8.345 -133.650 -8.175 -132.655 ;
        RECT -10.170 -133.770 -9.985 -133.665 ;
        RECT -10.765 -133.955 -9.985 -133.770 ;
        RECT -9.675 -133.845 -8.175 -133.650 ;
        RECT -10.765 -134.075 -10.580 -133.955 ;
        RECT -12.235 -134.260 -10.580 -134.075 ;
        RECT -7.855 -134.110 -7.685 -132.655 ;
        RECT -6.875 -132.740 -6.695 -132.470 ;
        RECT -6.875 -133.695 -6.705 -132.740 ;
        RECT -6.385 -134.110 -6.215 -132.655 ;
        RECT -5.325 -133.610 -5.155 -132.655 ;
        RECT -4.860 -132.690 -4.645 -132.270 ;
        RECT -5.350 -133.835 -5.135 -133.610 ;
        RECT -4.835 -133.695 -4.665 -132.690 ;
        RECT -3.780 -133.600 -3.610 -132.655 ;
        RECT -3.315 -132.700 -3.100 -132.270 ;
        RECT -5.830 -134.065 -5.135 -133.835 ;
        RECT -9.020 -134.280 -6.215 -134.110 ;
        RECT -9.020 -134.590 -8.850 -134.280 ;
        RECT -12.230 -134.935 -11.535 -134.665 ;
        RECT -9.580 -134.760 -8.850 -134.590 ;
        RECT -9.580 -135.335 -9.410 -134.760 ;
        RECT -8.485 -134.785 -7.790 -134.515 ;
        RECT -12.825 -135.505 -9.410 -135.335 ;
        RECT -9.105 -135.140 -6.705 -134.970 ;
        RECT -16.280 -136.725 -16.110 -135.770 ;
        RECT -24.725 -137.415 -21.085 -137.245 ;
        RECT -12.225 -137.245 -12.055 -135.685 ;
        RECT -11.735 -136.725 -11.565 -135.505 ;
        RECT -11.245 -137.245 -11.075 -135.685 ;
        RECT -10.645 -136.900 -10.475 -135.685 ;
        RECT -10.155 -136.725 -9.985 -135.505 ;
        RECT -9.665 -136.900 -9.495 -135.685 ;
        RECT -9.105 -136.900 -8.935 -135.140 ;
        RECT -10.645 -137.070 -8.935 -136.900 ;
        RECT -8.755 -135.510 -7.685 -135.340 ;
        RECT -8.755 -137.245 -8.585 -135.510 ;
        RECT -7.855 -136.725 -7.685 -135.510 ;
        RECT -6.875 -136.725 -6.705 -135.140 ;
        RECT -6.440 -135.155 -5.745 -134.885 ;
        RECT -5.350 -135.760 -5.135 -134.065 ;
        RECT -3.800 -134.555 -3.585 -133.600 ;
        RECT -3.290 -133.695 -3.120 -132.700 ;
        RECT 0.255 -132.715 0.450 -132.100 ;
        RECT 6.260 -132.270 9.420 -132.100 ;
        RECT 0.765 -132.470 5.805 -132.290 ;
        RECT -0.455 -133.500 -0.225 -132.820 ;
        RECT -4.300 -134.785 -3.585 -134.555 ;
        RECT -5.325 -136.725 -5.155 -135.760 ;
        RECT -3.800 -135.770 -3.585 -134.785 ;
        RECT -3.365 -135.125 -2.670 -134.855 ;
        RECT -0.425 -135.335 -0.255 -133.500 ;
        RECT 0.275 -133.660 0.445 -132.715 ;
        RECT 0.265 -134.075 0.450 -133.660 ;
        RECT 0.765 -133.695 0.935 -132.470 ;
        RECT 2.345 -133.665 2.515 -132.655 ;
        RECT 2.835 -133.650 3.005 -132.655 ;
        RECT 4.155 -133.650 4.325 -132.655 ;
        RECT 2.330 -133.770 2.515 -133.665 ;
        RECT 1.735 -133.955 2.515 -133.770 ;
        RECT 2.825 -133.845 4.325 -133.650 ;
        RECT 1.735 -134.075 1.920 -133.955 ;
        RECT 0.265 -134.260 1.920 -134.075 ;
        RECT 4.645 -134.110 4.815 -132.655 ;
        RECT 5.625 -132.740 5.805 -132.470 ;
        RECT 5.625 -133.695 5.795 -132.740 ;
        RECT 6.115 -134.110 6.285 -132.655 ;
        RECT 7.175 -133.610 7.345 -132.655 ;
        RECT 7.640 -132.690 7.855 -132.270 ;
        RECT 7.150 -133.835 7.365 -133.610 ;
        RECT 7.665 -133.695 7.835 -132.690 ;
        RECT 8.720 -133.600 8.890 -132.655 ;
        RECT 9.185 -132.700 9.400 -132.270 ;
        RECT 6.670 -134.065 7.365 -133.835 ;
        RECT 3.480 -134.280 6.285 -134.110 ;
        RECT 3.480 -134.590 3.650 -134.280 ;
        RECT 0.270 -134.935 0.965 -134.665 ;
        RECT 2.920 -134.760 3.650 -134.590 ;
        RECT 2.920 -135.335 3.090 -134.760 ;
        RECT 4.015 -134.785 4.710 -134.515 ;
        RECT -0.425 -135.505 3.090 -135.335 ;
        RECT 3.395 -135.140 5.795 -134.970 ;
        RECT -0.425 -135.510 -0.255 -135.505 ;
        RECT -3.780 -136.725 -3.610 -135.770 ;
        RECT -12.225 -137.415 -8.585 -137.245 ;
        RECT 0.275 -137.245 0.445 -135.685 ;
        RECT 0.765 -136.725 0.935 -135.505 ;
        RECT 1.255 -137.245 1.425 -135.685 ;
        RECT 1.855 -136.900 2.025 -135.685 ;
        RECT 2.345 -136.725 2.515 -135.505 ;
        RECT 2.835 -136.900 3.005 -135.685 ;
        RECT 3.395 -136.900 3.565 -135.140 ;
        RECT 1.855 -137.070 3.565 -136.900 ;
        RECT 3.745 -135.510 4.815 -135.340 ;
        RECT 3.745 -137.245 3.915 -135.510 ;
        RECT 4.645 -136.725 4.815 -135.510 ;
        RECT 5.625 -136.725 5.795 -135.140 ;
        RECT 6.060 -135.155 6.755 -134.885 ;
        RECT 7.150 -135.760 7.365 -134.065 ;
        RECT 8.700 -134.555 8.915 -133.600 ;
        RECT 9.210 -133.695 9.380 -132.700 ;
        RECT 12.755 -132.715 12.950 -132.100 ;
        RECT 18.760 -132.270 21.920 -132.100 ;
        RECT 13.265 -132.470 18.305 -132.290 ;
        RECT 11.630 -133.500 11.860 -132.820 ;
        RECT 11.655 -133.505 11.830 -133.500 ;
        RECT 8.200 -134.785 8.915 -134.555 ;
        RECT 7.175 -136.725 7.345 -135.760 ;
        RECT 8.700 -135.770 8.915 -134.785 ;
        RECT 9.135 -135.125 9.830 -134.855 ;
        RECT 11.655 -135.335 11.825 -133.505 ;
        RECT 12.775 -133.660 12.945 -132.715 ;
        RECT 12.765 -134.075 12.950 -133.660 ;
        RECT 13.265 -133.695 13.435 -132.470 ;
        RECT 14.845 -133.665 15.015 -132.655 ;
        RECT 15.335 -133.650 15.505 -132.655 ;
        RECT 16.655 -133.650 16.825 -132.655 ;
        RECT 14.830 -133.770 15.015 -133.665 ;
        RECT 14.235 -133.955 15.015 -133.770 ;
        RECT 15.325 -133.845 16.825 -133.650 ;
        RECT 14.235 -134.075 14.420 -133.955 ;
        RECT 12.765 -134.260 14.420 -134.075 ;
        RECT 17.145 -134.110 17.315 -132.655 ;
        RECT 18.125 -132.740 18.305 -132.470 ;
        RECT 18.125 -133.695 18.295 -132.740 ;
        RECT 18.615 -134.110 18.785 -132.655 ;
        RECT 19.675 -133.610 19.845 -132.655 ;
        RECT 20.140 -132.690 20.355 -132.270 ;
        RECT 19.650 -133.835 19.865 -133.610 ;
        RECT 20.165 -133.695 20.335 -132.690 ;
        RECT 21.220 -133.600 21.390 -132.655 ;
        RECT 21.685 -132.700 21.900 -132.270 ;
        RECT 19.170 -134.065 19.865 -133.835 ;
        RECT 15.980 -134.280 18.785 -134.110 ;
        RECT 15.980 -134.590 16.150 -134.280 ;
        RECT 12.770 -134.935 13.465 -134.665 ;
        RECT 15.420 -134.760 16.150 -134.590 ;
        RECT 15.420 -135.335 15.590 -134.760 ;
        RECT 16.515 -134.785 17.210 -134.515 ;
        RECT 11.655 -135.505 15.590 -135.335 ;
        RECT 15.895 -135.140 18.295 -134.970 ;
        RECT 8.720 -136.725 8.890 -135.770 ;
        RECT 0.275 -137.415 3.915 -137.245 ;
        RECT 12.775 -137.245 12.945 -135.685 ;
        RECT 13.265 -136.725 13.435 -135.505 ;
        RECT 13.755 -137.245 13.925 -135.685 ;
        RECT 14.355 -136.900 14.525 -135.685 ;
        RECT 14.845 -136.725 15.015 -135.505 ;
        RECT 15.335 -136.900 15.505 -135.685 ;
        RECT 15.895 -136.900 16.065 -135.140 ;
        RECT 14.355 -137.070 16.065 -136.900 ;
        RECT 16.245 -135.510 17.315 -135.340 ;
        RECT 16.245 -137.245 16.415 -135.510 ;
        RECT 17.145 -136.725 17.315 -135.510 ;
        RECT 18.125 -136.725 18.295 -135.140 ;
        RECT 18.560 -135.155 19.255 -134.885 ;
        RECT 19.650 -135.760 19.865 -134.065 ;
        RECT 21.200 -134.555 21.415 -133.600 ;
        RECT 21.710 -133.695 21.880 -132.700 ;
        RECT 27.755 -132.715 27.950 -132.100 ;
        RECT 28.265 -132.470 33.305 -132.290 ;
        RECT 33.680 -132.360 39.020 -132.100 ;
        RECT 26.155 -133.500 26.385 -132.820 ;
        RECT 20.700 -134.785 21.415 -134.555 ;
        RECT 19.675 -136.725 19.845 -135.760 ;
        RECT 21.200 -135.770 21.415 -134.785 ;
        RECT 21.635 -135.125 22.330 -134.855 ;
        RECT 26.185 -135.335 26.355 -133.500 ;
        RECT 27.775 -133.660 27.945 -132.715 ;
        RECT 27.765 -134.075 27.950 -133.660 ;
        RECT 28.265 -133.695 28.435 -132.470 ;
        RECT 29.845 -133.665 30.015 -132.655 ;
        RECT 30.335 -133.650 30.505 -132.655 ;
        RECT 31.655 -133.650 31.825 -132.655 ;
        RECT 29.830 -133.770 30.015 -133.665 ;
        RECT 29.235 -133.955 30.015 -133.770 ;
        RECT 30.325 -133.845 31.825 -133.650 ;
        RECT 29.235 -134.075 29.420 -133.955 ;
        RECT 27.765 -134.260 29.420 -134.075 ;
        RECT 32.145 -134.110 32.315 -132.655 ;
        RECT 33.125 -132.740 33.305 -132.470 ;
        RECT 33.125 -133.695 33.295 -132.740 ;
        RECT 33.615 -134.110 33.785 -132.655 ;
        RECT 34.675 -133.610 34.845 -132.655 ;
        RECT 35.140 -132.690 35.355 -132.360 ;
        RECT 34.650 -133.835 34.865 -133.610 ;
        RECT 35.165 -133.695 35.335 -132.690 ;
        RECT 36.220 -133.600 36.390 -132.655 ;
        RECT 36.685 -132.700 36.900 -132.360 ;
        RECT 34.170 -134.065 34.865 -133.835 ;
        RECT 30.980 -134.280 33.785 -134.110 ;
        RECT 30.980 -134.590 31.150 -134.280 ;
        RECT 27.770 -134.935 28.465 -134.665 ;
        RECT 30.420 -134.760 31.150 -134.590 ;
        RECT 30.420 -135.335 30.590 -134.760 ;
        RECT 31.515 -134.785 32.210 -134.515 ;
        RECT 26.185 -135.505 30.590 -135.335 ;
        RECT 30.895 -135.140 33.295 -134.970 ;
        RECT 21.220 -136.725 21.390 -135.770 ;
        RECT 12.775 -137.415 16.415 -137.245 ;
        RECT 27.775 -137.245 27.945 -135.685 ;
        RECT 28.265 -136.725 28.435 -135.505 ;
        RECT 28.755 -137.245 28.925 -135.685 ;
        RECT 29.355 -136.900 29.525 -135.685 ;
        RECT 29.845 -136.725 30.015 -135.505 ;
        RECT 30.335 -136.900 30.505 -135.685 ;
        RECT 30.895 -136.900 31.065 -135.140 ;
        RECT 29.355 -137.070 31.065 -136.900 ;
        RECT 31.245 -135.510 32.315 -135.340 ;
        RECT 31.245 -137.245 31.415 -135.510 ;
        RECT 32.145 -136.725 32.315 -135.510 ;
        RECT 33.125 -136.725 33.295 -135.140 ;
        RECT 33.560 -135.155 34.255 -134.885 ;
        RECT 34.650 -135.760 34.865 -134.065 ;
        RECT 36.200 -134.555 36.415 -133.600 ;
        RECT 36.710 -133.695 36.880 -132.700 ;
        RECT 35.700 -134.785 36.415 -134.555 ;
        RECT 34.675 -136.725 34.845 -135.760 ;
        RECT 36.200 -135.770 36.415 -134.785 ;
        RECT 36.635 -135.125 37.330 -134.855 ;
        RECT 36.220 -136.725 36.390 -135.770 ;
        RECT 27.775 -137.415 31.415 -137.245 ;
        RECT 44.545 -137.330 44.960 -128.005 ;
        RECT 45.730 -135.925 47.035 -127.025 ;
        RECT 60.810 -128.185 63.950 -128.015 ;
        RECT 53.350 -128.300 53.520 -128.280 ;
        RECT 53.320 -129.565 53.550 -128.300 ;
        RECT 54.330 -129.240 54.500 -128.280 ;
        RECT 55.310 -129.240 55.480 -128.280 ;
        RECT 57.760 -128.300 57.930 -128.280 ;
        RECT 56.655 -129.210 56.940 -128.390 ;
        RECT 54.300 -129.565 54.530 -129.240 ;
        RECT 55.280 -129.565 55.510 -129.240 ;
        RECT 53.320 -129.605 55.510 -129.565 ;
        RECT 57.730 -129.565 57.960 -128.300 ;
        RECT 58.740 -129.240 58.910 -128.280 ;
        RECT 59.720 -129.240 59.890 -128.280 ;
        RECT 60.810 -128.410 60.990 -128.185 ;
        RECT 58.710 -129.565 58.940 -129.240 ;
        RECT 59.690 -129.565 59.920 -129.240 ;
        RECT 57.730 -129.605 59.920 -129.565 ;
        RECT 60.195 -129.485 60.565 -128.645 ;
        RECT 60.815 -128.780 60.985 -128.410 ;
        RECT 60.195 -129.605 60.560 -129.485 ;
        RECT 52.300 -130.010 53.140 -129.640 ;
        RECT 53.320 -129.715 55.660 -129.605 ;
        RECT 56.710 -129.695 57.550 -129.640 ;
        RECT 55.950 -129.715 56.250 -129.695 ;
        RECT 56.535 -129.715 57.550 -129.695 ;
        RECT 53.320 -129.795 57.550 -129.715 ;
        RECT 49.295 -131.980 50.770 -131.490 ;
        RECT 52.400 -131.980 52.595 -130.010 ;
        RECT 52.860 -130.975 53.030 -130.180 ;
        RECT 53.320 -130.260 53.550 -129.795 ;
        RECT 53.350 -130.720 53.520 -130.260 ;
        RECT 53.840 -130.975 54.010 -130.180 ;
        RECT 54.300 -130.260 54.530 -129.795 ;
        RECT 55.280 -129.925 57.550 -129.795 ;
        RECT 55.280 -129.955 55.660 -129.925 ;
        RECT 54.330 -130.720 54.500 -130.260 ;
        RECT 54.820 -130.975 54.990 -130.180 ;
        RECT 55.280 -130.260 55.510 -129.955 ;
        RECT 55.310 -130.720 55.480 -130.260 ;
        RECT 55.950 -130.355 56.250 -129.925 ;
        RECT 56.535 -129.985 57.550 -129.925 ;
        RECT 56.710 -130.010 57.550 -129.985 ;
        RECT 57.730 -129.795 60.560 -129.605 ;
        RECT 57.270 -130.975 57.440 -130.180 ;
        RECT 57.730 -130.260 57.960 -129.795 ;
        RECT 57.760 -130.720 57.930 -130.260 ;
        RECT 58.250 -130.975 58.420 -130.180 ;
        RECT 58.710 -130.260 58.940 -129.795 ;
        RECT 59.690 -129.955 60.560 -129.795 ;
        RECT 60.785 -129.515 61.020 -128.780 ;
        RECT 61.305 -128.815 61.475 -128.355 ;
        RECT 61.790 -128.460 62.000 -128.185 ;
        RECT 61.300 -129.075 61.480 -128.815 ;
        RECT 61.795 -128.895 61.965 -128.460 ;
        RECT 62.285 -128.805 62.455 -128.355 ;
        RECT 62.760 -128.465 62.970 -128.185 ;
        RECT 62.285 -128.895 62.470 -128.805 ;
        RECT 62.775 -128.895 62.945 -128.465 ;
        RECT 63.265 -128.805 63.435 -128.355 ;
        RECT 63.740 -128.440 63.950 -128.185 ;
        RECT 74.310 -128.185 77.450 -128.015 ;
        RECT 66.475 -128.300 66.645 -128.280 ;
        RECT 62.290 -129.075 62.470 -128.895 ;
        RECT 63.260 -129.075 63.440 -128.805 ;
        RECT 63.755 -128.895 63.925 -128.440 ;
        RECT 64.245 -128.855 64.415 -128.355 ;
        RECT 64.230 -129.075 64.440 -128.855 ;
        RECT 61.300 -129.245 64.440 -129.075 ;
        RECT 60.785 -129.885 61.645 -129.515 ;
        RECT 63.565 -129.685 64.440 -129.245 ;
        RECT 66.445 -129.565 66.675 -128.300 ;
        RECT 67.455 -129.240 67.625 -128.280 ;
        RECT 68.435 -129.240 68.605 -128.280 ;
        RECT 71.260 -128.300 71.430 -128.280 ;
        RECT 70.155 -128.780 70.440 -128.390 ;
        RECT 69.135 -129.005 70.440 -128.780 ;
        RECT 67.425 -129.565 67.655 -129.240 ;
        RECT 68.405 -129.565 68.635 -129.240 ;
        RECT 66.445 -129.605 68.635 -129.565 ;
        RECT 65.425 -129.685 66.265 -129.640 ;
        RECT 58.740 -130.720 58.910 -130.260 ;
        RECT 59.230 -130.975 59.400 -130.180 ;
        RECT 59.690 -130.260 59.920 -129.955 ;
        RECT 59.720 -130.720 59.890 -130.260 ;
        RECT 60.785 -130.560 61.020 -129.885 ;
        RECT 63.565 -129.970 66.265 -129.685 ;
        RECT 63.565 -130.080 64.440 -129.970 ;
        RECT 65.425 -130.010 66.265 -129.970 ;
        RECT 66.445 -129.675 68.785 -129.605 ;
        RECT 69.135 -129.675 69.360 -129.005 ;
        RECT 70.155 -129.210 70.440 -129.005 ;
        RECT 71.230 -129.565 71.460 -128.300 ;
        RECT 72.240 -129.240 72.410 -128.280 ;
        RECT 73.220 -129.240 73.390 -128.280 ;
        RECT 74.310 -128.410 74.490 -128.185 ;
        RECT 72.210 -129.565 72.440 -129.240 ;
        RECT 73.190 -129.565 73.420 -129.240 ;
        RECT 71.230 -129.605 73.420 -129.565 ;
        RECT 73.695 -129.485 74.065 -128.645 ;
        RECT 74.315 -128.780 74.485 -128.410 ;
        RECT 73.695 -129.605 74.060 -129.485 ;
        RECT 66.445 -129.795 69.360 -129.675 ;
        RECT 61.285 -130.250 64.440 -130.080 ;
        RECT 61.285 -130.455 61.490 -130.250 ;
        RECT 60.815 -130.910 60.985 -130.560 ;
        RECT 52.815 -131.315 59.895 -130.975 ;
        RECT 60.790 -131.200 61.010 -130.910 ;
        RECT 61.305 -130.970 61.475 -130.455 ;
        RECT 61.795 -130.855 61.965 -130.430 ;
        RECT 62.275 -130.495 62.480 -130.250 ;
        RECT 61.770 -131.200 61.990 -130.855 ;
        RECT 62.285 -130.970 62.455 -130.495 ;
        RECT 62.775 -130.855 62.945 -130.430 ;
        RECT 63.245 -130.495 63.450 -130.250 ;
        RECT 64.230 -130.285 64.440 -130.250 ;
        RECT 62.750 -131.200 62.970 -130.855 ;
        RECT 63.265 -130.970 63.435 -130.495 ;
        RECT 63.755 -130.910 63.925 -130.430 ;
        RECT 64.230 -130.450 64.435 -130.285 ;
        RECT 64.200 -130.500 64.435 -130.450 ;
        RECT 63.735 -131.200 63.955 -130.910 ;
        RECT 64.200 -131.110 64.430 -130.500 ;
        RECT 65.985 -130.975 66.155 -130.180 ;
        RECT 66.445 -130.260 66.675 -129.795 ;
        RECT 66.475 -130.720 66.645 -130.260 ;
        RECT 66.965 -130.975 67.135 -130.180 ;
        RECT 67.425 -130.260 67.655 -129.795 ;
        RECT 68.405 -129.900 69.360 -129.795 ;
        RECT 69.610 -129.695 69.910 -129.690 ;
        RECT 70.210 -129.695 71.050 -129.640 ;
        RECT 68.405 -129.955 68.785 -129.900 ;
        RECT 67.455 -130.720 67.625 -130.260 ;
        RECT 67.945 -130.975 68.115 -130.180 ;
        RECT 68.405 -130.260 68.635 -129.955 ;
        RECT 68.435 -130.720 68.605 -130.260 ;
        RECT 69.035 -130.475 69.335 -129.900 ;
        RECT 69.610 -129.985 71.050 -129.695 ;
        RECT 69.610 -130.350 69.910 -129.985 ;
        RECT 70.210 -130.010 71.050 -129.985 ;
        RECT 71.230 -129.795 74.060 -129.605 ;
        RECT 70.770 -130.975 70.940 -130.180 ;
        RECT 71.230 -130.260 71.460 -129.795 ;
        RECT 71.260 -130.720 71.430 -130.260 ;
        RECT 71.750 -130.975 71.920 -130.180 ;
        RECT 72.210 -130.260 72.440 -129.795 ;
        RECT 73.190 -129.955 74.060 -129.795 ;
        RECT 74.285 -129.515 74.520 -128.780 ;
        RECT 74.805 -128.815 74.975 -128.355 ;
        RECT 75.290 -128.460 75.500 -128.185 ;
        RECT 74.800 -129.075 74.980 -128.815 ;
        RECT 75.295 -128.895 75.465 -128.460 ;
        RECT 75.785 -128.805 75.955 -128.355 ;
        RECT 76.260 -128.465 76.470 -128.185 ;
        RECT 75.785 -128.895 75.970 -128.805 ;
        RECT 76.275 -128.895 76.445 -128.465 ;
        RECT 76.765 -128.805 76.935 -128.355 ;
        RECT 77.240 -128.440 77.450 -128.185 ;
        RECT 79.975 -128.300 80.145 -128.280 ;
        RECT 75.790 -129.075 75.970 -128.895 ;
        RECT 76.760 -129.075 76.940 -128.805 ;
        RECT 77.255 -128.895 77.425 -128.440 ;
        RECT 77.745 -128.855 77.915 -128.355 ;
        RECT 77.730 -129.075 77.940 -128.855 ;
        RECT 74.800 -129.245 77.940 -129.075 ;
        RECT 74.285 -129.885 75.145 -129.515 ;
        RECT 77.065 -129.670 77.940 -129.245 ;
        RECT 79.945 -129.565 80.175 -128.300 ;
        RECT 80.955 -129.240 81.125 -128.280 ;
        RECT 81.935 -129.240 82.105 -128.280 ;
        RECT 80.925 -129.565 81.155 -129.240 ;
        RECT 81.905 -129.565 82.135 -129.240 ;
        RECT 79.945 -129.605 82.135 -129.565 ;
        RECT 78.925 -129.670 79.765 -129.640 ;
        RECT 72.240 -130.720 72.410 -130.260 ;
        RECT 72.730 -130.975 72.900 -130.180 ;
        RECT 73.190 -130.260 73.420 -129.955 ;
        RECT 73.220 -130.720 73.390 -130.260 ;
        RECT 74.285 -130.560 74.520 -129.885 ;
        RECT 77.065 -129.935 79.765 -129.670 ;
        RECT 77.065 -130.080 77.940 -129.935 ;
        RECT 78.925 -130.010 79.765 -129.935 ;
        RECT 79.945 -129.650 82.285 -129.605 ;
        RECT 79.945 -129.660 82.695 -129.650 ;
        RECT 79.945 -129.795 82.700 -129.660 ;
        RECT 74.785 -130.250 77.940 -130.080 ;
        RECT 74.785 -130.455 74.990 -130.250 ;
        RECT 74.315 -130.910 74.485 -130.560 ;
        RECT 60.790 -131.370 63.955 -131.200 ;
        RECT 65.940 -131.315 73.395 -130.975 ;
        RECT 74.290 -131.200 74.510 -130.910 ;
        RECT 74.805 -130.970 74.975 -130.455 ;
        RECT 75.295 -130.855 75.465 -130.430 ;
        RECT 75.775 -130.495 75.980 -130.250 ;
        RECT 75.270 -131.200 75.490 -130.855 ;
        RECT 75.785 -130.970 75.955 -130.495 ;
        RECT 76.275 -130.855 76.445 -130.430 ;
        RECT 76.745 -130.495 76.950 -130.250 ;
        RECT 77.730 -130.285 77.940 -130.250 ;
        RECT 76.250 -131.200 76.470 -130.855 ;
        RECT 76.765 -130.970 76.935 -130.495 ;
        RECT 77.255 -130.910 77.425 -130.430 ;
        RECT 77.730 -130.500 77.935 -130.285 ;
        RECT 77.235 -131.200 77.455 -130.910 ;
        RECT 77.745 -130.970 77.915 -130.500 ;
        RECT 79.485 -130.975 79.655 -130.180 ;
        RECT 79.945 -130.260 80.175 -129.795 ;
        RECT 79.975 -130.720 80.145 -130.260 ;
        RECT 80.465 -130.975 80.635 -130.180 ;
        RECT 80.925 -130.260 81.155 -129.795 ;
        RECT 81.905 -129.845 82.700 -129.795 ;
        RECT 81.905 -129.955 82.285 -129.845 ;
        RECT 80.955 -130.720 81.125 -130.260 ;
        RECT 81.445 -130.975 81.615 -130.180 ;
        RECT 81.905 -130.260 82.135 -129.955 ;
        RECT 81.935 -130.720 82.105 -130.260 ;
        RECT 74.290 -131.370 77.455 -131.200 ;
        RECT 79.440 -131.315 82.110 -130.975 ;
        RECT 55.745 -131.550 56.405 -131.495 ;
        RECT 78.360 -131.550 79.020 -131.485 ;
        RECT 55.745 -131.745 81.050 -131.550 ;
        RECT 82.460 -131.635 82.700 -129.845 ;
        RECT 55.745 -131.795 56.405 -131.745 ;
        RECT 78.360 -131.785 79.020 -131.745 ;
        RECT 64.765 -131.980 65.425 -131.925 ;
        RECT 69.470 -131.980 70.155 -131.930 ;
        RECT 49.295 -132.175 81.050 -131.980 ;
        RECT 49.295 -132.505 50.770 -132.175 ;
        RECT 64.765 -132.225 65.425 -132.175 ;
        RECT 69.470 -132.230 70.155 -132.175 ;
        RECT 82.405 -132.320 82.705 -131.635 ;
        RECT 54.130 -132.440 54.790 -132.345 ;
        RECT 67.295 -132.440 67.980 -132.345 ;
        RECT 80.280 -132.440 80.965 -132.375 ;
        RECT 54.125 -132.635 81.050 -132.440 ;
        RECT 54.130 -132.645 55.955 -132.635 ;
        RECT 54.650 -135.925 55.955 -132.645 ;
        RECT 57.735 -132.990 60.900 -132.820 ;
        RECT 62.920 -132.875 63.475 -132.635 ;
        RECT 67.295 -132.645 67.980 -132.635 ;
        RECT 64.350 -132.875 66.950 -132.865 ;
        RECT 67.310 -132.875 67.865 -132.645 ;
        RECT 57.275 -133.690 57.445 -133.220 ;
        RECT 57.735 -133.280 57.955 -132.990 ;
        RECT 57.255 -133.905 57.460 -133.690 ;
        RECT 57.765 -133.760 57.935 -133.280 ;
        RECT 58.255 -133.695 58.425 -133.220 ;
        RECT 58.720 -133.335 58.940 -132.990 ;
        RECT 57.250 -133.940 57.460 -133.905 ;
        RECT 58.240 -133.940 58.445 -133.695 ;
        RECT 58.745 -133.760 58.915 -133.335 ;
        RECT 59.235 -133.695 59.405 -133.220 ;
        RECT 59.700 -133.335 59.920 -132.990 ;
        RECT 59.210 -133.940 59.415 -133.695 ;
        RECT 59.725 -133.760 59.895 -133.335 ;
        RECT 60.215 -133.735 60.385 -133.220 ;
        RECT 60.680 -133.280 60.900 -132.990 ;
        RECT 61.795 -133.205 68.650 -132.875 ;
        RECT 61.795 -133.215 64.465 -133.205 ;
        RECT 65.980 -133.215 68.650 -133.205 ;
        RECT 71.235 -132.990 74.400 -132.820 ;
        RECT 76.300 -132.875 76.855 -132.635 ;
        RECT 80.280 -132.675 80.965 -132.635 ;
        RECT 80.355 -132.875 80.910 -132.675 ;
        RECT 60.705 -133.630 60.875 -133.280 ;
        RECT 60.200 -133.940 60.405 -133.735 ;
        RECT 57.250 -134.100 60.405 -133.940 ;
        RECT 56.875 -134.110 60.405 -134.100 ;
        RECT 56.875 -134.400 58.125 -134.110 ;
        RECT 60.670 -134.305 60.905 -133.630 ;
        RECT 61.800 -133.930 61.970 -133.470 ;
        RECT 61.770 -134.235 62.000 -133.930 ;
        RECT 62.290 -134.010 62.460 -133.215 ;
        RECT 62.780 -133.930 62.950 -133.470 ;
        RECT 57.250 -134.945 58.125 -134.400 ;
        RECT 60.045 -134.675 60.905 -134.305 ;
        RECT 57.250 -135.115 60.390 -134.945 ;
        RECT 57.250 -135.335 57.460 -135.115 ;
        RECT 57.275 -135.835 57.445 -135.335 ;
        RECT 57.765 -135.750 57.935 -135.295 ;
        RECT 58.250 -135.385 58.430 -135.115 ;
        RECT 59.220 -135.295 59.400 -135.115 ;
        RECT 45.730 -137.230 55.955 -135.925 ;
        RECT 57.740 -136.005 57.950 -135.750 ;
        RECT 58.255 -135.835 58.425 -135.385 ;
        RECT 58.745 -135.725 58.915 -135.295 ;
        RECT 59.220 -135.385 59.405 -135.295 ;
        RECT 58.720 -136.005 58.930 -135.725 ;
        RECT 59.235 -135.835 59.405 -135.385 ;
        RECT 59.725 -135.730 59.895 -135.295 ;
        RECT 60.210 -135.375 60.390 -135.115 ;
        RECT 59.690 -136.005 59.900 -135.730 ;
        RECT 60.215 -135.835 60.385 -135.375 ;
        RECT 60.670 -135.410 60.905 -134.675 ;
        RECT 61.130 -134.395 62.000 -134.235 ;
        RECT 62.750 -134.395 62.980 -133.930 ;
        RECT 63.270 -134.010 63.440 -133.215 ;
        RECT 63.760 -133.930 63.930 -133.470 ;
        RECT 63.730 -134.395 63.960 -133.930 ;
        RECT 64.250 -134.010 64.420 -133.215 ;
        RECT 64.980 -134.180 65.280 -133.385 ;
        RECT 65.985 -133.930 66.155 -133.470 ;
        RECT 61.130 -134.585 63.960 -134.395 ;
        RECT 64.140 -134.495 65.280 -134.180 ;
        RECT 65.955 -134.235 66.185 -133.930 ;
        RECT 66.475 -134.010 66.645 -133.215 ;
        RECT 66.965 -133.930 67.135 -133.470 ;
        RECT 65.465 -134.395 66.185 -134.235 ;
        RECT 66.935 -134.395 67.165 -133.930 ;
        RECT 67.455 -134.010 67.625 -133.215 ;
        RECT 67.945 -133.930 68.115 -133.470 ;
        RECT 67.915 -134.395 68.145 -133.930 ;
        RECT 68.435 -134.010 68.605 -133.215 ;
        RECT 70.775 -133.690 70.945 -133.220 ;
        RECT 71.235 -133.280 71.455 -132.990 ;
        RECT 70.755 -133.905 70.960 -133.690 ;
        RECT 71.265 -133.760 71.435 -133.280 ;
        RECT 71.755 -133.695 71.925 -133.220 ;
        RECT 72.220 -133.335 72.440 -132.990 ;
        RECT 70.750 -133.940 70.960 -133.905 ;
        RECT 71.740 -133.940 71.945 -133.695 ;
        RECT 72.245 -133.760 72.415 -133.335 ;
        RECT 72.735 -133.695 72.905 -133.220 ;
        RECT 73.200 -133.335 73.420 -132.990 ;
        RECT 72.710 -133.940 72.915 -133.695 ;
        RECT 73.225 -133.760 73.395 -133.335 ;
        RECT 73.715 -133.735 73.885 -133.220 ;
        RECT 74.180 -133.280 74.400 -132.990 ;
        RECT 75.295 -133.215 82.150 -132.875 ;
        RECT 74.205 -133.630 74.375 -133.280 ;
        RECT 73.700 -133.940 73.905 -133.735 ;
        RECT 70.750 -134.110 73.905 -133.940 ;
        RECT 64.140 -134.550 64.980 -134.495 ;
        RECT 61.130 -134.705 61.495 -134.585 ;
        RECT 60.705 -135.780 60.875 -135.410 ;
        RECT 61.125 -135.545 61.495 -134.705 ;
        RECT 61.770 -134.625 63.960 -134.585 ;
        RECT 61.770 -134.950 62.000 -134.625 ;
        RECT 62.750 -134.950 62.980 -134.625 ;
        RECT 60.700 -136.005 60.880 -135.780 ;
        RECT 61.800 -135.910 61.970 -134.950 ;
        RECT 62.780 -135.910 62.950 -134.950 ;
        RECT 63.730 -135.890 63.960 -134.625 ;
        RECT 65.465 -134.585 68.145 -134.395 ;
        RECT 68.325 -134.215 69.165 -134.180 ;
        RECT 68.325 -134.515 69.275 -134.215 ;
        RECT 70.295 -134.410 71.625 -134.110 ;
        RECT 74.170 -134.305 74.405 -133.630 ;
        RECT 75.300 -133.930 75.470 -133.470 ;
        RECT 75.270 -134.235 75.500 -133.930 ;
        RECT 75.790 -134.010 75.960 -133.215 ;
        RECT 76.280 -133.930 76.450 -133.470 ;
        RECT 68.325 -134.550 69.165 -134.515 ;
        RECT 64.750 -135.230 65.035 -134.980 ;
        RECT 65.465 -135.230 65.775 -134.585 ;
        RECT 65.955 -134.625 68.145 -134.585 ;
        RECT 65.955 -134.950 66.185 -134.625 ;
        RECT 66.935 -134.950 67.165 -134.625 ;
        RECT 64.750 -135.540 65.775 -135.230 ;
        RECT 64.750 -135.800 65.035 -135.540 ;
        RECT 63.760 -135.910 63.930 -135.890 ;
        RECT 65.985 -135.910 66.155 -134.950 ;
        RECT 66.965 -135.910 67.135 -134.950 ;
        RECT 67.915 -135.890 68.145 -134.625 ;
        RECT 70.750 -134.945 71.625 -134.410 ;
        RECT 73.545 -134.675 74.405 -134.305 ;
        RECT 70.750 -135.115 73.890 -134.945 ;
        RECT 70.750 -135.335 70.960 -135.115 ;
        RECT 70.775 -135.835 70.945 -135.335 ;
        RECT 71.265 -135.750 71.435 -135.295 ;
        RECT 71.750 -135.385 71.930 -135.115 ;
        RECT 72.720 -135.295 72.900 -135.115 ;
        RECT 67.945 -135.910 68.115 -135.890 ;
        RECT 57.740 -136.175 60.880 -136.005 ;
        RECT 71.240 -136.005 71.450 -135.750 ;
        RECT 71.755 -135.835 71.925 -135.385 ;
        RECT 72.245 -135.725 72.415 -135.295 ;
        RECT 72.720 -135.385 72.905 -135.295 ;
        RECT 72.220 -136.005 72.430 -135.725 ;
        RECT 72.735 -135.835 72.905 -135.385 ;
        RECT 73.225 -135.730 73.395 -135.295 ;
        RECT 73.710 -135.375 73.890 -135.115 ;
        RECT 73.190 -136.005 73.400 -135.730 ;
        RECT 73.715 -135.835 73.885 -135.375 ;
        RECT 74.170 -135.410 74.405 -134.675 ;
        RECT 74.630 -134.395 75.500 -134.235 ;
        RECT 76.250 -134.395 76.480 -133.930 ;
        RECT 76.770 -134.010 76.940 -133.215 ;
        RECT 77.260 -133.930 77.430 -133.470 ;
        RECT 77.230 -134.395 77.460 -133.930 ;
        RECT 77.750 -134.010 77.920 -133.215 ;
        RECT 78.540 -134.180 78.840 -133.460 ;
        RECT 79.485 -133.930 79.655 -133.470 ;
        RECT 74.630 -134.585 77.460 -134.395 ;
        RECT 77.640 -134.490 78.840 -134.180 ;
        RECT 79.455 -134.235 79.685 -133.930 ;
        RECT 79.975 -134.010 80.145 -133.215 ;
        RECT 80.465 -133.930 80.635 -133.470 ;
        RECT 79.020 -134.395 79.685 -134.235 ;
        RECT 80.435 -134.395 80.665 -133.930 ;
        RECT 80.955 -134.010 81.125 -133.215 ;
        RECT 81.445 -133.930 81.615 -133.470 ;
        RECT 81.415 -134.395 81.645 -133.930 ;
        RECT 81.935 -134.010 82.105 -133.215 ;
        RECT 82.460 -134.180 82.700 -132.320 ;
        RECT 77.640 -134.495 78.655 -134.490 ;
        RECT 77.640 -134.550 78.480 -134.495 ;
        RECT 74.630 -134.705 74.995 -134.585 ;
        RECT 74.205 -135.780 74.375 -135.410 ;
        RECT 74.625 -135.545 74.995 -134.705 ;
        RECT 75.270 -134.625 77.460 -134.585 ;
        RECT 75.270 -134.950 75.500 -134.625 ;
        RECT 76.250 -134.950 76.480 -134.625 ;
        RECT 74.200 -136.005 74.380 -135.780 ;
        RECT 75.300 -135.910 75.470 -134.950 ;
        RECT 76.280 -135.910 76.450 -134.950 ;
        RECT 77.230 -135.890 77.460 -134.625 ;
        RECT 79.020 -134.585 81.645 -134.395 ;
        RECT 81.825 -134.400 82.700 -134.180 ;
        RECT 81.825 -134.550 82.665 -134.400 ;
        RECT 78.250 -135.235 78.535 -134.980 ;
        RECT 79.020 -135.235 79.250 -134.585 ;
        RECT 79.455 -134.625 81.645 -134.585 ;
        RECT 79.455 -134.950 79.685 -134.625 ;
        RECT 80.435 -134.950 80.665 -134.625 ;
        RECT 78.250 -135.480 79.250 -135.235 ;
        RECT 78.250 -135.800 78.535 -135.480 ;
        RECT 77.260 -135.910 77.430 -135.890 ;
        RECT 79.485 -135.910 79.655 -134.950 ;
        RECT 80.465 -135.910 80.635 -134.950 ;
        RECT 81.415 -135.890 81.645 -134.625 ;
        RECT 129.445 -135.685 130.175 -116.935 ;
        RECT 133.425 -117.775 133.805 -116.935 ;
        RECT 133.425 -118.155 134.135 -117.775 ;
        RECT 133.755 -120.100 134.135 -118.155 ;
        RECT 138.800 -117.985 142.125 -117.845 ;
        RECT 138.800 -118.275 143.975 -117.985 ;
        RECT 147.845 -118.270 148.305 -117.845 ;
        RECT 138.800 -118.680 139.230 -118.275 ;
        RECT 140.100 -118.460 140.275 -118.275 ;
        RECT 141.725 -118.290 143.975 -118.275 ;
        RECT 134.540 -119.110 139.230 -118.680 ;
        RECT 133.755 -120.560 134.430 -120.100 ;
        RECT 135.240 -120.390 135.410 -119.110 ;
        RECT 135.730 -120.390 135.900 -119.350 ;
        RECT 136.220 -120.390 136.390 -119.110 ;
        RECT 136.710 -120.220 136.880 -119.350 ;
        RECT 139.615 -120.000 139.785 -118.460 ;
        RECT 140.105 -120.000 140.275 -118.460 ;
        RECT 140.595 -120.000 140.765 -118.460 ;
        RECT 141.085 -120.000 141.255 -118.460 ;
        RECT 141.575 -120.000 141.745 -118.460 ;
        RECT 139.455 -120.215 139.810 -120.210 ;
        RECT 141.515 -120.215 141.885 -120.185 ;
        RECT 139.455 -120.220 141.885 -120.215 ;
        RECT 136.710 -120.390 141.885 -120.220 ;
        RECT 143.670 -120.325 143.975 -118.290 ;
        RECT 136.715 -120.410 141.885 -120.390 ;
        RECT 136.715 -120.420 139.460 -120.410 ;
        RECT 134.650 -120.560 135.015 -120.530 ;
        RECT 141.515 -120.540 141.885 -120.410 ;
        RECT 133.755 -120.645 135.015 -120.560 ;
        RECT 133.780 -120.765 135.015 -120.645 ;
        RECT 139.190 -120.700 139.865 -120.660 ;
        RECT 139.090 -120.710 139.865 -120.700 ;
        RECT 133.780 -120.850 134.430 -120.765 ;
        RECT 134.650 -120.830 135.015 -120.765 ;
        RECT 138.055 -120.890 139.865 -120.710 ;
        RECT 142.450 -120.755 146.375 -120.325 ;
        RECT 139.090 -120.900 139.865 -120.890 ;
        RECT 139.190 -120.930 139.865 -120.900 ;
        RECT 140.105 -120.815 142.200 -120.775 ;
        RECT 140.105 -120.965 142.255 -120.815 ;
        RECT 135.240 -122.040 135.410 -121.000 ;
        RECT 136.220 -122.040 136.390 -121.000 ;
        RECT 137.200 -122.040 137.370 -121.000 ;
        RECT 140.105 -122.685 140.275 -120.965 ;
        RECT 141.085 -122.685 141.255 -120.965 ;
        RECT 141.950 -121.710 142.255 -120.965 ;
        RECT 143.150 -121.535 143.320 -120.755 ;
        RECT 143.640 -121.535 143.810 -120.995 ;
        RECT 144.130 -121.535 144.300 -120.755 ;
        RECT 144.620 -121.535 144.790 -120.995 ;
        RECT 142.560 -121.710 142.925 -121.680 ;
        RECT 141.950 -121.775 142.925 -121.710 ;
        RECT 142.060 -121.915 142.925 -121.775 ;
        RECT 142.560 -121.980 142.925 -121.915 ;
        RECT 145.110 -121.830 146.970 -121.480 ;
        RECT 143.150 -122.690 143.320 -122.150 ;
        RECT 144.130 -122.690 144.300 -122.150 ;
        RECT 145.110 -122.690 145.280 -121.830 ;
        RECT 143.380 -125.030 144.580 -124.860 ;
        RECT 135.110 -127.365 135.280 -125.645 ;
        RECT 136.090 -127.365 136.260 -125.645 ;
        RECT 138.155 -126.180 138.325 -125.640 ;
        RECT 139.135 -126.180 139.305 -125.640 ;
        RECT 137.565 -126.415 137.930 -126.350 ;
        RECT 137.065 -126.555 137.930 -126.415 ;
        RECT 136.955 -126.620 137.930 -126.555 ;
        RECT 136.955 -127.365 137.260 -126.620 ;
        RECT 137.565 -126.650 137.930 -126.620 ;
        RECT 140.115 -126.500 140.285 -125.640 ;
        RECT 135.110 -127.515 137.260 -127.365 ;
        RECT 135.110 -127.555 137.205 -127.515 ;
        RECT 138.155 -127.575 138.325 -126.795 ;
        RECT 138.645 -127.335 138.815 -126.795 ;
        RECT 139.135 -127.575 139.305 -126.795 ;
        RECT 139.625 -127.335 139.795 -126.795 ;
        RECT 140.115 -126.850 141.505 -126.500 ;
        RECT 133.330 -127.920 134.465 -127.910 ;
        RECT 136.520 -127.920 136.890 -127.790 ;
        RECT 133.330 -128.110 136.890 -127.920 ;
        RECT 137.455 -128.005 140.530 -127.575 ;
        RECT 134.460 -128.115 136.890 -128.110 ;
        RECT 134.460 -128.120 134.815 -128.115 ;
        RECT 136.520 -128.145 136.890 -128.115 ;
        RECT 134.620 -129.870 134.790 -128.330 ;
        RECT 135.110 -129.870 135.280 -128.330 ;
        RECT 135.600 -129.870 135.770 -128.330 ;
        RECT 136.090 -129.870 136.260 -128.330 ;
        RECT 136.580 -129.870 136.750 -128.330 ;
        RECT 135.105 -130.130 135.280 -129.870 ;
        RECT 138.675 -130.040 138.980 -128.005 ;
        RECT 141.125 -128.825 141.475 -126.850 ;
        RECT 142.345 -128.120 142.515 -125.200 ;
        RECT 143.380 -125.240 143.590 -125.030 ;
        RECT 142.325 -128.415 142.535 -128.120 ;
        RECT 143.400 -128.150 143.570 -125.240 ;
        RECT 143.890 -128.140 144.060 -125.200 ;
        RECT 144.370 -125.250 144.580 -125.030 ;
        RECT 143.385 -128.415 143.595 -128.150 ;
        RECT 142.325 -128.595 143.595 -128.415 ;
        RECT 143.870 -128.410 144.080 -128.140 ;
        RECT 144.380 -128.240 144.550 -125.250 ;
        RECT 145.440 -128.170 145.610 -125.200 ;
        RECT 143.870 -128.605 144.575 -128.410 ;
        RECT 144.360 -128.665 144.575 -128.605 ;
        RECT 143.150 -128.825 143.925 -128.775 ;
        RECT 141.125 -129.005 143.925 -128.825 ;
        RECT 141.125 -129.015 141.475 -129.005 ;
        RECT 143.150 -129.050 143.925 -129.005 ;
        RECT 144.360 -128.940 145.265 -128.665 ;
        RECT 144.360 -129.290 144.575 -128.940 ;
        RECT 141.800 -129.360 142.575 -129.315 ;
        RECT 141.615 -129.530 142.575 -129.360 ;
        RECT 141.800 -129.590 142.575 -129.530 ;
        RECT 142.805 -129.490 144.575 -129.290 ;
        RECT 145.435 -129.390 145.650 -128.170 ;
        RECT 146.620 -128.515 146.970 -121.830 ;
        RECT 147.960 -128.145 148.175 -118.270 ;
        RECT 149.595 -120.385 149.975 -116.865 ;
        RECT 151.105 -116.645 160.040 -116.455 ;
        RECT 151.105 -118.535 151.295 -116.645 ;
        RECT 157.140 -118.140 160.465 -118.000 ;
        RECT 157.140 -118.430 162.315 -118.140 ;
        RECT 150.990 -118.805 151.355 -118.535 ;
        RECT 157.140 -118.835 157.570 -118.430 ;
        RECT 158.440 -118.615 158.615 -118.430 ;
        RECT 160.065 -118.445 162.315 -118.430 ;
        RECT 152.880 -119.265 157.570 -118.835 ;
        RECT 152.120 -120.385 152.770 -120.255 ;
        RECT 149.595 -120.715 152.770 -120.385 ;
        RECT 153.580 -120.545 153.750 -119.265 ;
        RECT 154.070 -120.545 154.240 -119.505 ;
        RECT 154.560 -120.545 154.730 -119.265 ;
        RECT 155.050 -120.375 155.220 -119.505 ;
        RECT 157.955 -120.155 158.125 -118.615 ;
        RECT 158.445 -120.155 158.615 -118.615 ;
        RECT 158.935 -120.155 159.105 -118.615 ;
        RECT 159.425 -120.155 159.595 -118.615 ;
        RECT 159.915 -120.155 160.085 -118.615 ;
        RECT 157.795 -120.370 158.150 -120.365 ;
        RECT 159.855 -120.370 160.225 -120.340 ;
        RECT 157.795 -120.375 160.225 -120.370 ;
        RECT 155.050 -120.545 160.225 -120.375 ;
        RECT 162.010 -120.480 162.315 -118.445 ;
        RECT 155.055 -120.565 160.225 -120.545 ;
        RECT 155.055 -120.575 157.800 -120.565 ;
        RECT 152.990 -120.715 153.355 -120.685 ;
        RECT 159.855 -120.695 160.225 -120.565 ;
        RECT 149.595 -120.765 153.355 -120.715 ;
        RECT 152.120 -120.920 153.355 -120.765 ;
        RECT 157.530 -120.855 158.205 -120.815 ;
        RECT 157.430 -120.865 158.205 -120.855 ;
        RECT 152.120 -121.005 152.770 -120.920 ;
        RECT 152.990 -120.985 153.355 -120.920 ;
        RECT 152.255 -121.255 152.635 -121.005 ;
        RECT 156.395 -121.045 158.205 -120.865 ;
        RECT 160.790 -120.910 164.715 -120.480 ;
        RECT 157.430 -121.055 158.205 -121.045 ;
        RECT 157.530 -121.085 158.205 -121.055 ;
        RECT 158.445 -120.970 160.540 -120.930 ;
        RECT 158.445 -121.120 160.595 -120.970 ;
        RECT 153.580 -122.195 153.750 -121.155 ;
        RECT 154.560 -122.195 154.730 -121.155 ;
        RECT 155.540 -122.195 155.710 -121.155 ;
        RECT 158.445 -122.840 158.615 -121.120 ;
        RECT 159.425 -122.840 159.595 -121.120 ;
        RECT 160.290 -121.865 160.595 -121.120 ;
        RECT 161.490 -121.690 161.660 -120.910 ;
        RECT 161.980 -121.690 162.150 -121.150 ;
        RECT 162.470 -121.690 162.640 -120.910 ;
        RECT 162.960 -121.690 163.130 -121.150 ;
        RECT 160.900 -121.865 161.265 -121.835 ;
        RECT 160.290 -121.930 161.265 -121.865 ;
        RECT 160.400 -122.070 161.265 -121.930 ;
        RECT 160.900 -122.135 161.265 -122.070 ;
        RECT 163.450 -121.985 165.310 -121.635 ;
        RECT 161.490 -122.845 161.660 -122.305 ;
        RECT 162.470 -122.845 162.640 -122.305 ;
        RECT 163.450 -122.845 163.620 -121.985 ;
        RECT 161.720 -125.185 162.920 -125.015 ;
        RECT 153.450 -127.520 153.620 -125.800 ;
        RECT 154.430 -127.520 154.600 -125.800 ;
        RECT 156.495 -126.335 156.665 -125.795 ;
        RECT 157.475 -126.335 157.645 -125.795 ;
        RECT 155.905 -126.570 156.270 -126.505 ;
        RECT 155.405 -126.710 156.270 -126.570 ;
        RECT 155.295 -126.775 156.270 -126.710 ;
        RECT 155.295 -127.520 155.600 -126.775 ;
        RECT 155.905 -126.805 156.270 -126.775 ;
        RECT 158.455 -126.655 158.625 -125.795 ;
        RECT 153.450 -127.670 155.600 -127.520 ;
        RECT 153.450 -127.710 155.545 -127.670 ;
        RECT 156.495 -127.730 156.665 -126.950 ;
        RECT 156.985 -127.490 157.155 -126.950 ;
        RECT 157.475 -127.730 157.645 -126.950 ;
        RECT 157.965 -127.490 158.135 -126.950 ;
        RECT 158.455 -127.005 159.845 -126.655 ;
        RECT 151.670 -128.075 152.805 -128.065 ;
        RECT 154.860 -128.075 155.230 -127.945 ;
        RECT 147.960 -128.360 149.385 -128.145 ;
        RECT 151.670 -128.265 155.230 -128.075 ;
        RECT 155.795 -128.160 158.870 -127.730 ;
        RECT 152.800 -128.270 155.230 -128.265 ;
        RECT 152.800 -128.275 153.155 -128.270 ;
        RECT 154.860 -128.300 155.230 -128.270 ;
        RECT 146.565 -128.875 147.090 -128.515 ;
        RECT 149.170 -129.390 149.385 -128.360 ;
        RECT 136.730 -130.130 138.980 -130.040 ;
        RECT 134.520 -130.345 138.980 -130.130 ;
        RECT 134.520 -130.435 136.765 -130.345 ;
        RECT 138.675 -131.820 138.980 -130.345 ;
        RECT 142.345 -131.230 142.515 -129.760 ;
        RECT 142.805 -129.840 143.030 -129.490 ;
        RECT 144.765 -129.590 149.385 -129.390 ;
        RECT 145.005 -129.605 149.385 -129.590 ;
        RECT 142.310 -131.820 142.545 -131.230 ;
        RECT 142.835 -131.300 143.005 -129.840 ;
        RECT 143.325 -131.225 143.495 -129.760 ;
        RECT 144.535 -131.175 144.705 -129.760 ;
        RECT 145.005 -129.805 145.225 -129.605 ;
        RECT 143.290 -131.820 143.525 -131.225 ;
        RECT 144.500 -131.820 144.735 -131.175 ;
        RECT 145.025 -131.300 145.195 -129.805 ;
        RECT 152.960 -130.025 153.130 -128.485 ;
        RECT 153.450 -130.025 153.620 -128.485 ;
        RECT 153.940 -130.025 154.110 -128.485 ;
        RECT 154.430 -130.025 154.600 -128.485 ;
        RECT 154.920 -130.025 155.090 -128.485 ;
        RECT 153.445 -130.285 153.620 -130.025 ;
        RECT 157.015 -130.195 157.320 -128.160 ;
        RECT 159.465 -128.980 159.815 -127.005 ;
        RECT 160.685 -128.275 160.855 -125.355 ;
        RECT 161.720 -125.395 161.930 -125.185 ;
        RECT 160.665 -128.570 160.875 -128.275 ;
        RECT 161.740 -128.305 161.910 -125.395 ;
        RECT 162.230 -128.295 162.400 -125.355 ;
        RECT 162.710 -125.405 162.920 -125.185 ;
        RECT 161.725 -128.570 161.935 -128.305 ;
        RECT 160.665 -128.750 161.935 -128.570 ;
        RECT 162.210 -128.565 162.420 -128.295 ;
        RECT 162.720 -128.395 162.890 -125.405 ;
        RECT 163.780 -128.325 163.950 -125.355 ;
        RECT 162.210 -128.760 162.915 -128.565 ;
        RECT 162.700 -128.820 162.915 -128.760 ;
        RECT 161.490 -128.980 162.265 -128.930 ;
        RECT 159.465 -129.160 162.265 -128.980 ;
        RECT 159.465 -129.170 159.815 -129.160 ;
        RECT 161.490 -129.205 162.265 -129.160 ;
        RECT 162.700 -129.095 163.605 -128.820 ;
        RECT 162.700 -129.445 162.915 -129.095 ;
        RECT 160.140 -129.515 160.915 -129.470 ;
        RECT 159.955 -129.685 160.915 -129.515 ;
        RECT 160.140 -129.745 160.915 -129.685 ;
        RECT 161.145 -129.645 162.915 -129.445 ;
        RECT 163.775 -129.545 163.990 -128.325 ;
        RECT 164.960 -128.670 165.310 -121.985 ;
        RECT 164.905 -129.030 165.430 -128.670 ;
        RECT 167.435 -129.545 168.550 -129.095 ;
        RECT 155.070 -130.285 157.320 -130.195 ;
        RECT 152.860 -130.500 157.320 -130.285 ;
        RECT 152.860 -130.590 155.105 -130.500 ;
        RECT 138.675 -132.385 146.060 -131.820 ;
        RECT 157.015 -131.975 157.320 -130.500 ;
        RECT 160.685 -131.385 160.855 -129.915 ;
        RECT 161.145 -129.995 161.370 -129.645 ;
        RECT 163.105 -129.745 169.115 -129.545 ;
        RECT 163.345 -129.760 169.115 -129.745 ;
        RECT 160.650 -131.975 160.885 -131.385 ;
        RECT 161.175 -131.455 161.345 -129.995 ;
        RECT 161.665 -131.380 161.835 -129.915 ;
        RECT 162.875 -131.330 163.045 -129.915 ;
        RECT 163.345 -129.960 163.565 -129.760 ;
        RECT 167.435 -129.945 168.550 -129.760 ;
        RECT 161.630 -131.975 161.865 -131.380 ;
        RECT 162.840 -131.975 163.075 -131.330 ;
        RECT 163.365 -131.455 163.535 -129.960 ;
        RECT 157.015 -132.540 164.400 -131.975 ;
        RECT 120.115 -135.695 130.175 -135.685 ;
        RECT 81.445 -135.910 81.615 -135.890 ;
        RECT 71.240 -136.175 74.380 -136.005 ;
        RECT 120.115 -136.535 130.270 -135.695 ;
        RECT 120.115 -136.540 129.890 -136.535 ;
        RECT -40.045 -137.745 -39.230 -137.645 ;
        RECT -98.520 -138.425 -39.230 -137.745 ;
        RECT 44.425 -138.225 45.065 -137.330 ;
        RECT -98.520 -138.430 -97.830 -138.425 ;
        RECT -114.550 -138.655 -113.760 -138.490 ;
        RECT -40.045 -138.520 -39.230 -138.425 ;
        RECT 129.520 -138.505 130.625 -137.530 ;
        RECT 170.995 -137.605 171.725 -110.690 ;
        RECT 175.570 -110.710 176.705 -110.700 ;
        RECT 178.760 -110.710 179.130 -110.580 ;
        RECT 175.570 -110.900 179.130 -110.710 ;
        RECT 179.695 -110.795 182.770 -110.365 ;
        RECT 175.625 -115.150 176.005 -110.900 ;
        RECT 176.700 -110.905 179.130 -110.900 ;
        RECT 176.700 -110.910 177.055 -110.905 ;
        RECT 178.760 -110.935 179.130 -110.905 ;
        RECT 176.860 -112.660 177.030 -111.120 ;
        RECT 177.350 -112.660 177.520 -111.120 ;
        RECT 177.840 -112.660 178.010 -111.120 ;
        RECT 178.330 -112.660 178.500 -111.120 ;
        RECT 178.820 -112.660 178.990 -111.120 ;
        RECT 177.345 -112.920 177.520 -112.660 ;
        RECT 180.915 -112.830 181.220 -110.795 ;
        RECT 183.365 -111.615 183.715 -109.640 ;
        RECT 184.585 -110.910 184.755 -107.990 ;
        RECT 185.620 -108.030 185.830 -107.820 ;
        RECT 184.565 -111.205 184.775 -110.910 ;
        RECT 185.640 -110.940 185.810 -108.030 ;
        RECT 186.130 -110.930 186.300 -107.990 ;
        RECT 186.610 -108.040 186.820 -107.820 ;
        RECT 185.625 -111.205 185.835 -110.940 ;
        RECT 184.565 -111.385 185.835 -111.205 ;
        RECT 186.110 -111.200 186.320 -110.930 ;
        RECT 186.620 -111.030 186.790 -108.040 ;
        RECT 187.680 -110.960 187.850 -107.990 ;
        RECT 186.110 -111.395 186.815 -111.200 ;
        RECT 186.600 -111.455 186.815 -111.395 ;
        RECT 185.390 -111.615 186.165 -111.565 ;
        RECT 183.365 -111.795 186.165 -111.615 ;
        RECT 183.365 -111.805 183.715 -111.795 ;
        RECT 185.390 -111.840 186.165 -111.795 ;
        RECT 186.600 -111.730 187.505 -111.455 ;
        RECT 186.600 -112.080 186.815 -111.730 ;
        RECT 184.040 -112.150 184.815 -112.105 ;
        RECT 183.855 -112.320 184.815 -112.150 ;
        RECT 184.040 -112.380 184.815 -112.320 ;
        RECT 185.045 -112.280 186.815 -112.080 ;
        RECT 187.675 -112.180 187.890 -110.960 ;
        RECT 188.860 -111.305 189.210 -104.620 ;
        RECT 221.795 -105.025 221.965 -103.985 ;
        RECT 222.775 -105.025 222.945 -103.985 ;
        RECT 223.755 -105.025 223.925 -103.985 ;
        RECT 226.660 -105.670 226.830 -103.950 ;
        RECT 227.640 -105.670 227.810 -103.950 ;
        RECT 228.505 -104.695 228.810 -103.950 ;
        RECT 229.705 -104.520 229.875 -103.740 ;
        RECT 230.195 -104.520 230.365 -103.980 ;
        RECT 230.685 -104.520 230.855 -103.740 ;
        RECT 271.735 -103.745 272.410 -103.715 ;
        RECT 272.650 -103.630 274.745 -103.590 ;
        RECT 272.650 -103.780 274.800 -103.630 ;
        RECT 231.175 -104.520 231.345 -103.980 ;
        RECT 229.115 -104.695 229.480 -104.665 ;
        RECT 228.505 -104.760 229.480 -104.695 ;
        RECT 228.615 -104.900 229.480 -104.760 ;
        RECT 229.115 -104.965 229.480 -104.900 ;
        RECT 231.665 -104.815 233.525 -104.465 ;
        RECT 229.705 -105.675 229.875 -105.135 ;
        RECT 230.685 -105.675 230.855 -105.135 ;
        RECT 231.665 -105.675 231.835 -104.815 ;
        RECT 195.440 -107.100 197.045 -106.930 ;
        RECT 194.545 -109.780 194.715 -107.280 ;
        RECT 194.540 -110.010 194.715 -109.780 ;
        RECT 195.440 -110.010 195.640 -107.100 ;
        RECT 195.885 -107.300 196.060 -107.100 ;
        RECT 195.890 -109.820 196.060 -107.300 ;
        RECT 196.380 -109.785 196.550 -107.280 ;
        RECT 196.870 -107.295 197.045 -107.100 ;
        RECT 194.540 -110.210 195.640 -110.010 ;
        RECT 196.365 -110.385 196.555 -109.785 ;
        RECT 196.870 -109.820 197.040 -107.295 ;
        RECT 197.520 -110.200 197.690 -107.280 ;
        RECT 199.150 -109.850 199.320 -107.280 ;
        RECT 200.290 -108.730 200.460 -107.280 ;
        RECT 229.935 -108.015 231.135 -107.845 ;
        RECT 200.285 -109.195 200.470 -108.730 ;
        RECT 200.285 -109.380 200.970 -109.195 ;
        RECT 199.150 -110.020 199.945 -109.850 ;
        RECT 198.265 -110.200 198.955 -110.145 ;
        RECT 194.545 -110.575 196.555 -110.385 ;
        RECT 196.890 -110.370 198.955 -110.200 ;
        RECT 193.360 -110.630 194.050 -110.580 ;
        RECT 191.410 -110.800 194.050 -110.630 ;
        RECT 188.805 -111.665 189.330 -111.305 ;
        RECT 191.410 -112.180 191.625 -110.800 ;
        RECT 193.360 -110.850 194.050 -110.800 ;
        RECT 193.640 -111.305 194.330 -111.260 ;
        RECT 192.590 -111.475 194.330 -111.305 ;
        RECT 192.590 -112.110 192.950 -111.475 ;
        RECT 193.640 -111.530 194.330 -111.475 ;
        RECT 192.590 -112.155 193.010 -112.110 ;
        RECT 178.970 -112.920 181.220 -112.830 ;
        RECT 176.760 -113.135 181.220 -112.920 ;
        RECT 176.760 -113.225 179.005 -113.135 ;
        RECT 172.345 -115.880 176.005 -115.150 ;
        RECT 180.915 -114.610 181.220 -113.135 ;
        RECT 184.585 -114.020 184.755 -112.550 ;
        RECT 185.045 -112.630 185.270 -112.280 ;
        RECT 187.005 -112.380 191.625 -112.180 ;
        RECT 187.245 -112.395 191.625 -112.380 ;
        RECT 184.550 -114.610 184.785 -114.020 ;
        RECT 185.075 -114.090 185.245 -112.630 ;
        RECT 185.565 -114.015 185.735 -112.550 ;
        RECT 186.775 -113.965 186.945 -112.550 ;
        RECT 187.245 -112.595 187.465 -112.395 ;
        RECT 192.615 -112.505 193.010 -112.155 ;
        RECT 185.530 -114.610 185.765 -114.015 ;
        RECT 186.740 -114.610 186.975 -113.965 ;
        RECT 187.265 -114.090 187.435 -112.595 ;
        RECT 194.055 -113.715 194.225 -112.260 ;
        RECT 194.045 -114.270 194.230 -113.715 ;
        RECT 194.545 -113.800 194.715 -110.575 ;
        RECT 195.690 -110.925 195.880 -110.575 ;
        RECT 196.890 -110.765 197.060 -110.370 ;
        RECT 198.265 -110.415 198.955 -110.370 ;
        RECT 195.640 -111.615 195.910 -110.925 ;
        RECT 196.405 -110.935 197.060 -110.765 ;
        RECT 197.390 -110.850 198.080 -110.580 ;
        RECT 199.315 -110.925 199.585 -110.235 ;
        RECT 199.775 -110.240 199.945 -110.020 ;
        RECT 199.775 -110.510 200.605 -110.240 ;
        RECT 196.405 -113.800 196.575 -110.935 ;
        RECT 199.775 -111.085 199.945 -110.510 ;
        RECT 200.205 -111.085 200.475 -111.000 ;
        RECT 196.895 -111.280 197.690 -111.105 ;
        RECT 199.775 -111.110 200.475 -111.085 ;
        RECT 199.635 -111.255 200.475 -111.110 ;
        RECT 196.895 -113.800 197.065 -111.280 ;
        RECT 197.520 -113.800 197.690 -111.280 ;
        RECT 198.010 -113.715 198.180 -111.260 ;
        RECT 198.660 -113.710 198.830 -111.260 ;
        RECT 191.360 -114.290 194.415 -114.270 ;
        RECT 198.005 -114.290 198.190 -113.715 ;
        RECT 198.645 -114.290 198.830 -113.710 ;
        RECT 199.150 -113.800 199.320 -111.260 ;
        RECT 199.635 -111.280 199.945 -111.255 ;
        RECT 199.640 -113.800 199.810 -111.280 ;
        RECT 200.205 -111.295 200.475 -111.255 ;
        RECT 200.780 -111.845 200.970 -109.380 ;
        RECT 221.665 -110.350 221.835 -108.630 ;
        RECT 222.645 -110.350 222.815 -108.630 ;
        RECT 224.710 -109.165 224.880 -108.625 ;
        RECT 225.690 -109.165 225.860 -108.625 ;
        RECT 224.120 -109.400 224.485 -109.335 ;
        RECT 223.620 -109.540 224.485 -109.400 ;
        RECT 223.510 -109.605 224.485 -109.540 ;
        RECT 223.510 -110.350 223.815 -109.605 ;
        RECT 224.120 -109.635 224.485 -109.605 ;
        RECT 226.670 -109.485 226.840 -108.625 ;
        RECT 214.405 -110.425 218.240 -110.390 ;
        RECT 220.750 -110.415 221.425 -110.385 ;
        RECT 220.650 -110.425 221.425 -110.415 ;
        RECT 214.405 -110.605 221.425 -110.425 ;
        RECT 221.665 -110.500 223.815 -110.350 ;
        RECT 221.665 -110.540 223.760 -110.500 ;
        RECT 224.710 -110.560 224.880 -109.780 ;
        RECT 225.200 -110.320 225.370 -109.780 ;
        RECT 225.690 -110.560 225.860 -109.780 ;
        RECT 226.180 -110.320 226.350 -109.780 ;
        RECT 226.670 -109.835 228.060 -109.485 ;
        RECT 214.405 -111.120 218.240 -110.605 ;
        RECT 220.650 -110.615 221.425 -110.605 ;
        RECT 220.750 -110.655 221.425 -110.615 ;
        RECT 219.885 -110.905 221.020 -110.895 ;
        RECT 223.075 -110.905 223.445 -110.775 ;
        RECT 219.885 -111.095 223.445 -110.905 ;
        RECT 224.010 -110.990 227.085 -110.560 ;
        RECT 200.780 -112.035 202.240 -111.845 ;
        RECT 200.290 -113.705 200.460 -112.260 ;
        RECT 200.780 -112.285 200.970 -112.035 ;
        RECT 200.280 -114.290 200.465 -113.705 ;
        RECT 200.780 -113.800 200.950 -112.285 ;
        RECT 191.360 -114.610 201.030 -114.290 ;
        RECT 180.915 -114.835 201.030 -114.610 ;
        RECT 180.915 -115.175 191.925 -114.835 ;
        RECT 193.665 -115.095 201.030 -114.835 ;
        RECT 172.345 -135.795 173.075 -115.880 ;
        RECT 175.625 -116.540 176.005 -115.880 ;
        RECT 202.050 -116.510 202.240 -112.035 ;
        RECT 175.625 -116.920 192.175 -116.540 ;
        RECT 175.625 -117.830 176.005 -116.920 ;
        RECT 175.625 -118.210 176.335 -117.830 ;
        RECT 175.955 -120.155 176.335 -118.210 ;
        RECT 181.000 -118.040 184.325 -117.900 ;
        RECT 181.000 -118.330 186.175 -118.040 ;
        RECT 190.045 -118.325 190.505 -117.900 ;
        RECT 181.000 -118.735 181.430 -118.330 ;
        RECT 182.300 -118.515 182.475 -118.330 ;
        RECT 183.925 -118.345 186.175 -118.330 ;
        RECT 176.740 -119.165 181.430 -118.735 ;
        RECT 175.955 -120.615 176.630 -120.155 ;
        RECT 177.440 -120.445 177.610 -119.165 ;
        RECT 177.930 -120.445 178.100 -119.405 ;
        RECT 178.420 -120.445 178.590 -119.165 ;
        RECT 178.910 -120.275 179.080 -119.405 ;
        RECT 181.815 -120.055 181.985 -118.515 ;
        RECT 182.305 -120.055 182.475 -118.515 ;
        RECT 182.795 -120.055 182.965 -118.515 ;
        RECT 183.285 -120.055 183.455 -118.515 ;
        RECT 183.775 -120.055 183.945 -118.515 ;
        RECT 181.655 -120.270 182.010 -120.265 ;
        RECT 183.715 -120.270 184.085 -120.240 ;
        RECT 181.655 -120.275 184.085 -120.270 ;
        RECT 178.910 -120.445 184.085 -120.275 ;
        RECT 185.870 -120.380 186.175 -118.345 ;
        RECT 178.915 -120.465 184.085 -120.445 ;
        RECT 178.915 -120.475 181.660 -120.465 ;
        RECT 176.850 -120.615 177.215 -120.585 ;
        RECT 183.715 -120.595 184.085 -120.465 ;
        RECT 175.955 -120.700 177.215 -120.615 ;
        RECT 175.980 -120.820 177.215 -120.700 ;
        RECT 181.390 -120.755 182.065 -120.715 ;
        RECT 181.290 -120.765 182.065 -120.755 ;
        RECT 175.980 -120.905 176.630 -120.820 ;
        RECT 176.850 -120.885 177.215 -120.820 ;
        RECT 180.255 -120.945 182.065 -120.765 ;
        RECT 184.650 -120.810 188.575 -120.380 ;
        RECT 181.290 -120.955 182.065 -120.945 ;
        RECT 181.390 -120.985 182.065 -120.955 ;
        RECT 182.305 -120.870 184.400 -120.830 ;
        RECT 182.305 -121.020 184.455 -120.870 ;
        RECT 177.440 -122.095 177.610 -121.055 ;
        RECT 178.420 -122.095 178.590 -121.055 ;
        RECT 179.400 -122.095 179.570 -121.055 ;
        RECT 182.305 -122.740 182.475 -121.020 ;
        RECT 183.285 -122.740 183.455 -121.020 ;
        RECT 184.150 -121.765 184.455 -121.020 ;
        RECT 185.350 -121.590 185.520 -120.810 ;
        RECT 185.840 -121.590 186.010 -121.050 ;
        RECT 186.330 -121.590 186.500 -120.810 ;
        RECT 186.820 -121.590 186.990 -121.050 ;
        RECT 184.760 -121.765 185.125 -121.735 ;
        RECT 184.150 -121.830 185.125 -121.765 ;
        RECT 184.260 -121.970 185.125 -121.830 ;
        RECT 184.760 -122.035 185.125 -121.970 ;
        RECT 187.310 -121.885 189.170 -121.535 ;
        RECT 185.350 -122.745 185.520 -122.205 ;
        RECT 186.330 -122.745 186.500 -122.205 ;
        RECT 187.310 -122.745 187.480 -121.885 ;
        RECT 185.580 -125.085 186.780 -124.915 ;
        RECT 177.310 -127.420 177.480 -125.700 ;
        RECT 178.290 -127.420 178.460 -125.700 ;
        RECT 180.355 -126.235 180.525 -125.695 ;
        RECT 181.335 -126.235 181.505 -125.695 ;
        RECT 179.765 -126.470 180.130 -126.405 ;
        RECT 179.265 -126.610 180.130 -126.470 ;
        RECT 179.155 -126.675 180.130 -126.610 ;
        RECT 179.155 -127.420 179.460 -126.675 ;
        RECT 179.765 -126.705 180.130 -126.675 ;
        RECT 182.315 -126.555 182.485 -125.695 ;
        RECT 177.310 -127.570 179.460 -127.420 ;
        RECT 177.310 -127.610 179.405 -127.570 ;
        RECT 180.355 -127.630 180.525 -126.850 ;
        RECT 180.845 -127.390 181.015 -126.850 ;
        RECT 181.335 -127.630 181.505 -126.850 ;
        RECT 181.825 -127.390 181.995 -126.850 ;
        RECT 182.315 -126.905 183.705 -126.555 ;
        RECT 175.530 -127.975 176.665 -127.965 ;
        RECT 178.720 -127.975 179.090 -127.845 ;
        RECT 175.530 -128.165 179.090 -127.975 ;
        RECT 179.655 -128.060 182.730 -127.630 ;
        RECT 176.660 -128.170 179.090 -128.165 ;
        RECT 176.660 -128.175 177.015 -128.170 ;
        RECT 178.720 -128.200 179.090 -128.170 ;
        RECT 176.820 -129.925 176.990 -128.385 ;
        RECT 177.310 -129.925 177.480 -128.385 ;
        RECT 177.800 -129.925 177.970 -128.385 ;
        RECT 178.290 -129.925 178.460 -128.385 ;
        RECT 178.780 -129.925 178.950 -128.385 ;
        RECT 177.305 -130.185 177.480 -129.925 ;
        RECT 180.875 -130.095 181.180 -128.060 ;
        RECT 183.325 -128.880 183.675 -126.905 ;
        RECT 184.545 -128.175 184.715 -125.255 ;
        RECT 185.580 -125.295 185.790 -125.085 ;
        RECT 184.525 -128.470 184.735 -128.175 ;
        RECT 185.600 -128.205 185.770 -125.295 ;
        RECT 186.090 -128.195 186.260 -125.255 ;
        RECT 186.570 -125.305 186.780 -125.085 ;
        RECT 185.585 -128.470 185.795 -128.205 ;
        RECT 184.525 -128.650 185.795 -128.470 ;
        RECT 186.070 -128.465 186.280 -128.195 ;
        RECT 186.580 -128.295 186.750 -125.305 ;
        RECT 187.640 -128.225 187.810 -125.255 ;
        RECT 186.070 -128.660 186.775 -128.465 ;
        RECT 186.560 -128.720 186.775 -128.660 ;
        RECT 185.350 -128.880 186.125 -128.830 ;
        RECT 183.325 -129.060 186.125 -128.880 ;
        RECT 183.325 -129.070 183.675 -129.060 ;
        RECT 185.350 -129.105 186.125 -129.060 ;
        RECT 186.560 -128.995 187.465 -128.720 ;
        RECT 186.560 -129.345 186.775 -128.995 ;
        RECT 184.000 -129.415 184.775 -129.370 ;
        RECT 183.815 -129.585 184.775 -129.415 ;
        RECT 184.000 -129.645 184.775 -129.585 ;
        RECT 185.005 -129.545 186.775 -129.345 ;
        RECT 187.635 -129.445 187.850 -128.225 ;
        RECT 188.820 -128.570 189.170 -121.885 ;
        RECT 190.160 -128.200 190.375 -118.325 ;
        RECT 191.795 -120.440 192.175 -116.920 ;
        RECT 193.305 -116.700 202.240 -116.510 ;
        RECT 193.305 -118.590 193.495 -116.700 ;
        RECT 199.340 -118.195 202.665 -118.055 ;
        RECT 199.340 -118.485 204.515 -118.195 ;
        RECT 193.190 -118.860 193.555 -118.590 ;
        RECT 199.340 -118.890 199.770 -118.485 ;
        RECT 200.640 -118.670 200.815 -118.485 ;
        RECT 202.265 -118.500 204.515 -118.485 ;
        RECT 195.080 -119.320 199.770 -118.890 ;
        RECT 194.320 -120.440 194.970 -120.310 ;
        RECT 191.795 -120.770 194.970 -120.440 ;
        RECT 195.780 -120.600 195.950 -119.320 ;
        RECT 196.270 -120.600 196.440 -119.560 ;
        RECT 196.760 -120.600 196.930 -119.320 ;
        RECT 197.250 -120.430 197.420 -119.560 ;
        RECT 200.155 -120.210 200.325 -118.670 ;
        RECT 200.645 -120.210 200.815 -118.670 ;
        RECT 201.135 -120.210 201.305 -118.670 ;
        RECT 201.625 -120.210 201.795 -118.670 ;
        RECT 202.115 -120.210 202.285 -118.670 ;
        RECT 199.995 -120.425 200.350 -120.420 ;
        RECT 202.055 -120.425 202.425 -120.395 ;
        RECT 199.995 -120.430 202.425 -120.425 ;
        RECT 197.250 -120.600 202.425 -120.430 ;
        RECT 204.210 -120.535 204.515 -118.500 ;
        RECT 197.255 -120.620 202.425 -120.600 ;
        RECT 197.255 -120.630 200.000 -120.620 ;
        RECT 195.190 -120.770 195.555 -120.740 ;
        RECT 202.055 -120.750 202.425 -120.620 ;
        RECT 191.795 -120.820 195.555 -120.770 ;
        RECT 194.320 -120.975 195.555 -120.820 ;
        RECT 199.730 -120.910 200.405 -120.870 ;
        RECT 199.630 -120.920 200.405 -120.910 ;
        RECT 194.320 -121.060 194.970 -120.975 ;
        RECT 195.190 -121.040 195.555 -120.975 ;
        RECT 194.455 -121.310 194.835 -121.060 ;
        RECT 198.595 -121.100 200.405 -120.920 ;
        RECT 202.990 -120.965 206.915 -120.535 ;
        RECT 199.630 -121.110 200.405 -121.100 ;
        RECT 199.730 -121.140 200.405 -121.110 ;
        RECT 200.645 -121.025 202.740 -120.985 ;
        RECT 200.645 -121.175 202.795 -121.025 ;
        RECT 195.780 -122.250 195.950 -121.210 ;
        RECT 196.760 -122.250 196.930 -121.210 ;
        RECT 197.740 -122.250 197.910 -121.210 ;
        RECT 200.645 -122.895 200.815 -121.175 ;
        RECT 201.625 -122.895 201.795 -121.175 ;
        RECT 202.490 -121.920 202.795 -121.175 ;
        RECT 203.690 -121.745 203.860 -120.965 ;
        RECT 204.180 -121.745 204.350 -121.205 ;
        RECT 204.670 -121.745 204.840 -120.965 ;
        RECT 205.160 -121.745 205.330 -121.205 ;
        RECT 203.100 -121.920 203.465 -121.890 ;
        RECT 202.490 -121.985 203.465 -121.920 ;
        RECT 202.600 -122.125 203.465 -121.985 ;
        RECT 203.100 -122.190 203.465 -122.125 ;
        RECT 205.650 -122.040 207.510 -121.690 ;
        RECT 203.690 -122.900 203.860 -122.360 ;
        RECT 204.670 -122.900 204.840 -122.360 ;
        RECT 205.650 -122.900 205.820 -122.040 ;
        RECT 203.920 -125.240 205.120 -125.070 ;
        RECT 195.650 -127.575 195.820 -125.855 ;
        RECT 196.630 -127.575 196.800 -125.855 ;
        RECT 198.695 -126.390 198.865 -125.850 ;
        RECT 199.675 -126.390 199.845 -125.850 ;
        RECT 198.105 -126.625 198.470 -126.560 ;
        RECT 197.605 -126.765 198.470 -126.625 ;
        RECT 197.495 -126.830 198.470 -126.765 ;
        RECT 197.495 -127.575 197.800 -126.830 ;
        RECT 198.105 -126.860 198.470 -126.830 ;
        RECT 200.655 -126.710 200.825 -125.850 ;
        RECT 195.650 -127.725 197.800 -127.575 ;
        RECT 195.650 -127.765 197.745 -127.725 ;
        RECT 198.695 -127.785 198.865 -127.005 ;
        RECT 199.185 -127.545 199.355 -127.005 ;
        RECT 199.675 -127.785 199.845 -127.005 ;
        RECT 200.165 -127.545 200.335 -127.005 ;
        RECT 200.655 -127.060 202.045 -126.710 ;
        RECT 193.870 -128.130 195.005 -128.120 ;
        RECT 197.060 -128.130 197.430 -128.000 ;
        RECT 190.160 -128.415 191.585 -128.200 ;
        RECT 193.870 -128.320 197.430 -128.130 ;
        RECT 197.995 -128.215 201.070 -127.785 ;
        RECT 195.000 -128.325 197.430 -128.320 ;
        RECT 195.000 -128.330 195.355 -128.325 ;
        RECT 197.060 -128.355 197.430 -128.325 ;
        RECT 188.765 -128.930 189.290 -128.570 ;
        RECT 191.370 -129.445 191.585 -128.415 ;
        RECT 178.930 -130.185 181.180 -130.095 ;
        RECT 176.720 -130.400 181.180 -130.185 ;
        RECT 176.720 -130.490 178.965 -130.400 ;
        RECT 180.875 -131.875 181.180 -130.400 ;
        RECT 184.545 -131.285 184.715 -129.815 ;
        RECT 185.005 -129.895 185.230 -129.545 ;
        RECT 186.965 -129.645 191.585 -129.445 ;
        RECT 187.205 -129.660 191.585 -129.645 ;
        RECT 184.510 -131.875 184.745 -131.285 ;
        RECT 185.035 -131.355 185.205 -129.895 ;
        RECT 185.525 -131.280 185.695 -129.815 ;
        RECT 186.735 -131.230 186.905 -129.815 ;
        RECT 187.205 -129.860 187.425 -129.660 ;
        RECT 185.490 -131.875 185.725 -131.280 ;
        RECT 186.700 -131.875 186.935 -131.230 ;
        RECT 187.225 -131.355 187.395 -129.860 ;
        RECT 195.160 -130.080 195.330 -128.540 ;
        RECT 195.650 -130.080 195.820 -128.540 ;
        RECT 196.140 -130.080 196.310 -128.540 ;
        RECT 196.630 -130.080 196.800 -128.540 ;
        RECT 197.120 -130.080 197.290 -128.540 ;
        RECT 195.645 -130.340 195.820 -130.080 ;
        RECT 199.215 -130.250 199.520 -128.215 ;
        RECT 201.665 -129.035 202.015 -127.060 ;
        RECT 202.885 -128.330 203.055 -125.410 ;
        RECT 203.920 -125.450 204.130 -125.240 ;
        RECT 202.865 -128.625 203.075 -128.330 ;
        RECT 203.940 -128.360 204.110 -125.450 ;
        RECT 204.430 -128.350 204.600 -125.410 ;
        RECT 204.910 -125.460 205.120 -125.240 ;
        RECT 203.925 -128.625 204.135 -128.360 ;
        RECT 202.865 -128.805 204.135 -128.625 ;
        RECT 204.410 -128.620 204.620 -128.350 ;
        RECT 204.920 -128.450 205.090 -125.460 ;
        RECT 205.980 -128.380 206.150 -125.410 ;
        RECT 204.410 -128.815 205.115 -128.620 ;
        RECT 204.900 -128.875 205.115 -128.815 ;
        RECT 203.690 -129.035 204.465 -128.985 ;
        RECT 201.665 -129.215 204.465 -129.035 ;
        RECT 201.665 -129.225 202.015 -129.215 ;
        RECT 203.690 -129.260 204.465 -129.215 ;
        RECT 204.900 -129.150 205.805 -128.875 ;
        RECT 204.900 -129.500 205.115 -129.150 ;
        RECT 202.340 -129.570 203.115 -129.525 ;
        RECT 202.155 -129.740 203.115 -129.570 ;
        RECT 202.340 -129.800 203.115 -129.740 ;
        RECT 203.345 -129.700 205.115 -129.500 ;
        RECT 205.975 -129.600 206.190 -128.380 ;
        RECT 207.160 -128.725 207.510 -122.040 ;
        RECT 207.105 -129.085 207.630 -128.725 ;
        RECT 209.680 -129.600 211.365 -128.785 ;
        RECT 197.270 -130.340 199.520 -130.250 ;
        RECT 195.060 -130.555 199.520 -130.340 ;
        RECT 195.060 -130.645 197.305 -130.555 ;
        RECT 180.875 -132.440 188.260 -131.875 ;
        RECT 199.215 -132.030 199.520 -130.555 ;
        RECT 202.885 -131.440 203.055 -129.970 ;
        RECT 203.345 -130.050 203.570 -129.700 ;
        RECT 205.305 -129.800 211.365 -129.600 ;
        RECT 205.545 -129.815 211.365 -129.800 ;
        RECT 202.850 -132.030 203.085 -131.440 ;
        RECT 203.375 -131.510 203.545 -130.050 ;
        RECT 203.865 -131.435 204.035 -129.970 ;
        RECT 205.075 -131.385 205.245 -129.970 ;
        RECT 205.545 -130.015 205.765 -129.815 ;
        RECT 203.830 -132.030 204.065 -131.435 ;
        RECT 205.040 -132.030 205.275 -131.385 ;
        RECT 205.565 -131.510 205.735 -130.015 ;
        RECT 209.680 -130.440 211.365 -129.815 ;
        RECT 199.215 -132.595 206.600 -132.030 ;
        RECT 172.230 -136.530 173.245 -135.795 ;
        RECT 207.885 -136.700 209.470 -135.245 ;
        RECT 170.650 -138.620 172.020 -137.605 ;
        RECT -99.210 -138.655 -98.525 -138.630 ;
        RECT -114.550 -138.915 -98.525 -138.655 ;
        RECT -114.550 -139.070 -113.760 -138.915 ;
        RECT -99.210 -138.920 -98.525 -138.915 ;
        RECT 207.970 -140.600 209.300 -136.700 ;
        RECT 214.405 -137.695 215.135 -111.120 ;
        RECT 219.940 -115.785 220.320 -111.095 ;
        RECT 221.015 -111.100 223.445 -111.095 ;
        RECT 221.015 -111.105 221.370 -111.100 ;
        RECT 223.075 -111.130 223.445 -111.100 ;
        RECT 221.175 -112.855 221.345 -111.315 ;
        RECT 221.665 -112.855 221.835 -111.315 ;
        RECT 222.155 -112.855 222.325 -111.315 ;
        RECT 222.645 -112.855 222.815 -111.315 ;
        RECT 223.135 -112.855 223.305 -111.315 ;
        RECT 221.660 -113.115 221.835 -112.855 ;
        RECT 225.230 -113.025 225.535 -110.990 ;
        RECT 227.680 -111.810 228.030 -109.835 ;
        RECT 228.900 -111.105 229.070 -108.185 ;
        RECT 229.935 -108.225 230.145 -108.015 ;
        RECT 228.880 -111.400 229.090 -111.105 ;
        RECT 229.955 -111.135 230.125 -108.225 ;
        RECT 230.445 -111.125 230.615 -108.185 ;
        RECT 230.925 -108.235 231.135 -108.015 ;
        RECT 229.940 -111.400 230.150 -111.135 ;
        RECT 228.880 -111.580 230.150 -111.400 ;
        RECT 230.425 -111.395 230.635 -111.125 ;
        RECT 230.935 -111.225 231.105 -108.235 ;
        RECT 231.995 -111.155 232.165 -108.185 ;
        RECT 230.425 -111.590 231.130 -111.395 ;
        RECT 230.915 -111.650 231.130 -111.590 ;
        RECT 229.705 -111.810 230.480 -111.760 ;
        RECT 227.680 -111.990 230.480 -111.810 ;
        RECT 227.680 -112.000 228.030 -111.990 ;
        RECT 229.705 -112.035 230.480 -111.990 ;
        RECT 230.915 -111.925 231.820 -111.650 ;
        RECT 230.915 -112.275 231.130 -111.925 ;
        RECT 228.355 -112.345 229.130 -112.300 ;
        RECT 228.170 -112.515 229.130 -112.345 ;
        RECT 228.355 -112.575 229.130 -112.515 ;
        RECT 229.360 -112.475 231.130 -112.275 ;
        RECT 231.990 -112.375 232.205 -111.155 ;
        RECT 233.175 -111.500 233.525 -104.815 ;
        RECT 267.785 -104.855 267.955 -103.815 ;
        RECT 268.765 -104.855 268.935 -103.815 ;
        RECT 269.745 -104.855 269.915 -103.815 ;
        RECT 272.650 -105.500 272.820 -103.780 ;
        RECT 273.630 -105.500 273.800 -103.780 ;
        RECT 274.495 -104.525 274.800 -103.780 ;
        RECT 275.695 -104.350 275.865 -103.570 ;
        RECT 276.185 -104.350 276.355 -103.810 ;
        RECT 276.675 -104.350 276.845 -103.570 ;
        RECT 277.165 -104.350 277.335 -103.810 ;
        RECT 275.105 -104.525 275.470 -104.495 ;
        RECT 274.495 -104.590 275.470 -104.525 ;
        RECT 274.605 -104.730 275.470 -104.590 ;
        RECT 275.105 -104.795 275.470 -104.730 ;
        RECT 277.655 -104.645 279.515 -104.295 ;
        RECT 311.555 -104.525 311.725 -103.485 ;
        RECT 312.535 -104.525 312.705 -103.485 ;
        RECT 313.515 -104.525 313.685 -103.485 ;
        RECT 275.695 -105.505 275.865 -104.965 ;
        RECT 276.675 -105.505 276.845 -104.965 ;
        RECT 277.655 -105.505 277.825 -104.645 ;
        RECT 239.755 -107.295 241.360 -107.125 ;
        RECT 238.860 -109.975 239.030 -107.475 ;
        RECT 238.855 -110.205 239.030 -109.975 ;
        RECT 239.755 -110.205 239.955 -107.295 ;
        RECT 240.200 -107.495 240.375 -107.295 ;
        RECT 240.205 -110.015 240.375 -107.495 ;
        RECT 240.695 -109.980 240.865 -107.475 ;
        RECT 241.185 -107.490 241.360 -107.295 ;
        RECT 238.855 -110.405 239.955 -110.205 ;
        RECT 240.680 -110.580 240.870 -109.980 ;
        RECT 241.185 -110.015 241.355 -107.490 ;
        RECT 241.835 -110.395 242.005 -107.475 ;
        RECT 243.465 -110.045 243.635 -107.475 ;
        RECT 244.605 -108.925 244.775 -107.475 ;
        RECT 275.925 -107.845 277.125 -107.675 ;
        RECT 244.600 -109.390 244.785 -108.925 ;
        RECT 244.600 -109.575 245.285 -109.390 ;
        RECT 243.465 -110.215 244.260 -110.045 ;
        RECT 242.580 -110.395 243.270 -110.340 ;
        RECT 238.860 -110.770 240.870 -110.580 ;
        RECT 241.205 -110.565 243.270 -110.395 ;
        RECT 237.675 -110.825 238.365 -110.775 ;
        RECT 235.725 -110.995 238.365 -110.825 ;
        RECT 233.120 -111.860 233.645 -111.500 ;
        RECT 235.725 -112.375 235.940 -110.995 ;
        RECT 237.675 -111.045 238.365 -110.995 ;
        RECT 237.955 -111.500 238.645 -111.455 ;
        RECT 236.905 -111.670 238.645 -111.500 ;
        RECT 236.905 -112.305 237.265 -111.670 ;
        RECT 237.955 -111.725 238.645 -111.670 ;
        RECT 236.905 -112.350 237.325 -112.305 ;
        RECT 223.285 -113.115 225.535 -113.025 ;
        RECT 221.075 -113.330 225.535 -113.115 ;
        RECT 221.075 -113.420 223.320 -113.330 ;
        RECT 225.230 -114.805 225.535 -113.330 ;
        RECT 228.900 -114.215 229.070 -112.745 ;
        RECT 229.360 -112.825 229.585 -112.475 ;
        RECT 231.320 -112.575 235.940 -112.375 ;
        RECT 231.560 -112.590 235.940 -112.575 ;
        RECT 228.865 -114.805 229.100 -114.215 ;
        RECT 229.390 -114.285 229.560 -112.825 ;
        RECT 229.880 -114.210 230.050 -112.745 ;
        RECT 231.090 -114.160 231.260 -112.745 ;
        RECT 231.560 -112.790 231.780 -112.590 ;
        RECT 236.930 -112.700 237.325 -112.350 ;
        RECT 229.845 -114.805 230.080 -114.210 ;
        RECT 231.055 -114.805 231.290 -114.160 ;
        RECT 231.580 -114.285 231.750 -112.790 ;
        RECT 238.370 -113.910 238.540 -112.455 ;
        RECT 238.360 -114.465 238.545 -113.910 ;
        RECT 238.860 -113.995 239.030 -110.770 ;
        RECT 240.005 -111.120 240.195 -110.770 ;
        RECT 241.205 -110.960 241.375 -110.565 ;
        RECT 242.580 -110.610 243.270 -110.565 ;
        RECT 239.955 -111.810 240.225 -111.120 ;
        RECT 240.720 -111.130 241.375 -110.960 ;
        RECT 241.705 -111.045 242.395 -110.775 ;
        RECT 243.630 -111.120 243.900 -110.430 ;
        RECT 244.090 -110.435 244.260 -110.215 ;
        RECT 244.090 -110.705 244.920 -110.435 ;
        RECT 240.720 -113.995 240.890 -111.130 ;
        RECT 244.090 -111.280 244.260 -110.705 ;
        RECT 244.520 -111.280 244.790 -111.195 ;
        RECT 241.210 -111.475 242.005 -111.300 ;
        RECT 244.090 -111.305 244.790 -111.280 ;
        RECT 243.950 -111.450 244.790 -111.305 ;
        RECT 241.210 -113.995 241.380 -111.475 ;
        RECT 241.835 -113.995 242.005 -111.475 ;
        RECT 242.325 -113.910 242.495 -111.455 ;
        RECT 242.975 -113.905 243.145 -111.455 ;
        RECT 235.675 -114.485 238.730 -114.465 ;
        RECT 242.320 -114.485 242.505 -113.910 ;
        RECT 242.960 -114.485 243.145 -113.905 ;
        RECT 243.465 -113.995 243.635 -111.455 ;
        RECT 243.950 -111.475 244.260 -111.450 ;
        RECT 243.955 -113.995 244.125 -111.475 ;
        RECT 244.520 -111.490 244.790 -111.450 ;
        RECT 245.095 -112.040 245.285 -109.575 ;
        RECT 261.000 -110.255 264.645 -109.930 ;
        RECT 267.655 -110.180 267.825 -108.460 ;
        RECT 268.635 -110.180 268.805 -108.460 ;
        RECT 270.700 -108.995 270.870 -108.455 ;
        RECT 271.680 -108.995 271.850 -108.455 ;
        RECT 270.110 -109.230 270.475 -109.165 ;
        RECT 269.610 -109.370 270.475 -109.230 ;
        RECT 269.500 -109.435 270.475 -109.370 ;
        RECT 269.500 -110.180 269.805 -109.435 ;
        RECT 270.110 -109.465 270.475 -109.435 ;
        RECT 272.660 -109.315 272.830 -108.455 ;
        RECT 266.740 -110.245 267.415 -110.215 ;
        RECT 266.640 -110.255 267.415 -110.245 ;
        RECT 261.000 -110.435 267.415 -110.255 ;
        RECT 267.655 -110.330 269.805 -110.180 ;
        RECT 267.655 -110.370 269.750 -110.330 ;
        RECT 270.700 -110.390 270.870 -109.610 ;
        RECT 271.190 -110.150 271.360 -109.610 ;
        RECT 271.680 -110.390 271.850 -109.610 ;
        RECT 272.170 -110.150 272.340 -109.610 ;
        RECT 272.660 -109.665 274.050 -109.315 ;
        RECT 261.000 -110.660 264.645 -110.435 ;
        RECT 266.640 -110.445 267.415 -110.435 ;
        RECT 266.740 -110.485 267.415 -110.445 ;
        RECT 245.095 -112.230 246.555 -112.040 ;
        RECT 244.605 -113.900 244.775 -112.455 ;
        RECT 245.095 -112.480 245.285 -112.230 ;
        RECT 244.595 -114.485 244.780 -113.900 ;
        RECT 245.095 -113.995 245.265 -112.480 ;
        RECT 235.675 -114.805 245.345 -114.485 ;
        RECT 225.230 -115.030 245.345 -114.805 ;
        RECT 225.230 -115.370 236.240 -115.030 ;
        RECT 237.980 -115.290 245.345 -115.030 ;
        RECT 216.690 -116.515 220.320 -115.785 ;
        RECT 216.690 -136.520 217.420 -116.515 ;
        RECT 219.940 -116.735 220.320 -116.515 ;
        RECT 246.365 -116.705 246.555 -112.230 ;
        RECT 219.940 -117.115 236.490 -116.735 ;
        RECT 219.940 -118.025 220.320 -117.115 ;
        RECT 219.940 -118.405 220.650 -118.025 ;
        RECT 220.270 -120.350 220.650 -118.405 ;
        RECT 225.315 -118.235 228.640 -118.095 ;
        RECT 225.315 -118.525 230.490 -118.235 ;
        RECT 234.360 -118.520 234.820 -118.095 ;
        RECT 225.315 -118.930 225.745 -118.525 ;
        RECT 226.615 -118.710 226.790 -118.525 ;
        RECT 228.240 -118.540 230.490 -118.525 ;
        RECT 221.055 -119.360 225.745 -118.930 ;
        RECT 220.270 -120.810 220.945 -120.350 ;
        RECT 221.755 -120.640 221.925 -119.360 ;
        RECT 222.245 -120.640 222.415 -119.600 ;
        RECT 222.735 -120.640 222.905 -119.360 ;
        RECT 223.225 -120.470 223.395 -119.600 ;
        RECT 226.130 -120.250 226.300 -118.710 ;
        RECT 226.620 -120.250 226.790 -118.710 ;
        RECT 227.110 -120.250 227.280 -118.710 ;
        RECT 227.600 -120.250 227.770 -118.710 ;
        RECT 228.090 -120.250 228.260 -118.710 ;
        RECT 225.970 -120.465 226.325 -120.460 ;
        RECT 228.030 -120.465 228.400 -120.435 ;
        RECT 225.970 -120.470 228.400 -120.465 ;
        RECT 223.225 -120.640 228.400 -120.470 ;
        RECT 230.185 -120.575 230.490 -118.540 ;
        RECT 223.230 -120.660 228.400 -120.640 ;
        RECT 223.230 -120.670 225.975 -120.660 ;
        RECT 221.165 -120.810 221.530 -120.780 ;
        RECT 228.030 -120.790 228.400 -120.660 ;
        RECT 220.270 -120.895 221.530 -120.810 ;
        RECT 220.295 -121.015 221.530 -120.895 ;
        RECT 225.705 -120.950 226.380 -120.910 ;
        RECT 225.605 -120.960 226.380 -120.950 ;
        RECT 220.295 -121.100 220.945 -121.015 ;
        RECT 221.165 -121.080 221.530 -121.015 ;
        RECT 224.570 -121.140 226.380 -120.960 ;
        RECT 228.965 -121.005 232.890 -120.575 ;
        RECT 225.605 -121.150 226.380 -121.140 ;
        RECT 225.705 -121.180 226.380 -121.150 ;
        RECT 226.620 -121.065 228.715 -121.025 ;
        RECT 226.620 -121.215 228.770 -121.065 ;
        RECT 221.755 -122.290 221.925 -121.250 ;
        RECT 222.735 -122.290 222.905 -121.250 ;
        RECT 223.715 -122.290 223.885 -121.250 ;
        RECT 226.620 -122.935 226.790 -121.215 ;
        RECT 227.600 -122.935 227.770 -121.215 ;
        RECT 228.465 -121.960 228.770 -121.215 ;
        RECT 229.665 -121.785 229.835 -121.005 ;
        RECT 230.155 -121.785 230.325 -121.245 ;
        RECT 230.645 -121.785 230.815 -121.005 ;
        RECT 231.135 -121.785 231.305 -121.245 ;
        RECT 229.075 -121.960 229.440 -121.930 ;
        RECT 228.465 -122.025 229.440 -121.960 ;
        RECT 228.575 -122.165 229.440 -122.025 ;
        RECT 229.075 -122.230 229.440 -122.165 ;
        RECT 231.625 -122.080 233.485 -121.730 ;
        RECT 229.665 -122.940 229.835 -122.400 ;
        RECT 230.645 -122.940 230.815 -122.400 ;
        RECT 231.625 -122.940 231.795 -122.080 ;
        RECT 229.895 -125.280 231.095 -125.110 ;
        RECT 221.625 -127.615 221.795 -125.895 ;
        RECT 222.605 -127.615 222.775 -125.895 ;
        RECT 224.670 -126.430 224.840 -125.890 ;
        RECT 225.650 -126.430 225.820 -125.890 ;
        RECT 224.080 -126.665 224.445 -126.600 ;
        RECT 223.580 -126.805 224.445 -126.665 ;
        RECT 223.470 -126.870 224.445 -126.805 ;
        RECT 223.470 -127.615 223.775 -126.870 ;
        RECT 224.080 -126.900 224.445 -126.870 ;
        RECT 226.630 -126.750 226.800 -125.890 ;
        RECT 221.625 -127.765 223.775 -127.615 ;
        RECT 221.625 -127.805 223.720 -127.765 ;
        RECT 224.670 -127.825 224.840 -127.045 ;
        RECT 225.160 -127.585 225.330 -127.045 ;
        RECT 225.650 -127.825 225.820 -127.045 ;
        RECT 226.140 -127.585 226.310 -127.045 ;
        RECT 226.630 -127.100 228.020 -126.750 ;
        RECT 219.845 -128.170 220.980 -128.160 ;
        RECT 223.035 -128.170 223.405 -128.040 ;
        RECT 219.845 -128.360 223.405 -128.170 ;
        RECT 223.970 -128.255 227.045 -127.825 ;
        RECT 220.975 -128.365 223.405 -128.360 ;
        RECT 220.975 -128.370 221.330 -128.365 ;
        RECT 223.035 -128.395 223.405 -128.365 ;
        RECT 221.135 -130.120 221.305 -128.580 ;
        RECT 221.625 -130.120 221.795 -128.580 ;
        RECT 222.115 -130.120 222.285 -128.580 ;
        RECT 222.605 -130.120 222.775 -128.580 ;
        RECT 223.095 -130.120 223.265 -128.580 ;
        RECT 221.620 -130.380 221.795 -130.120 ;
        RECT 225.190 -130.290 225.495 -128.255 ;
        RECT 227.640 -129.075 227.990 -127.100 ;
        RECT 228.860 -128.370 229.030 -125.450 ;
        RECT 229.895 -125.490 230.105 -125.280 ;
        RECT 228.840 -128.665 229.050 -128.370 ;
        RECT 229.915 -128.400 230.085 -125.490 ;
        RECT 230.405 -128.390 230.575 -125.450 ;
        RECT 230.885 -125.500 231.095 -125.280 ;
        RECT 229.900 -128.665 230.110 -128.400 ;
        RECT 228.840 -128.845 230.110 -128.665 ;
        RECT 230.385 -128.660 230.595 -128.390 ;
        RECT 230.895 -128.490 231.065 -125.500 ;
        RECT 231.955 -128.420 232.125 -125.450 ;
        RECT 230.385 -128.855 231.090 -128.660 ;
        RECT 230.875 -128.915 231.090 -128.855 ;
        RECT 229.665 -129.075 230.440 -129.025 ;
        RECT 227.640 -129.255 230.440 -129.075 ;
        RECT 227.640 -129.265 227.990 -129.255 ;
        RECT 229.665 -129.300 230.440 -129.255 ;
        RECT 230.875 -129.190 231.780 -128.915 ;
        RECT 230.875 -129.540 231.090 -129.190 ;
        RECT 228.315 -129.610 229.090 -129.565 ;
        RECT 228.130 -129.780 229.090 -129.610 ;
        RECT 228.315 -129.840 229.090 -129.780 ;
        RECT 229.320 -129.740 231.090 -129.540 ;
        RECT 231.950 -129.640 232.165 -128.420 ;
        RECT 233.135 -128.765 233.485 -122.080 ;
        RECT 234.475 -128.395 234.690 -118.520 ;
        RECT 236.110 -120.635 236.490 -117.115 ;
        RECT 237.620 -116.895 246.555 -116.705 ;
        RECT 237.620 -118.785 237.810 -116.895 ;
        RECT 243.655 -118.390 246.980 -118.250 ;
        RECT 243.655 -118.680 248.830 -118.390 ;
        RECT 237.505 -119.055 237.870 -118.785 ;
        RECT 243.655 -119.085 244.085 -118.680 ;
        RECT 244.955 -118.865 245.130 -118.680 ;
        RECT 246.580 -118.695 248.830 -118.680 ;
        RECT 239.395 -119.515 244.085 -119.085 ;
        RECT 238.635 -120.635 239.285 -120.505 ;
        RECT 236.110 -120.965 239.285 -120.635 ;
        RECT 240.095 -120.795 240.265 -119.515 ;
        RECT 240.585 -120.795 240.755 -119.755 ;
        RECT 241.075 -120.795 241.245 -119.515 ;
        RECT 241.565 -120.625 241.735 -119.755 ;
        RECT 244.470 -120.405 244.640 -118.865 ;
        RECT 244.960 -120.405 245.130 -118.865 ;
        RECT 245.450 -120.405 245.620 -118.865 ;
        RECT 245.940 -120.405 246.110 -118.865 ;
        RECT 246.430 -120.405 246.600 -118.865 ;
        RECT 244.310 -120.620 244.665 -120.615 ;
        RECT 246.370 -120.620 246.740 -120.590 ;
        RECT 244.310 -120.625 246.740 -120.620 ;
        RECT 241.565 -120.795 246.740 -120.625 ;
        RECT 248.525 -120.730 248.830 -118.695 ;
        RECT 241.570 -120.815 246.740 -120.795 ;
        RECT 241.570 -120.825 244.315 -120.815 ;
        RECT 239.505 -120.965 239.870 -120.935 ;
        RECT 246.370 -120.945 246.740 -120.815 ;
        RECT 236.110 -121.015 239.870 -120.965 ;
        RECT 238.635 -121.170 239.870 -121.015 ;
        RECT 244.045 -121.105 244.720 -121.065 ;
        RECT 243.945 -121.115 244.720 -121.105 ;
        RECT 238.635 -121.255 239.285 -121.170 ;
        RECT 239.505 -121.235 239.870 -121.170 ;
        RECT 238.770 -121.505 239.150 -121.255 ;
        RECT 242.910 -121.295 244.720 -121.115 ;
        RECT 247.305 -121.160 251.230 -120.730 ;
        RECT 243.945 -121.305 244.720 -121.295 ;
        RECT 244.045 -121.335 244.720 -121.305 ;
        RECT 244.960 -121.220 247.055 -121.180 ;
        RECT 244.960 -121.370 247.110 -121.220 ;
        RECT 240.095 -122.445 240.265 -121.405 ;
        RECT 241.075 -122.445 241.245 -121.405 ;
        RECT 242.055 -122.445 242.225 -121.405 ;
        RECT 244.960 -123.090 245.130 -121.370 ;
        RECT 245.940 -123.090 246.110 -121.370 ;
        RECT 246.805 -122.115 247.110 -121.370 ;
        RECT 248.005 -121.940 248.175 -121.160 ;
        RECT 248.495 -121.940 248.665 -121.400 ;
        RECT 248.985 -121.940 249.155 -121.160 ;
        RECT 249.475 -121.940 249.645 -121.400 ;
        RECT 247.415 -122.115 247.780 -122.085 ;
        RECT 246.805 -122.180 247.780 -122.115 ;
        RECT 246.915 -122.320 247.780 -122.180 ;
        RECT 247.415 -122.385 247.780 -122.320 ;
        RECT 249.965 -122.235 251.825 -121.885 ;
        RECT 248.005 -123.095 248.175 -122.555 ;
        RECT 248.985 -123.095 249.155 -122.555 ;
        RECT 249.965 -123.095 250.135 -122.235 ;
        RECT 248.235 -125.435 249.435 -125.265 ;
        RECT 239.965 -127.770 240.135 -126.050 ;
        RECT 240.945 -127.770 241.115 -126.050 ;
        RECT 243.010 -126.585 243.180 -126.045 ;
        RECT 243.990 -126.585 244.160 -126.045 ;
        RECT 242.420 -126.820 242.785 -126.755 ;
        RECT 241.920 -126.960 242.785 -126.820 ;
        RECT 241.810 -127.025 242.785 -126.960 ;
        RECT 241.810 -127.770 242.115 -127.025 ;
        RECT 242.420 -127.055 242.785 -127.025 ;
        RECT 244.970 -126.905 245.140 -126.045 ;
        RECT 239.965 -127.920 242.115 -127.770 ;
        RECT 239.965 -127.960 242.060 -127.920 ;
        RECT 243.010 -127.980 243.180 -127.200 ;
        RECT 243.500 -127.740 243.670 -127.200 ;
        RECT 243.990 -127.980 244.160 -127.200 ;
        RECT 244.480 -127.740 244.650 -127.200 ;
        RECT 244.970 -127.255 246.360 -126.905 ;
        RECT 238.185 -128.325 239.320 -128.315 ;
        RECT 241.375 -128.325 241.745 -128.195 ;
        RECT 234.475 -128.610 235.900 -128.395 ;
        RECT 238.185 -128.515 241.745 -128.325 ;
        RECT 242.310 -128.410 245.385 -127.980 ;
        RECT 239.315 -128.520 241.745 -128.515 ;
        RECT 239.315 -128.525 239.670 -128.520 ;
        RECT 241.375 -128.550 241.745 -128.520 ;
        RECT 233.080 -129.125 233.605 -128.765 ;
        RECT 235.685 -129.640 235.900 -128.610 ;
        RECT 223.245 -130.380 225.495 -130.290 ;
        RECT 221.035 -130.595 225.495 -130.380 ;
        RECT 221.035 -130.685 223.280 -130.595 ;
        RECT 225.190 -132.070 225.495 -130.595 ;
        RECT 228.860 -131.480 229.030 -130.010 ;
        RECT 229.320 -130.090 229.545 -129.740 ;
        RECT 231.280 -129.840 235.900 -129.640 ;
        RECT 231.520 -129.855 235.900 -129.840 ;
        RECT 228.825 -132.070 229.060 -131.480 ;
        RECT 229.350 -131.550 229.520 -130.090 ;
        RECT 229.840 -131.475 230.010 -130.010 ;
        RECT 231.050 -131.425 231.220 -130.010 ;
        RECT 231.520 -130.055 231.740 -129.855 ;
        RECT 229.805 -132.070 230.040 -131.475 ;
        RECT 231.015 -132.070 231.250 -131.425 ;
        RECT 231.540 -131.550 231.710 -130.055 ;
        RECT 239.475 -130.275 239.645 -128.735 ;
        RECT 239.965 -130.275 240.135 -128.735 ;
        RECT 240.455 -130.275 240.625 -128.735 ;
        RECT 240.945 -130.275 241.115 -128.735 ;
        RECT 241.435 -130.275 241.605 -128.735 ;
        RECT 239.960 -130.535 240.135 -130.275 ;
        RECT 243.530 -130.445 243.835 -128.410 ;
        RECT 245.980 -129.230 246.330 -127.255 ;
        RECT 247.200 -128.525 247.370 -125.605 ;
        RECT 248.235 -125.645 248.445 -125.435 ;
        RECT 247.180 -128.820 247.390 -128.525 ;
        RECT 248.255 -128.555 248.425 -125.645 ;
        RECT 248.745 -128.545 248.915 -125.605 ;
        RECT 249.225 -125.655 249.435 -125.435 ;
        RECT 248.240 -128.820 248.450 -128.555 ;
        RECT 247.180 -129.000 248.450 -128.820 ;
        RECT 248.725 -128.815 248.935 -128.545 ;
        RECT 249.235 -128.645 249.405 -125.655 ;
        RECT 250.295 -128.575 250.465 -125.605 ;
        RECT 248.725 -129.010 249.430 -128.815 ;
        RECT 249.215 -129.070 249.430 -129.010 ;
        RECT 248.005 -129.230 248.780 -129.180 ;
        RECT 245.980 -129.410 248.780 -129.230 ;
        RECT 245.980 -129.420 246.330 -129.410 ;
        RECT 248.005 -129.455 248.780 -129.410 ;
        RECT 249.215 -129.345 250.120 -129.070 ;
        RECT 249.215 -129.695 249.430 -129.345 ;
        RECT 246.655 -129.765 247.430 -129.720 ;
        RECT 246.470 -129.935 247.430 -129.765 ;
        RECT 246.655 -129.995 247.430 -129.935 ;
        RECT 247.660 -129.895 249.430 -129.695 ;
        RECT 250.290 -129.795 250.505 -128.575 ;
        RECT 251.475 -128.920 251.825 -122.235 ;
        RECT 251.420 -129.280 251.945 -128.920 ;
        RECT 254.070 -129.795 255.140 -129.220 ;
        RECT 241.585 -130.535 243.835 -130.445 ;
        RECT 239.375 -130.750 243.835 -130.535 ;
        RECT 239.375 -130.840 241.620 -130.750 ;
        RECT 225.190 -132.635 232.575 -132.070 ;
        RECT 243.530 -132.225 243.835 -130.750 ;
        RECT 247.200 -131.635 247.370 -130.165 ;
        RECT 247.660 -130.245 247.885 -129.895 ;
        RECT 249.620 -129.995 255.630 -129.795 ;
        RECT 249.860 -130.010 255.630 -129.995 ;
        RECT 247.165 -132.225 247.400 -131.635 ;
        RECT 247.690 -131.705 247.860 -130.245 ;
        RECT 248.180 -131.630 248.350 -130.165 ;
        RECT 249.390 -131.580 249.560 -130.165 ;
        RECT 249.860 -130.210 250.080 -130.010 ;
        RECT 248.145 -132.225 248.380 -131.630 ;
        RECT 249.355 -132.225 249.590 -131.580 ;
        RECT 249.880 -131.705 250.050 -130.210 ;
        RECT 254.070 -130.320 255.140 -130.010 ;
        RECT 243.530 -132.790 250.915 -132.225 ;
        RECT 261.000 -137.500 261.730 -110.660 ;
        RECT 265.875 -110.735 267.010 -110.725 ;
        RECT 269.065 -110.735 269.435 -110.605 ;
        RECT 265.875 -110.925 269.435 -110.735 ;
        RECT 270.000 -110.820 273.075 -110.390 ;
        RECT 265.930 -115.280 266.310 -110.925 ;
        RECT 267.005 -110.930 269.435 -110.925 ;
        RECT 267.005 -110.935 267.360 -110.930 ;
        RECT 269.065 -110.960 269.435 -110.930 ;
        RECT 267.165 -112.685 267.335 -111.145 ;
        RECT 267.655 -112.685 267.825 -111.145 ;
        RECT 268.145 -112.685 268.315 -111.145 ;
        RECT 268.635 -112.685 268.805 -111.145 ;
        RECT 269.125 -112.685 269.295 -111.145 ;
        RECT 267.650 -112.945 267.825 -112.685 ;
        RECT 271.220 -112.855 271.525 -110.820 ;
        RECT 273.670 -111.640 274.020 -109.665 ;
        RECT 274.890 -110.935 275.060 -108.015 ;
        RECT 275.925 -108.055 276.135 -107.845 ;
        RECT 274.870 -111.230 275.080 -110.935 ;
        RECT 275.945 -110.965 276.115 -108.055 ;
        RECT 276.435 -110.955 276.605 -108.015 ;
        RECT 276.915 -108.065 277.125 -107.845 ;
        RECT 275.930 -111.230 276.140 -110.965 ;
        RECT 274.870 -111.410 276.140 -111.230 ;
        RECT 276.415 -111.225 276.625 -110.955 ;
        RECT 276.925 -111.055 277.095 -108.065 ;
        RECT 277.985 -110.985 278.155 -108.015 ;
        RECT 276.415 -111.420 277.120 -111.225 ;
        RECT 276.905 -111.480 277.120 -111.420 ;
        RECT 275.695 -111.640 276.470 -111.590 ;
        RECT 273.670 -111.820 276.470 -111.640 ;
        RECT 273.670 -111.830 274.020 -111.820 ;
        RECT 275.695 -111.865 276.470 -111.820 ;
        RECT 276.905 -111.755 277.810 -111.480 ;
        RECT 276.905 -112.105 277.120 -111.755 ;
        RECT 274.345 -112.175 275.120 -112.130 ;
        RECT 274.160 -112.345 275.120 -112.175 ;
        RECT 274.345 -112.405 275.120 -112.345 ;
        RECT 275.350 -112.305 277.120 -112.105 ;
        RECT 277.980 -112.205 278.195 -110.985 ;
        RECT 279.165 -111.330 279.515 -104.645 ;
        RECT 316.420 -105.170 316.590 -103.450 ;
        RECT 317.400 -105.170 317.570 -103.450 ;
        RECT 318.265 -104.195 318.570 -103.450 ;
        RECT 319.465 -104.020 319.635 -103.240 ;
        RECT 319.955 -104.020 320.125 -103.480 ;
        RECT 320.445 -104.020 320.615 -103.240 ;
        RECT 355.860 -103.250 356.510 -103.165 ;
        RECT 356.730 -103.230 357.095 -103.165 ;
        RECT 360.135 -103.290 361.945 -103.110 ;
        RECT 364.530 -103.155 368.455 -102.725 ;
        RECT 402.680 -102.770 403.330 -102.310 ;
        RECT 404.140 -102.600 404.310 -101.320 ;
        RECT 404.630 -102.600 404.800 -101.560 ;
        RECT 405.120 -102.600 405.290 -101.320 ;
        RECT 405.610 -102.430 405.780 -101.560 ;
        RECT 408.515 -102.210 408.685 -100.670 ;
        RECT 409.005 -102.210 409.175 -100.670 ;
        RECT 409.495 -102.210 409.665 -100.670 ;
        RECT 409.985 -102.210 410.155 -100.670 ;
        RECT 410.475 -102.210 410.645 -100.670 ;
        RECT 408.355 -102.425 408.710 -102.420 ;
        RECT 410.415 -102.425 410.785 -102.395 ;
        RECT 408.355 -102.430 410.785 -102.425 ;
        RECT 405.610 -102.600 410.785 -102.430 ;
        RECT 412.570 -102.535 412.875 -100.500 ;
        RECT 405.615 -102.620 410.785 -102.600 ;
        RECT 405.615 -102.630 408.360 -102.620 ;
        RECT 403.550 -102.770 403.915 -102.740 ;
        RECT 410.415 -102.750 410.785 -102.620 ;
        RECT 402.680 -102.975 403.915 -102.770 ;
        RECT 408.090 -102.910 408.765 -102.870 ;
        RECT 407.990 -102.920 408.765 -102.910 ;
        RECT 402.680 -103.060 403.330 -102.975 ;
        RECT 403.550 -103.040 403.915 -102.975 ;
        RECT 406.955 -103.100 408.765 -102.920 ;
        RECT 411.350 -102.965 415.275 -102.535 ;
        RECT 407.990 -103.110 408.765 -103.100 ;
        RECT 408.090 -103.140 408.765 -103.110 ;
        RECT 409.005 -103.025 411.100 -102.985 ;
        RECT 361.170 -103.300 361.945 -103.290 ;
        RECT 361.270 -103.330 361.945 -103.300 ;
        RECT 362.185 -103.215 364.280 -103.175 ;
        RECT 362.185 -103.365 364.335 -103.215 ;
        RECT 320.935 -104.020 321.105 -103.480 ;
        RECT 318.875 -104.195 319.240 -104.165 ;
        RECT 318.265 -104.260 319.240 -104.195 ;
        RECT 318.375 -104.400 319.240 -104.260 ;
        RECT 318.875 -104.465 319.240 -104.400 ;
        RECT 321.425 -104.315 323.285 -103.965 ;
        RECT 319.465 -105.175 319.635 -104.635 ;
        RECT 320.445 -105.175 320.615 -104.635 ;
        RECT 321.425 -105.175 321.595 -104.315 ;
        RECT 285.745 -107.125 287.350 -106.955 ;
        RECT 284.850 -109.805 285.020 -107.305 ;
        RECT 284.845 -110.035 285.020 -109.805 ;
        RECT 285.745 -110.035 285.945 -107.125 ;
        RECT 286.190 -107.325 286.365 -107.125 ;
        RECT 286.195 -109.845 286.365 -107.325 ;
        RECT 286.685 -109.810 286.855 -107.305 ;
        RECT 287.175 -107.320 287.350 -107.125 ;
        RECT 284.845 -110.235 285.945 -110.035 ;
        RECT 286.670 -110.410 286.860 -109.810 ;
        RECT 287.175 -109.845 287.345 -107.320 ;
        RECT 287.825 -110.225 287.995 -107.305 ;
        RECT 289.455 -109.875 289.625 -107.305 ;
        RECT 290.595 -108.755 290.765 -107.305 ;
        RECT 319.695 -107.515 320.895 -107.345 ;
        RECT 290.590 -109.220 290.775 -108.755 ;
        RECT 290.590 -109.405 291.275 -109.220 ;
        RECT 289.455 -110.045 290.250 -109.875 ;
        RECT 288.570 -110.225 289.260 -110.170 ;
        RECT 284.850 -110.600 286.860 -110.410 ;
        RECT 287.195 -110.395 289.260 -110.225 ;
        RECT 283.665 -110.655 284.355 -110.605 ;
        RECT 281.715 -110.825 284.355 -110.655 ;
        RECT 279.110 -111.690 279.635 -111.330 ;
        RECT 281.715 -112.205 281.930 -110.825 ;
        RECT 283.665 -110.875 284.355 -110.825 ;
        RECT 283.945 -111.330 284.635 -111.285 ;
        RECT 282.895 -111.500 284.635 -111.330 ;
        RECT 282.895 -112.135 283.255 -111.500 ;
        RECT 283.945 -111.555 284.635 -111.500 ;
        RECT 282.895 -112.180 283.315 -112.135 ;
        RECT 269.275 -112.945 271.525 -112.855 ;
        RECT 267.065 -113.160 271.525 -112.945 ;
        RECT 267.065 -113.250 269.310 -113.160 ;
        RECT 271.220 -114.635 271.525 -113.160 ;
        RECT 274.890 -114.045 275.060 -112.575 ;
        RECT 275.350 -112.655 275.575 -112.305 ;
        RECT 277.310 -112.405 281.930 -112.205 ;
        RECT 277.550 -112.420 281.930 -112.405 ;
        RECT 274.855 -114.635 275.090 -114.045 ;
        RECT 275.380 -114.115 275.550 -112.655 ;
        RECT 275.870 -114.040 276.040 -112.575 ;
        RECT 277.080 -113.990 277.250 -112.575 ;
        RECT 277.550 -112.620 277.770 -112.420 ;
        RECT 282.920 -112.530 283.315 -112.180 ;
        RECT 275.835 -114.635 276.070 -114.040 ;
        RECT 277.045 -114.635 277.280 -113.990 ;
        RECT 277.570 -114.115 277.740 -112.620 ;
        RECT 284.360 -113.740 284.530 -112.285 ;
        RECT 284.350 -114.295 284.535 -113.740 ;
        RECT 284.850 -113.825 285.020 -110.600 ;
        RECT 285.995 -110.950 286.185 -110.600 ;
        RECT 287.195 -110.790 287.365 -110.395 ;
        RECT 288.570 -110.440 289.260 -110.395 ;
        RECT 285.945 -111.640 286.215 -110.950 ;
        RECT 286.710 -110.960 287.365 -110.790 ;
        RECT 287.695 -110.875 288.385 -110.605 ;
        RECT 289.620 -110.950 289.890 -110.260 ;
        RECT 290.080 -110.265 290.250 -110.045 ;
        RECT 290.080 -110.535 290.910 -110.265 ;
        RECT 286.710 -113.825 286.880 -110.960 ;
        RECT 290.080 -111.110 290.250 -110.535 ;
        RECT 290.510 -111.110 290.780 -111.025 ;
        RECT 287.200 -111.305 287.995 -111.130 ;
        RECT 290.080 -111.135 290.780 -111.110 ;
        RECT 289.940 -111.280 290.780 -111.135 ;
        RECT 287.200 -113.825 287.370 -111.305 ;
        RECT 287.825 -113.825 287.995 -111.305 ;
        RECT 288.315 -113.740 288.485 -111.285 ;
        RECT 288.965 -113.735 289.135 -111.285 ;
        RECT 281.665 -114.315 284.720 -114.295 ;
        RECT 288.310 -114.315 288.495 -113.740 ;
        RECT 288.950 -114.315 289.135 -113.735 ;
        RECT 289.455 -113.825 289.625 -111.285 ;
        RECT 289.940 -111.305 290.250 -111.280 ;
        RECT 289.945 -113.825 290.115 -111.305 ;
        RECT 290.510 -111.320 290.780 -111.280 ;
        RECT 291.085 -111.870 291.275 -109.405 ;
        RECT 303.635 -109.925 308.265 -109.305 ;
        RECT 311.425 -109.850 311.595 -108.130 ;
        RECT 312.405 -109.850 312.575 -108.130 ;
        RECT 314.470 -108.665 314.640 -108.125 ;
        RECT 315.450 -108.665 315.620 -108.125 ;
        RECT 313.880 -108.900 314.245 -108.835 ;
        RECT 313.380 -109.040 314.245 -108.900 ;
        RECT 313.270 -109.105 314.245 -109.040 ;
        RECT 313.270 -109.850 313.575 -109.105 ;
        RECT 313.880 -109.135 314.245 -109.105 ;
        RECT 316.430 -108.985 316.600 -108.125 ;
        RECT 310.510 -109.915 311.185 -109.885 ;
        RECT 310.410 -109.925 311.185 -109.915 ;
        RECT 303.635 -110.105 311.185 -109.925 ;
        RECT 311.425 -110.000 313.575 -109.850 ;
        RECT 311.425 -110.040 313.520 -110.000 ;
        RECT 314.470 -110.060 314.640 -109.280 ;
        RECT 314.960 -109.820 315.130 -109.280 ;
        RECT 315.450 -110.060 315.620 -109.280 ;
        RECT 315.940 -109.820 316.110 -109.280 ;
        RECT 316.430 -109.335 317.820 -108.985 ;
        RECT 303.635 -110.500 308.265 -110.105 ;
        RECT 310.410 -110.115 311.185 -110.105 ;
        RECT 310.510 -110.155 311.185 -110.115 ;
        RECT 309.645 -110.405 310.780 -110.395 ;
        RECT 312.835 -110.405 313.205 -110.275 ;
        RECT 291.085 -112.060 292.545 -111.870 ;
        RECT 290.595 -113.730 290.765 -112.285 ;
        RECT 291.085 -112.310 291.275 -112.060 ;
        RECT 290.585 -114.315 290.770 -113.730 ;
        RECT 291.085 -113.825 291.255 -112.310 ;
        RECT 281.665 -114.635 291.335 -114.315 ;
        RECT 271.220 -114.860 291.335 -114.635 ;
        RECT 271.220 -115.200 282.230 -114.860 ;
        RECT 283.970 -115.120 291.335 -114.860 ;
        RECT 262.375 -116.085 266.310 -115.280 ;
        RECT 262.375 -135.690 263.180 -116.085 ;
        RECT 265.930 -116.565 266.310 -116.085 ;
        RECT 292.355 -116.535 292.545 -112.060 ;
        RECT 265.930 -116.945 282.480 -116.565 ;
        RECT 265.930 -117.855 266.310 -116.945 ;
        RECT 265.930 -118.235 266.640 -117.855 ;
        RECT 266.260 -120.180 266.640 -118.235 ;
        RECT 271.305 -118.065 274.630 -117.925 ;
        RECT 271.305 -118.355 276.480 -118.065 ;
        RECT 280.350 -118.350 280.810 -117.925 ;
        RECT 271.305 -118.760 271.735 -118.355 ;
        RECT 272.605 -118.540 272.780 -118.355 ;
        RECT 274.230 -118.370 276.480 -118.355 ;
        RECT 267.045 -119.190 271.735 -118.760 ;
        RECT 266.260 -120.640 266.935 -120.180 ;
        RECT 267.745 -120.470 267.915 -119.190 ;
        RECT 268.235 -120.470 268.405 -119.430 ;
        RECT 268.725 -120.470 268.895 -119.190 ;
        RECT 269.215 -120.300 269.385 -119.430 ;
        RECT 272.120 -120.080 272.290 -118.540 ;
        RECT 272.610 -120.080 272.780 -118.540 ;
        RECT 273.100 -120.080 273.270 -118.540 ;
        RECT 273.590 -120.080 273.760 -118.540 ;
        RECT 274.080 -120.080 274.250 -118.540 ;
        RECT 271.960 -120.295 272.315 -120.290 ;
        RECT 274.020 -120.295 274.390 -120.265 ;
        RECT 271.960 -120.300 274.390 -120.295 ;
        RECT 269.215 -120.470 274.390 -120.300 ;
        RECT 276.175 -120.405 276.480 -118.370 ;
        RECT 269.220 -120.490 274.390 -120.470 ;
        RECT 269.220 -120.500 271.965 -120.490 ;
        RECT 267.155 -120.640 267.520 -120.610 ;
        RECT 274.020 -120.620 274.390 -120.490 ;
        RECT 266.260 -120.725 267.520 -120.640 ;
        RECT 266.285 -120.845 267.520 -120.725 ;
        RECT 271.695 -120.780 272.370 -120.740 ;
        RECT 271.595 -120.790 272.370 -120.780 ;
        RECT 266.285 -120.930 266.935 -120.845 ;
        RECT 267.155 -120.910 267.520 -120.845 ;
        RECT 270.560 -120.970 272.370 -120.790 ;
        RECT 274.955 -120.835 278.880 -120.405 ;
        RECT 271.595 -120.980 272.370 -120.970 ;
        RECT 271.695 -121.010 272.370 -120.980 ;
        RECT 272.610 -120.895 274.705 -120.855 ;
        RECT 272.610 -121.045 274.760 -120.895 ;
        RECT 267.745 -122.120 267.915 -121.080 ;
        RECT 268.725 -122.120 268.895 -121.080 ;
        RECT 269.705 -122.120 269.875 -121.080 ;
        RECT 272.610 -122.765 272.780 -121.045 ;
        RECT 273.590 -122.765 273.760 -121.045 ;
        RECT 274.455 -121.790 274.760 -121.045 ;
        RECT 275.655 -121.615 275.825 -120.835 ;
        RECT 276.145 -121.615 276.315 -121.075 ;
        RECT 276.635 -121.615 276.805 -120.835 ;
        RECT 277.125 -121.615 277.295 -121.075 ;
        RECT 275.065 -121.790 275.430 -121.760 ;
        RECT 274.455 -121.855 275.430 -121.790 ;
        RECT 274.565 -121.995 275.430 -121.855 ;
        RECT 275.065 -122.060 275.430 -121.995 ;
        RECT 277.615 -121.910 279.475 -121.560 ;
        RECT 275.655 -122.770 275.825 -122.230 ;
        RECT 276.635 -122.770 276.805 -122.230 ;
        RECT 277.615 -122.770 277.785 -121.910 ;
        RECT 275.885 -125.110 277.085 -124.940 ;
        RECT 267.615 -127.445 267.785 -125.725 ;
        RECT 268.595 -127.445 268.765 -125.725 ;
        RECT 270.660 -126.260 270.830 -125.720 ;
        RECT 271.640 -126.260 271.810 -125.720 ;
        RECT 270.070 -126.495 270.435 -126.430 ;
        RECT 269.570 -126.635 270.435 -126.495 ;
        RECT 269.460 -126.700 270.435 -126.635 ;
        RECT 269.460 -127.445 269.765 -126.700 ;
        RECT 270.070 -126.730 270.435 -126.700 ;
        RECT 272.620 -126.580 272.790 -125.720 ;
        RECT 267.615 -127.595 269.765 -127.445 ;
        RECT 267.615 -127.635 269.710 -127.595 ;
        RECT 270.660 -127.655 270.830 -126.875 ;
        RECT 271.150 -127.415 271.320 -126.875 ;
        RECT 271.640 -127.655 271.810 -126.875 ;
        RECT 272.130 -127.415 272.300 -126.875 ;
        RECT 272.620 -126.930 274.010 -126.580 ;
        RECT 265.835 -128.000 266.970 -127.990 ;
        RECT 269.025 -128.000 269.395 -127.870 ;
        RECT 265.835 -128.190 269.395 -128.000 ;
        RECT 269.960 -128.085 273.035 -127.655 ;
        RECT 266.965 -128.195 269.395 -128.190 ;
        RECT 266.965 -128.200 267.320 -128.195 ;
        RECT 269.025 -128.225 269.395 -128.195 ;
        RECT 267.125 -129.950 267.295 -128.410 ;
        RECT 267.615 -129.950 267.785 -128.410 ;
        RECT 268.105 -129.950 268.275 -128.410 ;
        RECT 268.595 -129.950 268.765 -128.410 ;
        RECT 269.085 -129.950 269.255 -128.410 ;
        RECT 267.610 -130.210 267.785 -129.950 ;
        RECT 271.180 -130.120 271.485 -128.085 ;
        RECT 273.630 -128.905 273.980 -126.930 ;
        RECT 274.850 -128.200 275.020 -125.280 ;
        RECT 275.885 -125.320 276.095 -125.110 ;
        RECT 274.830 -128.495 275.040 -128.200 ;
        RECT 275.905 -128.230 276.075 -125.320 ;
        RECT 276.395 -128.220 276.565 -125.280 ;
        RECT 276.875 -125.330 277.085 -125.110 ;
        RECT 275.890 -128.495 276.100 -128.230 ;
        RECT 274.830 -128.675 276.100 -128.495 ;
        RECT 276.375 -128.490 276.585 -128.220 ;
        RECT 276.885 -128.320 277.055 -125.330 ;
        RECT 277.945 -128.250 278.115 -125.280 ;
        RECT 276.375 -128.685 277.080 -128.490 ;
        RECT 276.865 -128.745 277.080 -128.685 ;
        RECT 275.655 -128.905 276.430 -128.855 ;
        RECT 273.630 -129.085 276.430 -128.905 ;
        RECT 273.630 -129.095 273.980 -129.085 ;
        RECT 275.655 -129.130 276.430 -129.085 ;
        RECT 276.865 -129.020 277.770 -128.745 ;
        RECT 276.865 -129.370 277.080 -129.020 ;
        RECT 274.305 -129.440 275.080 -129.395 ;
        RECT 274.120 -129.610 275.080 -129.440 ;
        RECT 274.305 -129.670 275.080 -129.610 ;
        RECT 275.310 -129.570 277.080 -129.370 ;
        RECT 277.940 -129.470 278.155 -128.250 ;
        RECT 279.125 -128.595 279.475 -121.910 ;
        RECT 280.465 -128.225 280.680 -118.350 ;
        RECT 282.100 -120.465 282.480 -116.945 ;
        RECT 283.610 -116.725 292.545 -116.535 ;
        RECT 283.610 -118.615 283.800 -116.725 ;
        RECT 289.645 -118.220 292.970 -118.080 ;
        RECT 289.645 -118.510 294.820 -118.220 ;
        RECT 283.495 -118.885 283.860 -118.615 ;
        RECT 289.645 -118.915 290.075 -118.510 ;
        RECT 290.945 -118.695 291.120 -118.510 ;
        RECT 292.570 -118.525 294.820 -118.510 ;
        RECT 285.385 -119.345 290.075 -118.915 ;
        RECT 284.625 -120.465 285.275 -120.335 ;
        RECT 282.100 -120.795 285.275 -120.465 ;
        RECT 286.085 -120.625 286.255 -119.345 ;
        RECT 286.575 -120.625 286.745 -119.585 ;
        RECT 287.065 -120.625 287.235 -119.345 ;
        RECT 287.555 -120.455 287.725 -119.585 ;
        RECT 290.460 -120.235 290.630 -118.695 ;
        RECT 290.950 -120.235 291.120 -118.695 ;
        RECT 291.440 -120.235 291.610 -118.695 ;
        RECT 291.930 -120.235 292.100 -118.695 ;
        RECT 292.420 -120.235 292.590 -118.695 ;
        RECT 290.300 -120.450 290.655 -120.445 ;
        RECT 292.360 -120.450 292.730 -120.420 ;
        RECT 290.300 -120.455 292.730 -120.450 ;
        RECT 287.555 -120.625 292.730 -120.455 ;
        RECT 294.515 -120.560 294.820 -118.525 ;
        RECT 287.560 -120.645 292.730 -120.625 ;
        RECT 287.560 -120.655 290.305 -120.645 ;
        RECT 285.495 -120.795 285.860 -120.765 ;
        RECT 292.360 -120.775 292.730 -120.645 ;
        RECT 282.100 -120.845 285.860 -120.795 ;
        RECT 284.625 -121.000 285.860 -120.845 ;
        RECT 290.035 -120.935 290.710 -120.895 ;
        RECT 289.935 -120.945 290.710 -120.935 ;
        RECT 284.625 -121.085 285.275 -121.000 ;
        RECT 285.495 -121.065 285.860 -121.000 ;
        RECT 284.760 -121.335 285.140 -121.085 ;
        RECT 288.900 -121.125 290.710 -120.945 ;
        RECT 293.295 -120.990 297.220 -120.560 ;
        RECT 289.935 -121.135 290.710 -121.125 ;
        RECT 290.035 -121.165 290.710 -121.135 ;
        RECT 290.950 -121.050 293.045 -121.010 ;
        RECT 290.950 -121.200 293.100 -121.050 ;
        RECT 286.085 -122.275 286.255 -121.235 ;
        RECT 287.065 -122.275 287.235 -121.235 ;
        RECT 288.045 -122.275 288.215 -121.235 ;
        RECT 290.950 -122.920 291.120 -121.200 ;
        RECT 291.930 -122.920 292.100 -121.200 ;
        RECT 292.795 -121.945 293.100 -121.200 ;
        RECT 293.995 -121.770 294.165 -120.990 ;
        RECT 294.485 -121.770 294.655 -121.230 ;
        RECT 294.975 -121.770 295.145 -120.990 ;
        RECT 295.465 -121.770 295.635 -121.230 ;
        RECT 293.405 -121.945 293.770 -121.915 ;
        RECT 292.795 -122.010 293.770 -121.945 ;
        RECT 292.905 -122.150 293.770 -122.010 ;
        RECT 293.405 -122.215 293.770 -122.150 ;
        RECT 295.955 -122.065 297.815 -121.715 ;
        RECT 293.995 -122.925 294.165 -122.385 ;
        RECT 294.975 -122.925 295.145 -122.385 ;
        RECT 295.955 -122.925 296.125 -122.065 ;
        RECT 294.225 -125.265 295.425 -125.095 ;
        RECT 285.955 -127.600 286.125 -125.880 ;
        RECT 286.935 -127.600 287.105 -125.880 ;
        RECT 289.000 -126.415 289.170 -125.875 ;
        RECT 289.980 -126.415 290.150 -125.875 ;
        RECT 288.410 -126.650 288.775 -126.585 ;
        RECT 287.910 -126.790 288.775 -126.650 ;
        RECT 287.800 -126.855 288.775 -126.790 ;
        RECT 287.800 -127.600 288.105 -126.855 ;
        RECT 288.410 -126.885 288.775 -126.855 ;
        RECT 290.960 -126.735 291.130 -125.875 ;
        RECT 285.955 -127.750 288.105 -127.600 ;
        RECT 285.955 -127.790 288.050 -127.750 ;
        RECT 289.000 -127.810 289.170 -127.030 ;
        RECT 289.490 -127.570 289.660 -127.030 ;
        RECT 289.980 -127.810 290.150 -127.030 ;
        RECT 290.470 -127.570 290.640 -127.030 ;
        RECT 290.960 -127.085 292.350 -126.735 ;
        RECT 284.175 -128.155 285.310 -128.145 ;
        RECT 287.365 -128.155 287.735 -128.025 ;
        RECT 280.465 -128.440 281.890 -128.225 ;
        RECT 284.175 -128.345 287.735 -128.155 ;
        RECT 288.300 -128.240 291.375 -127.810 ;
        RECT 285.305 -128.350 287.735 -128.345 ;
        RECT 285.305 -128.355 285.660 -128.350 ;
        RECT 287.365 -128.380 287.735 -128.350 ;
        RECT 279.070 -128.955 279.595 -128.595 ;
        RECT 281.675 -129.470 281.890 -128.440 ;
        RECT 269.235 -130.210 271.485 -130.120 ;
        RECT 267.025 -130.425 271.485 -130.210 ;
        RECT 267.025 -130.515 269.270 -130.425 ;
        RECT 271.180 -131.900 271.485 -130.425 ;
        RECT 274.850 -131.310 275.020 -129.840 ;
        RECT 275.310 -129.920 275.535 -129.570 ;
        RECT 277.270 -129.670 281.890 -129.470 ;
        RECT 277.510 -129.685 281.890 -129.670 ;
        RECT 274.815 -131.900 275.050 -131.310 ;
        RECT 275.340 -131.380 275.510 -129.920 ;
        RECT 275.830 -131.305 276.000 -129.840 ;
        RECT 277.040 -131.255 277.210 -129.840 ;
        RECT 277.510 -129.885 277.730 -129.685 ;
        RECT 275.795 -131.900 276.030 -131.305 ;
        RECT 277.005 -131.900 277.240 -131.255 ;
        RECT 277.530 -131.380 277.700 -129.885 ;
        RECT 285.465 -130.105 285.635 -128.565 ;
        RECT 285.955 -130.105 286.125 -128.565 ;
        RECT 286.445 -130.105 286.615 -128.565 ;
        RECT 286.935 -130.105 287.105 -128.565 ;
        RECT 287.425 -130.105 287.595 -128.565 ;
        RECT 285.950 -130.365 286.125 -130.105 ;
        RECT 289.520 -130.275 289.825 -128.240 ;
        RECT 291.970 -129.060 292.320 -127.085 ;
        RECT 293.190 -128.355 293.360 -125.435 ;
        RECT 294.225 -125.475 294.435 -125.265 ;
        RECT 293.170 -128.650 293.380 -128.355 ;
        RECT 294.245 -128.385 294.415 -125.475 ;
        RECT 294.735 -128.375 294.905 -125.435 ;
        RECT 295.215 -125.485 295.425 -125.265 ;
        RECT 294.230 -128.650 294.440 -128.385 ;
        RECT 293.170 -128.830 294.440 -128.650 ;
        RECT 294.715 -128.645 294.925 -128.375 ;
        RECT 295.225 -128.475 295.395 -125.485 ;
        RECT 296.285 -128.405 296.455 -125.435 ;
        RECT 294.715 -128.840 295.420 -128.645 ;
        RECT 295.205 -128.900 295.420 -128.840 ;
        RECT 293.995 -129.060 294.770 -129.010 ;
        RECT 291.970 -129.240 294.770 -129.060 ;
        RECT 291.970 -129.250 292.320 -129.240 ;
        RECT 293.995 -129.285 294.770 -129.240 ;
        RECT 295.205 -129.175 296.110 -128.900 ;
        RECT 295.205 -129.525 295.420 -129.175 ;
        RECT 292.645 -129.595 293.420 -129.550 ;
        RECT 292.460 -129.765 293.420 -129.595 ;
        RECT 292.645 -129.825 293.420 -129.765 ;
        RECT 293.650 -129.725 295.420 -129.525 ;
        RECT 296.280 -129.625 296.495 -128.405 ;
        RECT 297.465 -128.750 297.815 -122.065 ;
        RECT 297.410 -129.110 297.935 -128.750 ;
        RECT 299.700 -129.625 301.160 -128.780 ;
        RECT 287.575 -130.365 289.825 -130.275 ;
        RECT 285.365 -130.580 289.825 -130.365 ;
        RECT 285.365 -130.670 287.610 -130.580 ;
        RECT 271.180 -132.465 278.565 -131.900 ;
        RECT 289.520 -132.055 289.825 -130.580 ;
        RECT 293.190 -131.465 293.360 -129.995 ;
        RECT 293.650 -130.075 293.875 -129.725 ;
        RECT 295.610 -129.825 301.620 -129.625 ;
        RECT 295.850 -129.840 301.620 -129.825 ;
        RECT 293.155 -132.055 293.390 -131.465 ;
        RECT 293.680 -131.535 293.850 -130.075 ;
        RECT 294.170 -131.460 294.340 -129.995 ;
        RECT 295.380 -131.410 295.550 -129.995 ;
        RECT 295.850 -130.040 296.070 -129.840 ;
        RECT 294.135 -132.055 294.370 -131.460 ;
        RECT 295.345 -132.055 295.580 -131.410 ;
        RECT 295.870 -131.535 296.040 -130.040 ;
        RECT 299.700 -130.275 301.160 -129.840 ;
        RECT 289.520 -132.620 296.905 -132.055 ;
        RECT 262.285 -136.525 263.255 -135.690 ;
        RECT 303.635 -137.425 304.830 -110.500 ;
        RECT 309.645 -110.595 313.205 -110.405 ;
        RECT 313.770 -110.490 316.845 -110.060 ;
        RECT 309.700 -115.415 310.080 -110.595 ;
        RECT 310.775 -110.600 313.205 -110.595 ;
        RECT 310.775 -110.605 311.130 -110.600 ;
        RECT 312.835 -110.630 313.205 -110.600 ;
        RECT 310.935 -112.355 311.105 -110.815 ;
        RECT 311.425 -112.355 311.595 -110.815 ;
        RECT 311.915 -112.355 312.085 -110.815 ;
        RECT 312.405 -112.355 312.575 -110.815 ;
        RECT 312.895 -112.355 313.065 -110.815 ;
        RECT 311.420 -112.615 311.595 -112.355 ;
        RECT 314.990 -112.525 315.295 -110.490 ;
        RECT 317.440 -111.310 317.790 -109.335 ;
        RECT 318.660 -110.605 318.830 -107.685 ;
        RECT 319.695 -107.725 319.905 -107.515 ;
        RECT 318.640 -110.900 318.850 -110.605 ;
        RECT 319.715 -110.635 319.885 -107.725 ;
        RECT 320.205 -110.625 320.375 -107.685 ;
        RECT 320.685 -107.735 320.895 -107.515 ;
        RECT 319.700 -110.900 319.910 -110.635 ;
        RECT 318.640 -111.080 319.910 -110.900 ;
        RECT 320.185 -110.895 320.395 -110.625 ;
        RECT 320.695 -110.725 320.865 -107.735 ;
        RECT 321.755 -110.655 321.925 -107.685 ;
        RECT 320.185 -111.090 320.890 -110.895 ;
        RECT 320.675 -111.150 320.890 -111.090 ;
        RECT 319.465 -111.310 320.240 -111.260 ;
        RECT 317.440 -111.490 320.240 -111.310 ;
        RECT 317.440 -111.500 317.790 -111.490 ;
        RECT 319.465 -111.535 320.240 -111.490 ;
        RECT 320.675 -111.425 321.580 -111.150 ;
        RECT 320.675 -111.775 320.890 -111.425 ;
        RECT 318.115 -111.845 318.890 -111.800 ;
        RECT 317.930 -112.015 318.890 -111.845 ;
        RECT 318.115 -112.075 318.890 -112.015 ;
        RECT 319.120 -111.975 320.890 -111.775 ;
        RECT 321.750 -111.875 321.965 -110.655 ;
        RECT 322.935 -111.000 323.285 -104.315 ;
        RECT 357.320 -104.440 357.490 -103.400 ;
        RECT 358.300 -104.440 358.470 -103.400 ;
        RECT 359.280 -104.440 359.450 -103.400 ;
        RECT 362.185 -105.085 362.355 -103.365 ;
        RECT 363.165 -105.085 363.335 -103.365 ;
        RECT 364.030 -104.110 364.335 -103.365 ;
        RECT 365.230 -103.935 365.400 -103.155 ;
        RECT 365.720 -103.935 365.890 -103.395 ;
        RECT 366.210 -103.935 366.380 -103.155 ;
        RECT 409.005 -103.175 411.155 -103.025 ;
        RECT 366.700 -103.935 366.870 -103.395 ;
        RECT 364.640 -104.110 365.005 -104.080 ;
        RECT 364.030 -104.175 365.005 -104.110 ;
        RECT 364.140 -104.315 365.005 -104.175 ;
        RECT 364.640 -104.380 365.005 -104.315 ;
        RECT 367.190 -104.230 369.050 -103.880 ;
        RECT 365.230 -105.090 365.400 -104.550 ;
        RECT 366.210 -105.090 366.380 -104.550 ;
        RECT 367.190 -105.090 367.360 -104.230 ;
        RECT 329.515 -106.795 331.120 -106.625 ;
        RECT 328.620 -109.475 328.790 -106.975 ;
        RECT 328.615 -109.705 328.790 -109.475 ;
        RECT 329.515 -109.705 329.715 -106.795 ;
        RECT 329.960 -106.995 330.135 -106.795 ;
        RECT 329.965 -109.515 330.135 -106.995 ;
        RECT 330.455 -109.480 330.625 -106.975 ;
        RECT 330.945 -106.990 331.120 -106.795 ;
        RECT 328.615 -109.905 329.715 -109.705 ;
        RECT 330.440 -110.080 330.630 -109.480 ;
        RECT 330.945 -109.515 331.115 -106.990 ;
        RECT 331.595 -109.895 331.765 -106.975 ;
        RECT 333.225 -109.545 333.395 -106.975 ;
        RECT 334.365 -108.425 334.535 -106.975 ;
        RECT 365.460 -107.430 366.660 -107.260 ;
        RECT 334.360 -108.890 334.545 -108.425 ;
        RECT 334.360 -109.075 335.045 -108.890 ;
        RECT 333.225 -109.715 334.020 -109.545 ;
        RECT 332.340 -109.895 333.030 -109.840 ;
        RECT 328.620 -110.270 330.630 -110.080 ;
        RECT 330.965 -110.065 333.030 -109.895 ;
        RECT 327.435 -110.325 328.125 -110.275 ;
        RECT 325.485 -110.495 328.125 -110.325 ;
        RECT 322.880 -111.360 323.405 -111.000 ;
        RECT 325.485 -111.875 325.700 -110.495 ;
        RECT 327.435 -110.545 328.125 -110.495 ;
        RECT 327.715 -111.000 328.405 -110.955 ;
        RECT 326.665 -111.170 328.405 -111.000 ;
        RECT 326.665 -111.805 327.025 -111.170 ;
        RECT 327.715 -111.225 328.405 -111.170 ;
        RECT 326.665 -111.850 327.085 -111.805 ;
        RECT 313.045 -112.615 315.295 -112.525 ;
        RECT 310.835 -112.830 315.295 -112.615 ;
        RECT 310.835 -112.920 313.080 -112.830 ;
        RECT 314.990 -114.305 315.295 -112.830 ;
        RECT 318.660 -113.715 318.830 -112.245 ;
        RECT 319.120 -112.325 319.345 -111.975 ;
        RECT 321.080 -112.075 325.700 -111.875 ;
        RECT 321.320 -112.090 325.700 -112.075 ;
        RECT 318.625 -114.305 318.860 -113.715 ;
        RECT 319.150 -113.785 319.320 -112.325 ;
        RECT 319.640 -113.710 319.810 -112.245 ;
        RECT 320.850 -113.660 321.020 -112.245 ;
        RECT 321.320 -112.290 321.540 -112.090 ;
        RECT 326.690 -112.200 327.085 -111.850 ;
        RECT 319.605 -114.305 319.840 -113.710 ;
        RECT 320.815 -114.305 321.050 -113.660 ;
        RECT 321.340 -113.785 321.510 -112.290 ;
        RECT 328.130 -113.410 328.300 -111.955 ;
        RECT 328.120 -113.965 328.305 -113.410 ;
        RECT 328.620 -113.495 328.790 -110.270 ;
        RECT 329.765 -110.620 329.955 -110.270 ;
        RECT 330.965 -110.460 331.135 -110.065 ;
        RECT 332.340 -110.110 333.030 -110.065 ;
        RECT 329.715 -111.310 329.985 -110.620 ;
        RECT 330.480 -110.630 331.135 -110.460 ;
        RECT 331.465 -110.545 332.155 -110.275 ;
        RECT 333.390 -110.620 333.660 -109.930 ;
        RECT 333.850 -109.935 334.020 -109.715 ;
        RECT 333.850 -110.205 334.680 -109.935 ;
        RECT 330.480 -113.495 330.650 -110.630 ;
        RECT 333.850 -110.780 334.020 -110.205 ;
        RECT 334.280 -110.780 334.550 -110.695 ;
        RECT 330.970 -110.975 331.765 -110.800 ;
        RECT 333.850 -110.805 334.550 -110.780 ;
        RECT 333.710 -110.950 334.550 -110.805 ;
        RECT 330.970 -113.495 331.140 -110.975 ;
        RECT 331.595 -113.495 331.765 -110.975 ;
        RECT 332.085 -113.410 332.255 -110.955 ;
        RECT 332.735 -113.405 332.905 -110.955 ;
        RECT 325.435 -113.985 328.490 -113.965 ;
        RECT 332.080 -113.985 332.265 -113.410 ;
        RECT 332.720 -113.985 332.905 -113.405 ;
        RECT 333.225 -113.495 333.395 -110.955 ;
        RECT 333.710 -110.975 334.020 -110.950 ;
        RECT 333.715 -113.495 333.885 -110.975 ;
        RECT 334.280 -110.990 334.550 -110.950 ;
        RECT 334.855 -111.540 335.045 -109.075 ;
        RECT 350.275 -109.840 353.595 -109.445 ;
        RECT 357.190 -109.765 357.360 -108.045 ;
        RECT 358.170 -109.765 358.340 -108.045 ;
        RECT 360.235 -108.580 360.405 -108.040 ;
        RECT 361.215 -108.580 361.385 -108.040 ;
        RECT 359.645 -108.815 360.010 -108.750 ;
        RECT 359.145 -108.955 360.010 -108.815 ;
        RECT 359.035 -109.020 360.010 -108.955 ;
        RECT 359.035 -109.765 359.340 -109.020 ;
        RECT 359.645 -109.050 360.010 -109.020 ;
        RECT 362.195 -108.900 362.365 -108.040 ;
        RECT 356.275 -109.830 356.950 -109.800 ;
        RECT 356.175 -109.840 356.950 -109.830 ;
        RECT 350.275 -110.020 356.950 -109.840 ;
        RECT 357.190 -109.915 359.340 -109.765 ;
        RECT 357.190 -109.955 359.285 -109.915 ;
        RECT 360.235 -109.975 360.405 -109.195 ;
        RECT 360.725 -109.735 360.895 -109.195 ;
        RECT 361.215 -109.975 361.385 -109.195 ;
        RECT 361.705 -109.735 361.875 -109.195 ;
        RECT 362.195 -109.250 363.585 -108.900 ;
        RECT 350.275 -110.370 353.595 -110.020 ;
        RECT 356.175 -110.030 356.950 -110.020 ;
        RECT 356.275 -110.070 356.950 -110.030 ;
        RECT 355.410 -110.320 356.545 -110.310 ;
        RECT 358.600 -110.320 358.970 -110.190 ;
        RECT 334.855 -111.730 336.315 -111.540 ;
        RECT 334.365 -113.400 334.535 -111.955 ;
        RECT 334.855 -111.980 335.045 -111.730 ;
        RECT 334.355 -113.985 334.540 -113.400 ;
        RECT 334.855 -113.495 335.025 -111.980 ;
        RECT 325.435 -114.305 335.105 -113.985 ;
        RECT 314.990 -114.530 335.105 -114.305 ;
        RECT 314.990 -114.870 326.000 -114.530 ;
        RECT 327.740 -114.790 335.105 -114.530 ;
        RECT 306.135 -116.235 310.080 -115.415 ;
        RECT 336.125 -116.205 336.315 -111.730 ;
        RECT 306.135 -116.500 326.250 -116.235 ;
        RECT 214.135 -138.390 215.395 -137.695 ;
        RECT 260.830 -138.525 261.990 -137.500 ;
        RECT 303.325 -138.585 305.065 -137.425 ;
        RECT 306.135 -139.350 307.220 -116.500 ;
        RECT 309.700 -116.615 326.250 -116.500 ;
        RECT 309.700 -117.525 310.080 -116.615 ;
        RECT 309.700 -117.905 310.410 -117.525 ;
        RECT 310.030 -119.850 310.410 -117.905 ;
        RECT 315.075 -117.735 318.400 -117.595 ;
        RECT 315.075 -118.025 320.250 -117.735 ;
        RECT 324.120 -118.020 324.580 -117.595 ;
        RECT 315.075 -118.430 315.505 -118.025 ;
        RECT 316.375 -118.210 316.550 -118.025 ;
        RECT 318.000 -118.040 320.250 -118.025 ;
        RECT 310.815 -118.860 315.505 -118.430 ;
        RECT 310.030 -120.310 310.705 -119.850 ;
        RECT 311.515 -120.140 311.685 -118.860 ;
        RECT 312.005 -120.140 312.175 -119.100 ;
        RECT 312.495 -120.140 312.665 -118.860 ;
        RECT 312.985 -119.970 313.155 -119.100 ;
        RECT 315.890 -119.750 316.060 -118.210 ;
        RECT 316.380 -119.750 316.550 -118.210 ;
        RECT 316.870 -119.750 317.040 -118.210 ;
        RECT 317.360 -119.750 317.530 -118.210 ;
        RECT 317.850 -119.750 318.020 -118.210 ;
        RECT 315.730 -119.965 316.085 -119.960 ;
        RECT 317.790 -119.965 318.160 -119.935 ;
        RECT 315.730 -119.970 318.160 -119.965 ;
        RECT 312.985 -120.140 318.160 -119.970 ;
        RECT 319.945 -120.075 320.250 -118.040 ;
        RECT 312.990 -120.160 318.160 -120.140 ;
        RECT 312.990 -120.170 315.735 -120.160 ;
        RECT 310.925 -120.310 311.290 -120.280 ;
        RECT 317.790 -120.290 318.160 -120.160 ;
        RECT 310.030 -120.395 311.290 -120.310 ;
        RECT 310.055 -120.515 311.290 -120.395 ;
        RECT 315.465 -120.450 316.140 -120.410 ;
        RECT 315.365 -120.460 316.140 -120.450 ;
        RECT 310.055 -120.600 310.705 -120.515 ;
        RECT 310.925 -120.580 311.290 -120.515 ;
        RECT 314.330 -120.640 316.140 -120.460 ;
        RECT 318.725 -120.505 322.650 -120.075 ;
        RECT 315.365 -120.650 316.140 -120.640 ;
        RECT 315.465 -120.680 316.140 -120.650 ;
        RECT 316.380 -120.565 318.475 -120.525 ;
        RECT 316.380 -120.715 318.530 -120.565 ;
        RECT 311.515 -121.790 311.685 -120.750 ;
        RECT 312.495 -121.790 312.665 -120.750 ;
        RECT 313.475 -121.790 313.645 -120.750 ;
        RECT 316.380 -122.435 316.550 -120.715 ;
        RECT 317.360 -122.435 317.530 -120.715 ;
        RECT 318.225 -121.460 318.530 -120.715 ;
        RECT 319.425 -121.285 319.595 -120.505 ;
        RECT 319.915 -121.285 320.085 -120.745 ;
        RECT 320.405 -121.285 320.575 -120.505 ;
        RECT 320.895 -121.285 321.065 -120.745 ;
        RECT 318.835 -121.460 319.200 -121.430 ;
        RECT 318.225 -121.525 319.200 -121.460 ;
        RECT 318.335 -121.665 319.200 -121.525 ;
        RECT 318.835 -121.730 319.200 -121.665 ;
        RECT 321.385 -121.580 323.245 -121.230 ;
        RECT 319.425 -122.440 319.595 -121.900 ;
        RECT 320.405 -122.440 320.575 -121.900 ;
        RECT 321.385 -122.440 321.555 -121.580 ;
        RECT 319.655 -124.780 320.855 -124.610 ;
        RECT 311.385 -127.115 311.555 -125.395 ;
        RECT 312.365 -127.115 312.535 -125.395 ;
        RECT 314.430 -125.930 314.600 -125.390 ;
        RECT 315.410 -125.930 315.580 -125.390 ;
        RECT 313.840 -126.165 314.205 -126.100 ;
        RECT 313.340 -126.305 314.205 -126.165 ;
        RECT 313.230 -126.370 314.205 -126.305 ;
        RECT 313.230 -127.115 313.535 -126.370 ;
        RECT 313.840 -126.400 314.205 -126.370 ;
        RECT 316.390 -126.250 316.560 -125.390 ;
        RECT 311.385 -127.265 313.535 -127.115 ;
        RECT 311.385 -127.305 313.480 -127.265 ;
        RECT 314.430 -127.325 314.600 -126.545 ;
        RECT 314.920 -127.085 315.090 -126.545 ;
        RECT 315.410 -127.325 315.580 -126.545 ;
        RECT 315.900 -127.085 316.070 -126.545 ;
        RECT 316.390 -126.600 317.780 -126.250 ;
        RECT 309.605 -127.670 310.740 -127.660 ;
        RECT 312.795 -127.670 313.165 -127.540 ;
        RECT 309.605 -127.860 313.165 -127.670 ;
        RECT 313.730 -127.755 316.805 -127.325 ;
        RECT 310.735 -127.865 313.165 -127.860 ;
        RECT 310.735 -127.870 311.090 -127.865 ;
        RECT 312.795 -127.895 313.165 -127.865 ;
        RECT 310.895 -129.620 311.065 -128.080 ;
        RECT 311.385 -129.620 311.555 -128.080 ;
        RECT 311.875 -129.620 312.045 -128.080 ;
        RECT 312.365 -129.620 312.535 -128.080 ;
        RECT 312.855 -129.620 313.025 -128.080 ;
        RECT 311.380 -129.880 311.555 -129.620 ;
        RECT 314.950 -129.790 315.255 -127.755 ;
        RECT 317.400 -128.575 317.750 -126.600 ;
        RECT 318.620 -127.870 318.790 -124.950 ;
        RECT 319.655 -124.990 319.865 -124.780 ;
        RECT 318.600 -128.165 318.810 -127.870 ;
        RECT 319.675 -127.900 319.845 -124.990 ;
        RECT 320.165 -127.890 320.335 -124.950 ;
        RECT 320.645 -125.000 320.855 -124.780 ;
        RECT 319.660 -128.165 319.870 -127.900 ;
        RECT 318.600 -128.345 319.870 -128.165 ;
        RECT 320.145 -128.160 320.355 -127.890 ;
        RECT 320.655 -127.990 320.825 -125.000 ;
        RECT 321.715 -127.920 321.885 -124.950 ;
        RECT 320.145 -128.355 320.850 -128.160 ;
        RECT 320.635 -128.415 320.850 -128.355 ;
        RECT 319.425 -128.575 320.200 -128.525 ;
        RECT 317.400 -128.755 320.200 -128.575 ;
        RECT 317.400 -128.765 317.750 -128.755 ;
        RECT 319.425 -128.800 320.200 -128.755 ;
        RECT 320.635 -128.690 321.540 -128.415 ;
        RECT 320.635 -129.040 320.850 -128.690 ;
        RECT 318.075 -129.110 318.850 -129.065 ;
        RECT 317.890 -129.280 318.850 -129.110 ;
        RECT 318.075 -129.340 318.850 -129.280 ;
        RECT 319.080 -129.240 320.850 -129.040 ;
        RECT 321.710 -129.140 321.925 -127.920 ;
        RECT 322.895 -128.265 323.245 -121.580 ;
        RECT 324.235 -127.895 324.450 -118.020 ;
        RECT 325.870 -120.135 326.250 -116.615 ;
        RECT 327.380 -116.395 336.315 -116.205 ;
        RECT 327.380 -118.285 327.570 -116.395 ;
        RECT 333.415 -117.890 336.740 -117.750 ;
        RECT 333.415 -118.180 338.590 -117.890 ;
        RECT 327.265 -118.555 327.630 -118.285 ;
        RECT 333.415 -118.585 333.845 -118.180 ;
        RECT 334.715 -118.365 334.890 -118.180 ;
        RECT 336.340 -118.195 338.590 -118.180 ;
        RECT 329.155 -119.015 333.845 -118.585 ;
        RECT 328.395 -120.135 329.045 -120.005 ;
        RECT 325.870 -120.465 329.045 -120.135 ;
        RECT 329.855 -120.295 330.025 -119.015 ;
        RECT 330.345 -120.295 330.515 -119.255 ;
        RECT 330.835 -120.295 331.005 -119.015 ;
        RECT 331.325 -120.125 331.495 -119.255 ;
        RECT 334.230 -119.905 334.400 -118.365 ;
        RECT 334.720 -119.905 334.890 -118.365 ;
        RECT 335.210 -119.905 335.380 -118.365 ;
        RECT 335.700 -119.905 335.870 -118.365 ;
        RECT 336.190 -119.905 336.360 -118.365 ;
        RECT 334.070 -120.120 334.425 -120.115 ;
        RECT 336.130 -120.120 336.500 -120.090 ;
        RECT 334.070 -120.125 336.500 -120.120 ;
        RECT 331.325 -120.295 336.500 -120.125 ;
        RECT 338.285 -120.230 338.590 -118.195 ;
        RECT 331.330 -120.315 336.500 -120.295 ;
        RECT 331.330 -120.325 334.075 -120.315 ;
        RECT 329.265 -120.465 329.630 -120.435 ;
        RECT 336.130 -120.445 336.500 -120.315 ;
        RECT 325.870 -120.515 329.630 -120.465 ;
        RECT 328.395 -120.670 329.630 -120.515 ;
        RECT 333.805 -120.605 334.480 -120.565 ;
        RECT 333.705 -120.615 334.480 -120.605 ;
        RECT 328.395 -120.755 329.045 -120.670 ;
        RECT 329.265 -120.735 329.630 -120.670 ;
        RECT 328.530 -121.005 328.910 -120.755 ;
        RECT 332.670 -120.795 334.480 -120.615 ;
        RECT 337.065 -120.660 340.990 -120.230 ;
        RECT 333.705 -120.805 334.480 -120.795 ;
        RECT 333.805 -120.835 334.480 -120.805 ;
        RECT 334.720 -120.720 336.815 -120.680 ;
        RECT 334.720 -120.870 336.870 -120.720 ;
        RECT 329.855 -121.945 330.025 -120.905 ;
        RECT 330.835 -121.945 331.005 -120.905 ;
        RECT 331.815 -121.945 331.985 -120.905 ;
        RECT 334.720 -122.590 334.890 -120.870 ;
        RECT 335.700 -122.590 335.870 -120.870 ;
        RECT 336.565 -121.615 336.870 -120.870 ;
        RECT 337.765 -121.440 337.935 -120.660 ;
        RECT 338.255 -121.440 338.425 -120.900 ;
        RECT 338.745 -121.440 338.915 -120.660 ;
        RECT 339.235 -121.440 339.405 -120.900 ;
        RECT 337.175 -121.615 337.540 -121.585 ;
        RECT 336.565 -121.680 337.540 -121.615 ;
        RECT 336.675 -121.820 337.540 -121.680 ;
        RECT 337.175 -121.885 337.540 -121.820 ;
        RECT 339.725 -121.735 341.585 -121.385 ;
        RECT 337.765 -122.595 337.935 -122.055 ;
        RECT 338.745 -122.595 338.915 -122.055 ;
        RECT 339.725 -122.595 339.895 -121.735 ;
        RECT 337.995 -124.935 339.195 -124.765 ;
        RECT 329.725 -127.270 329.895 -125.550 ;
        RECT 330.705 -127.270 330.875 -125.550 ;
        RECT 332.770 -126.085 332.940 -125.545 ;
        RECT 333.750 -126.085 333.920 -125.545 ;
        RECT 332.180 -126.320 332.545 -126.255 ;
        RECT 331.680 -126.460 332.545 -126.320 ;
        RECT 331.570 -126.525 332.545 -126.460 ;
        RECT 331.570 -127.270 331.875 -126.525 ;
        RECT 332.180 -126.555 332.545 -126.525 ;
        RECT 334.730 -126.405 334.900 -125.545 ;
        RECT 329.725 -127.420 331.875 -127.270 ;
        RECT 329.725 -127.460 331.820 -127.420 ;
        RECT 332.770 -127.480 332.940 -126.700 ;
        RECT 333.260 -127.240 333.430 -126.700 ;
        RECT 333.750 -127.480 333.920 -126.700 ;
        RECT 334.240 -127.240 334.410 -126.700 ;
        RECT 334.730 -126.755 336.120 -126.405 ;
        RECT 327.945 -127.825 329.080 -127.815 ;
        RECT 331.135 -127.825 331.505 -127.695 ;
        RECT 324.235 -128.110 325.660 -127.895 ;
        RECT 327.945 -128.015 331.505 -127.825 ;
        RECT 332.070 -127.910 335.145 -127.480 ;
        RECT 329.075 -128.020 331.505 -128.015 ;
        RECT 329.075 -128.025 329.430 -128.020 ;
        RECT 331.135 -128.050 331.505 -128.020 ;
        RECT 322.840 -128.625 323.365 -128.265 ;
        RECT 325.445 -129.140 325.660 -128.110 ;
        RECT 313.005 -129.880 315.255 -129.790 ;
        RECT 310.795 -130.095 315.255 -129.880 ;
        RECT 310.795 -130.185 313.040 -130.095 ;
        RECT 314.950 -131.570 315.255 -130.095 ;
        RECT 318.620 -130.980 318.790 -129.510 ;
        RECT 319.080 -129.590 319.305 -129.240 ;
        RECT 321.040 -129.340 325.660 -129.140 ;
        RECT 321.280 -129.355 325.660 -129.340 ;
        RECT 318.585 -131.570 318.820 -130.980 ;
        RECT 319.110 -131.050 319.280 -129.590 ;
        RECT 319.600 -130.975 319.770 -129.510 ;
        RECT 320.810 -130.925 320.980 -129.510 ;
        RECT 321.280 -129.555 321.500 -129.355 ;
        RECT 319.565 -131.570 319.800 -130.975 ;
        RECT 320.775 -131.570 321.010 -130.925 ;
        RECT 321.300 -131.050 321.470 -129.555 ;
        RECT 329.235 -129.775 329.405 -128.235 ;
        RECT 329.725 -129.775 329.895 -128.235 ;
        RECT 330.215 -129.775 330.385 -128.235 ;
        RECT 330.705 -129.775 330.875 -128.235 ;
        RECT 331.195 -129.775 331.365 -128.235 ;
        RECT 329.720 -130.035 329.895 -129.775 ;
        RECT 333.290 -129.945 333.595 -127.910 ;
        RECT 335.740 -128.730 336.090 -126.755 ;
        RECT 336.960 -128.025 337.130 -125.105 ;
        RECT 337.995 -125.145 338.205 -124.935 ;
        RECT 336.940 -128.320 337.150 -128.025 ;
        RECT 338.015 -128.055 338.185 -125.145 ;
        RECT 338.505 -128.045 338.675 -125.105 ;
        RECT 338.985 -125.155 339.195 -124.935 ;
        RECT 338.000 -128.320 338.210 -128.055 ;
        RECT 336.940 -128.500 338.210 -128.320 ;
        RECT 338.485 -128.315 338.695 -128.045 ;
        RECT 338.995 -128.145 339.165 -125.155 ;
        RECT 340.055 -128.075 340.225 -125.105 ;
        RECT 338.485 -128.510 339.190 -128.315 ;
        RECT 338.975 -128.570 339.190 -128.510 ;
        RECT 337.765 -128.730 338.540 -128.680 ;
        RECT 335.740 -128.910 338.540 -128.730 ;
        RECT 335.740 -128.920 336.090 -128.910 ;
        RECT 337.765 -128.955 338.540 -128.910 ;
        RECT 338.975 -128.845 339.880 -128.570 ;
        RECT 338.975 -129.195 339.190 -128.845 ;
        RECT 336.415 -129.265 337.190 -129.220 ;
        RECT 336.230 -129.435 337.190 -129.265 ;
        RECT 336.415 -129.495 337.190 -129.435 ;
        RECT 337.420 -129.395 339.190 -129.195 ;
        RECT 340.050 -129.295 340.265 -128.075 ;
        RECT 341.235 -128.420 341.585 -121.735 ;
        RECT 341.180 -128.780 341.705 -128.420 ;
        RECT 343.525 -129.295 344.830 -128.490 ;
        RECT 331.345 -130.035 333.595 -129.945 ;
        RECT 329.135 -130.250 333.595 -130.035 ;
        RECT 329.135 -130.340 331.380 -130.250 ;
        RECT 314.950 -132.135 322.335 -131.570 ;
        RECT 333.290 -131.725 333.595 -130.250 ;
        RECT 336.960 -131.135 337.130 -129.665 ;
        RECT 337.420 -129.745 337.645 -129.395 ;
        RECT 339.380 -129.495 345.390 -129.295 ;
        RECT 339.620 -129.510 345.390 -129.495 ;
        RECT 336.925 -131.725 337.160 -131.135 ;
        RECT 337.450 -131.205 337.620 -129.745 ;
        RECT 337.940 -131.130 338.110 -129.665 ;
        RECT 339.150 -131.080 339.320 -129.665 ;
        RECT 339.620 -129.710 339.840 -129.510 ;
        RECT 337.905 -131.725 338.140 -131.130 ;
        RECT 339.115 -131.725 339.350 -131.080 ;
        RECT 339.640 -131.205 339.810 -129.710 ;
        RECT 343.525 -130.010 344.830 -129.510 ;
        RECT 333.290 -132.290 340.675 -131.725 ;
        RECT 350.275 -137.410 351.200 -110.370 ;
        RECT 355.410 -110.510 358.970 -110.320 ;
        RECT 359.535 -110.405 362.610 -109.975 ;
        RECT 355.465 -115.620 355.845 -110.510 ;
        RECT 356.540 -110.515 358.970 -110.510 ;
        RECT 356.540 -110.520 356.895 -110.515 ;
        RECT 358.600 -110.545 358.970 -110.515 ;
        RECT 356.700 -112.270 356.870 -110.730 ;
        RECT 357.190 -112.270 357.360 -110.730 ;
        RECT 357.680 -112.270 357.850 -110.730 ;
        RECT 358.170 -112.270 358.340 -110.730 ;
        RECT 358.660 -112.270 358.830 -110.730 ;
        RECT 357.185 -112.530 357.360 -112.270 ;
        RECT 360.755 -112.440 361.060 -110.405 ;
        RECT 363.205 -111.225 363.555 -109.250 ;
        RECT 364.425 -110.520 364.595 -107.600 ;
        RECT 365.460 -107.640 365.670 -107.430 ;
        RECT 364.405 -110.815 364.615 -110.520 ;
        RECT 365.480 -110.550 365.650 -107.640 ;
        RECT 365.970 -110.540 366.140 -107.600 ;
        RECT 366.450 -107.650 366.660 -107.430 ;
        RECT 365.465 -110.815 365.675 -110.550 ;
        RECT 364.405 -110.995 365.675 -110.815 ;
        RECT 365.950 -110.810 366.160 -110.540 ;
        RECT 366.460 -110.640 366.630 -107.650 ;
        RECT 367.520 -110.570 367.690 -107.600 ;
        RECT 365.950 -111.005 366.655 -110.810 ;
        RECT 366.440 -111.065 366.655 -111.005 ;
        RECT 365.230 -111.225 366.005 -111.175 ;
        RECT 363.205 -111.405 366.005 -111.225 ;
        RECT 363.205 -111.415 363.555 -111.405 ;
        RECT 365.230 -111.450 366.005 -111.405 ;
        RECT 366.440 -111.340 367.345 -111.065 ;
        RECT 366.440 -111.690 366.655 -111.340 ;
        RECT 363.880 -111.760 364.655 -111.715 ;
        RECT 363.695 -111.930 364.655 -111.760 ;
        RECT 363.880 -111.990 364.655 -111.930 ;
        RECT 364.885 -111.890 366.655 -111.690 ;
        RECT 367.515 -111.790 367.730 -110.570 ;
        RECT 368.700 -110.915 369.050 -104.230 ;
        RECT 404.140 -104.250 404.310 -103.210 ;
        RECT 405.120 -104.250 405.290 -103.210 ;
        RECT 406.100 -104.250 406.270 -103.210 ;
        RECT 409.005 -104.895 409.175 -103.175 ;
        RECT 409.985 -104.895 410.155 -103.175 ;
        RECT 410.850 -103.920 411.155 -103.175 ;
        RECT 412.050 -103.745 412.220 -102.965 ;
        RECT 412.540 -103.745 412.710 -103.205 ;
        RECT 413.030 -103.745 413.200 -102.965 ;
        RECT 413.520 -103.745 413.690 -103.205 ;
        RECT 411.460 -103.920 411.825 -103.890 ;
        RECT 410.850 -103.985 411.825 -103.920 ;
        RECT 410.960 -104.125 411.825 -103.985 ;
        RECT 411.460 -104.190 411.825 -104.125 ;
        RECT 414.010 -104.040 415.870 -103.690 ;
        RECT 412.050 -104.900 412.220 -104.360 ;
        RECT 413.030 -104.900 413.200 -104.360 ;
        RECT 414.010 -104.900 414.180 -104.040 ;
        RECT 375.280 -106.710 376.885 -106.540 ;
        RECT 374.385 -109.390 374.555 -106.890 ;
        RECT 374.380 -109.620 374.555 -109.390 ;
        RECT 375.280 -109.620 375.480 -106.710 ;
        RECT 375.725 -106.910 375.900 -106.710 ;
        RECT 375.730 -109.430 375.900 -106.910 ;
        RECT 376.220 -109.395 376.390 -106.890 ;
        RECT 376.710 -106.905 376.885 -106.710 ;
        RECT 374.380 -109.820 375.480 -109.620 ;
        RECT 376.205 -109.995 376.395 -109.395 ;
        RECT 376.710 -109.430 376.880 -106.905 ;
        RECT 377.360 -109.810 377.530 -106.890 ;
        RECT 378.990 -109.460 379.160 -106.890 ;
        RECT 380.130 -108.340 380.300 -106.890 ;
        RECT 412.280 -107.240 413.480 -107.070 ;
        RECT 380.125 -108.805 380.310 -108.340 ;
        RECT 380.125 -108.990 380.810 -108.805 ;
        RECT 378.990 -109.630 379.785 -109.460 ;
        RECT 378.105 -109.810 378.795 -109.755 ;
        RECT 374.385 -110.185 376.395 -109.995 ;
        RECT 376.730 -109.980 378.795 -109.810 ;
        RECT 373.200 -110.240 373.890 -110.190 ;
        RECT 371.250 -110.410 373.890 -110.240 ;
        RECT 368.645 -111.275 369.170 -110.915 ;
        RECT 371.250 -111.790 371.465 -110.410 ;
        RECT 373.200 -110.460 373.890 -110.410 ;
        RECT 373.480 -110.915 374.170 -110.870 ;
        RECT 372.430 -111.085 374.170 -110.915 ;
        RECT 372.430 -111.720 372.790 -111.085 ;
        RECT 373.480 -111.140 374.170 -111.085 ;
        RECT 372.430 -111.765 372.850 -111.720 ;
        RECT 358.810 -112.530 361.060 -112.440 ;
        RECT 356.600 -112.745 361.060 -112.530 ;
        RECT 356.600 -112.835 358.845 -112.745 ;
        RECT 360.755 -114.220 361.060 -112.745 ;
        RECT 364.425 -113.630 364.595 -112.160 ;
        RECT 364.885 -112.240 365.110 -111.890 ;
        RECT 366.845 -111.990 371.465 -111.790 ;
        RECT 367.085 -112.005 371.465 -111.990 ;
        RECT 364.390 -114.220 364.625 -113.630 ;
        RECT 364.915 -113.700 365.085 -112.240 ;
        RECT 365.405 -113.625 365.575 -112.160 ;
        RECT 366.615 -113.575 366.785 -112.160 ;
        RECT 367.085 -112.205 367.305 -112.005 ;
        RECT 372.455 -112.115 372.850 -111.765 ;
        RECT 365.370 -114.220 365.605 -113.625 ;
        RECT 366.580 -114.220 366.815 -113.575 ;
        RECT 367.105 -113.700 367.275 -112.205 ;
        RECT 373.895 -113.325 374.065 -111.870 ;
        RECT 373.885 -113.880 374.070 -113.325 ;
        RECT 374.385 -113.410 374.555 -110.185 ;
        RECT 375.530 -110.535 375.720 -110.185 ;
        RECT 376.730 -110.375 376.900 -109.980 ;
        RECT 378.105 -110.025 378.795 -109.980 ;
        RECT 375.480 -111.225 375.750 -110.535 ;
        RECT 376.245 -110.545 376.900 -110.375 ;
        RECT 377.230 -110.460 377.920 -110.190 ;
        RECT 379.155 -110.535 379.425 -109.845 ;
        RECT 379.615 -109.850 379.785 -109.630 ;
        RECT 379.615 -110.120 380.445 -109.850 ;
        RECT 376.245 -113.410 376.415 -110.545 ;
        RECT 379.615 -110.695 379.785 -110.120 ;
        RECT 380.045 -110.695 380.315 -110.610 ;
        RECT 376.735 -110.890 377.530 -110.715 ;
        RECT 379.615 -110.720 380.315 -110.695 ;
        RECT 379.475 -110.865 380.315 -110.720 ;
        RECT 376.735 -113.410 376.905 -110.890 ;
        RECT 377.360 -113.410 377.530 -110.890 ;
        RECT 377.850 -113.325 378.020 -110.870 ;
        RECT 378.500 -113.320 378.670 -110.870 ;
        RECT 371.200 -113.900 374.255 -113.880 ;
        RECT 377.845 -113.900 378.030 -113.325 ;
        RECT 378.485 -113.900 378.670 -113.320 ;
        RECT 378.990 -113.410 379.160 -110.870 ;
        RECT 379.475 -110.890 379.785 -110.865 ;
        RECT 379.480 -113.410 379.650 -110.890 ;
        RECT 380.045 -110.905 380.315 -110.865 ;
        RECT 380.620 -111.455 380.810 -108.990 ;
        RECT 394.860 -109.650 400.900 -108.735 ;
        RECT 404.010 -109.575 404.180 -107.855 ;
        RECT 404.990 -109.575 405.160 -107.855 ;
        RECT 407.055 -108.390 407.225 -107.850 ;
        RECT 408.035 -108.390 408.205 -107.850 ;
        RECT 406.465 -108.625 406.830 -108.560 ;
        RECT 405.965 -108.765 406.830 -108.625 ;
        RECT 405.855 -108.830 406.830 -108.765 ;
        RECT 405.855 -109.575 406.160 -108.830 ;
        RECT 406.465 -108.860 406.830 -108.830 ;
        RECT 409.015 -108.710 409.185 -107.850 ;
        RECT 403.095 -109.640 403.770 -109.610 ;
        RECT 402.995 -109.650 403.770 -109.640 ;
        RECT 394.860 -109.830 403.770 -109.650 ;
        RECT 404.010 -109.725 406.160 -109.575 ;
        RECT 404.010 -109.765 406.105 -109.725 ;
        RECT 407.055 -109.785 407.225 -109.005 ;
        RECT 407.545 -109.545 407.715 -109.005 ;
        RECT 408.035 -109.785 408.205 -109.005 ;
        RECT 408.525 -109.545 408.695 -109.005 ;
        RECT 409.015 -109.060 410.405 -108.710 ;
        RECT 394.860 -110.205 400.900 -109.830 ;
        RECT 402.995 -109.840 403.770 -109.830 ;
        RECT 403.095 -109.880 403.770 -109.840 ;
        RECT 402.230 -110.130 403.365 -110.120 ;
        RECT 405.420 -110.130 405.790 -110.000 ;
        RECT 380.620 -111.645 382.080 -111.455 ;
        RECT 380.130 -113.315 380.300 -111.870 ;
        RECT 380.620 -111.895 380.810 -111.645 ;
        RECT 380.120 -113.900 380.305 -113.315 ;
        RECT 380.620 -113.410 380.790 -111.895 ;
        RECT 371.200 -114.220 380.870 -113.900 ;
        RECT 360.755 -114.445 380.870 -114.220 ;
        RECT 360.755 -114.785 371.765 -114.445 ;
        RECT 373.505 -114.705 380.870 -114.445 ;
        RECT 352.090 -116.150 355.845 -115.620 ;
        RECT 381.890 -116.120 382.080 -111.645 ;
        RECT 352.090 -116.470 372.015 -116.150 ;
        RECT 352.090 -135.650 352.940 -116.470 ;
        RECT 355.465 -116.530 372.015 -116.470 ;
        RECT 355.465 -117.440 355.845 -116.530 ;
        RECT 355.465 -117.820 356.175 -117.440 ;
        RECT 355.795 -119.765 356.175 -117.820 ;
        RECT 360.840 -117.650 364.165 -117.510 ;
        RECT 360.840 -117.940 366.015 -117.650 ;
        RECT 369.885 -117.935 370.345 -117.510 ;
        RECT 360.840 -118.345 361.270 -117.940 ;
        RECT 362.140 -118.125 362.315 -117.940 ;
        RECT 363.765 -117.955 366.015 -117.940 ;
        RECT 356.580 -118.775 361.270 -118.345 ;
        RECT 355.795 -120.225 356.470 -119.765 ;
        RECT 357.280 -120.055 357.450 -118.775 ;
        RECT 357.770 -120.055 357.940 -119.015 ;
        RECT 358.260 -120.055 358.430 -118.775 ;
        RECT 358.750 -119.885 358.920 -119.015 ;
        RECT 361.655 -119.665 361.825 -118.125 ;
        RECT 362.145 -119.665 362.315 -118.125 ;
        RECT 362.635 -119.665 362.805 -118.125 ;
        RECT 363.125 -119.665 363.295 -118.125 ;
        RECT 363.615 -119.665 363.785 -118.125 ;
        RECT 361.495 -119.880 361.850 -119.875 ;
        RECT 363.555 -119.880 363.925 -119.850 ;
        RECT 361.495 -119.885 363.925 -119.880 ;
        RECT 358.750 -120.055 363.925 -119.885 ;
        RECT 365.710 -119.990 366.015 -117.955 ;
        RECT 358.755 -120.075 363.925 -120.055 ;
        RECT 358.755 -120.085 361.500 -120.075 ;
        RECT 356.690 -120.225 357.055 -120.195 ;
        RECT 363.555 -120.205 363.925 -120.075 ;
        RECT 355.795 -120.310 357.055 -120.225 ;
        RECT 355.820 -120.430 357.055 -120.310 ;
        RECT 361.230 -120.365 361.905 -120.325 ;
        RECT 361.130 -120.375 361.905 -120.365 ;
        RECT 355.820 -120.515 356.470 -120.430 ;
        RECT 356.690 -120.495 357.055 -120.430 ;
        RECT 360.095 -120.555 361.905 -120.375 ;
        RECT 364.490 -120.420 368.415 -119.990 ;
        RECT 361.130 -120.565 361.905 -120.555 ;
        RECT 361.230 -120.595 361.905 -120.565 ;
        RECT 362.145 -120.480 364.240 -120.440 ;
        RECT 362.145 -120.630 364.295 -120.480 ;
        RECT 357.280 -121.705 357.450 -120.665 ;
        RECT 358.260 -121.705 358.430 -120.665 ;
        RECT 359.240 -121.705 359.410 -120.665 ;
        RECT 362.145 -122.350 362.315 -120.630 ;
        RECT 363.125 -122.350 363.295 -120.630 ;
        RECT 363.990 -121.375 364.295 -120.630 ;
        RECT 365.190 -121.200 365.360 -120.420 ;
        RECT 365.680 -121.200 365.850 -120.660 ;
        RECT 366.170 -121.200 366.340 -120.420 ;
        RECT 366.660 -121.200 366.830 -120.660 ;
        RECT 364.600 -121.375 364.965 -121.345 ;
        RECT 363.990 -121.440 364.965 -121.375 ;
        RECT 364.100 -121.580 364.965 -121.440 ;
        RECT 364.600 -121.645 364.965 -121.580 ;
        RECT 367.150 -121.495 369.010 -121.145 ;
        RECT 365.190 -122.355 365.360 -121.815 ;
        RECT 366.170 -122.355 366.340 -121.815 ;
        RECT 367.150 -122.355 367.320 -121.495 ;
        RECT 365.420 -124.695 366.620 -124.525 ;
        RECT 357.150 -127.030 357.320 -125.310 ;
        RECT 358.130 -127.030 358.300 -125.310 ;
        RECT 360.195 -125.845 360.365 -125.305 ;
        RECT 361.175 -125.845 361.345 -125.305 ;
        RECT 359.605 -126.080 359.970 -126.015 ;
        RECT 359.105 -126.220 359.970 -126.080 ;
        RECT 358.995 -126.285 359.970 -126.220 ;
        RECT 358.995 -127.030 359.300 -126.285 ;
        RECT 359.605 -126.315 359.970 -126.285 ;
        RECT 362.155 -126.165 362.325 -125.305 ;
        RECT 357.150 -127.180 359.300 -127.030 ;
        RECT 357.150 -127.220 359.245 -127.180 ;
        RECT 360.195 -127.240 360.365 -126.460 ;
        RECT 360.685 -127.000 360.855 -126.460 ;
        RECT 361.175 -127.240 361.345 -126.460 ;
        RECT 361.665 -127.000 361.835 -126.460 ;
        RECT 362.155 -126.515 363.545 -126.165 ;
        RECT 355.370 -127.585 356.505 -127.575 ;
        RECT 358.560 -127.585 358.930 -127.455 ;
        RECT 355.370 -127.775 358.930 -127.585 ;
        RECT 359.495 -127.670 362.570 -127.240 ;
        RECT 356.500 -127.780 358.930 -127.775 ;
        RECT 356.500 -127.785 356.855 -127.780 ;
        RECT 358.560 -127.810 358.930 -127.780 ;
        RECT 356.660 -129.535 356.830 -127.995 ;
        RECT 357.150 -129.535 357.320 -127.995 ;
        RECT 357.640 -129.535 357.810 -127.995 ;
        RECT 358.130 -129.535 358.300 -127.995 ;
        RECT 358.620 -129.535 358.790 -127.995 ;
        RECT 357.145 -129.795 357.320 -129.535 ;
        RECT 360.715 -129.705 361.020 -127.670 ;
        RECT 363.165 -128.490 363.515 -126.515 ;
        RECT 364.385 -127.785 364.555 -124.865 ;
        RECT 365.420 -124.905 365.630 -124.695 ;
        RECT 364.365 -128.080 364.575 -127.785 ;
        RECT 365.440 -127.815 365.610 -124.905 ;
        RECT 365.930 -127.805 366.100 -124.865 ;
        RECT 366.410 -124.915 366.620 -124.695 ;
        RECT 365.425 -128.080 365.635 -127.815 ;
        RECT 364.365 -128.260 365.635 -128.080 ;
        RECT 365.910 -128.075 366.120 -127.805 ;
        RECT 366.420 -127.905 366.590 -124.915 ;
        RECT 367.480 -127.835 367.650 -124.865 ;
        RECT 365.910 -128.270 366.615 -128.075 ;
        RECT 366.400 -128.330 366.615 -128.270 ;
        RECT 365.190 -128.490 365.965 -128.440 ;
        RECT 363.165 -128.670 365.965 -128.490 ;
        RECT 363.165 -128.680 363.515 -128.670 ;
        RECT 365.190 -128.715 365.965 -128.670 ;
        RECT 366.400 -128.605 367.305 -128.330 ;
        RECT 366.400 -128.955 366.615 -128.605 ;
        RECT 363.840 -129.025 364.615 -128.980 ;
        RECT 363.655 -129.195 364.615 -129.025 ;
        RECT 363.840 -129.255 364.615 -129.195 ;
        RECT 364.845 -129.155 366.615 -128.955 ;
        RECT 367.475 -129.055 367.690 -127.835 ;
        RECT 368.660 -128.180 369.010 -121.495 ;
        RECT 370.000 -127.810 370.215 -117.935 ;
        RECT 371.635 -120.050 372.015 -116.530 ;
        RECT 373.145 -116.310 382.080 -116.120 ;
        RECT 373.145 -118.200 373.335 -116.310 ;
        RECT 379.180 -117.805 382.505 -117.665 ;
        RECT 379.180 -118.095 384.355 -117.805 ;
        RECT 373.030 -118.470 373.395 -118.200 ;
        RECT 379.180 -118.500 379.610 -118.095 ;
        RECT 380.480 -118.280 380.655 -118.095 ;
        RECT 382.105 -118.110 384.355 -118.095 ;
        RECT 374.920 -118.930 379.610 -118.500 ;
        RECT 374.160 -120.050 374.810 -119.920 ;
        RECT 371.635 -120.380 374.810 -120.050 ;
        RECT 375.620 -120.210 375.790 -118.930 ;
        RECT 376.110 -120.210 376.280 -119.170 ;
        RECT 376.600 -120.210 376.770 -118.930 ;
        RECT 377.090 -120.040 377.260 -119.170 ;
        RECT 379.995 -119.820 380.165 -118.280 ;
        RECT 380.485 -119.820 380.655 -118.280 ;
        RECT 380.975 -119.820 381.145 -118.280 ;
        RECT 381.465 -119.820 381.635 -118.280 ;
        RECT 381.955 -119.820 382.125 -118.280 ;
        RECT 379.835 -120.035 380.190 -120.030 ;
        RECT 381.895 -120.035 382.265 -120.005 ;
        RECT 379.835 -120.040 382.265 -120.035 ;
        RECT 377.090 -120.210 382.265 -120.040 ;
        RECT 384.050 -120.145 384.355 -118.110 ;
        RECT 377.095 -120.230 382.265 -120.210 ;
        RECT 377.095 -120.240 379.840 -120.230 ;
        RECT 375.030 -120.380 375.395 -120.350 ;
        RECT 381.895 -120.360 382.265 -120.230 ;
        RECT 371.635 -120.430 375.395 -120.380 ;
        RECT 374.160 -120.585 375.395 -120.430 ;
        RECT 379.570 -120.520 380.245 -120.480 ;
        RECT 379.470 -120.530 380.245 -120.520 ;
        RECT 374.160 -120.670 374.810 -120.585 ;
        RECT 375.030 -120.650 375.395 -120.585 ;
        RECT 374.295 -120.920 374.675 -120.670 ;
        RECT 378.435 -120.710 380.245 -120.530 ;
        RECT 382.830 -120.575 386.755 -120.145 ;
        RECT 379.470 -120.720 380.245 -120.710 ;
        RECT 379.570 -120.750 380.245 -120.720 ;
        RECT 380.485 -120.635 382.580 -120.595 ;
        RECT 380.485 -120.785 382.635 -120.635 ;
        RECT 375.620 -121.860 375.790 -120.820 ;
        RECT 376.600 -121.860 376.770 -120.820 ;
        RECT 377.580 -121.860 377.750 -120.820 ;
        RECT 380.485 -122.505 380.655 -120.785 ;
        RECT 381.465 -122.505 381.635 -120.785 ;
        RECT 382.330 -121.530 382.635 -120.785 ;
        RECT 383.530 -121.355 383.700 -120.575 ;
        RECT 384.020 -121.355 384.190 -120.815 ;
        RECT 384.510 -121.355 384.680 -120.575 ;
        RECT 385.000 -121.355 385.170 -120.815 ;
        RECT 382.940 -121.530 383.305 -121.500 ;
        RECT 382.330 -121.595 383.305 -121.530 ;
        RECT 382.440 -121.735 383.305 -121.595 ;
        RECT 382.940 -121.800 383.305 -121.735 ;
        RECT 385.490 -121.650 387.350 -121.300 ;
        RECT 383.530 -122.510 383.700 -121.970 ;
        RECT 384.510 -122.510 384.680 -121.970 ;
        RECT 385.490 -122.510 385.660 -121.650 ;
        RECT 383.760 -124.850 384.960 -124.680 ;
        RECT 375.490 -127.185 375.660 -125.465 ;
        RECT 376.470 -127.185 376.640 -125.465 ;
        RECT 378.535 -126.000 378.705 -125.460 ;
        RECT 379.515 -126.000 379.685 -125.460 ;
        RECT 377.945 -126.235 378.310 -126.170 ;
        RECT 377.445 -126.375 378.310 -126.235 ;
        RECT 377.335 -126.440 378.310 -126.375 ;
        RECT 377.335 -127.185 377.640 -126.440 ;
        RECT 377.945 -126.470 378.310 -126.440 ;
        RECT 380.495 -126.320 380.665 -125.460 ;
        RECT 375.490 -127.335 377.640 -127.185 ;
        RECT 375.490 -127.375 377.585 -127.335 ;
        RECT 378.535 -127.395 378.705 -126.615 ;
        RECT 379.025 -127.155 379.195 -126.615 ;
        RECT 379.515 -127.395 379.685 -126.615 ;
        RECT 380.005 -127.155 380.175 -126.615 ;
        RECT 380.495 -126.670 381.885 -126.320 ;
        RECT 373.710 -127.740 374.845 -127.730 ;
        RECT 376.900 -127.740 377.270 -127.610 ;
        RECT 370.000 -128.025 371.425 -127.810 ;
        RECT 373.710 -127.930 377.270 -127.740 ;
        RECT 377.835 -127.825 380.910 -127.395 ;
        RECT 374.840 -127.935 377.270 -127.930 ;
        RECT 374.840 -127.940 375.195 -127.935 ;
        RECT 376.900 -127.965 377.270 -127.935 ;
        RECT 368.605 -128.540 369.130 -128.180 ;
        RECT 371.210 -129.055 371.425 -128.025 ;
        RECT 358.770 -129.795 361.020 -129.705 ;
        RECT 356.560 -130.010 361.020 -129.795 ;
        RECT 356.560 -130.100 358.805 -130.010 ;
        RECT 360.715 -131.485 361.020 -130.010 ;
        RECT 364.385 -130.895 364.555 -129.425 ;
        RECT 364.845 -129.505 365.070 -129.155 ;
        RECT 366.805 -129.255 371.425 -129.055 ;
        RECT 367.045 -129.270 371.425 -129.255 ;
        RECT 364.350 -131.485 364.585 -130.895 ;
        RECT 364.875 -130.965 365.045 -129.505 ;
        RECT 365.365 -130.890 365.535 -129.425 ;
        RECT 366.575 -130.840 366.745 -129.425 ;
        RECT 367.045 -129.470 367.265 -129.270 ;
        RECT 365.330 -131.485 365.565 -130.890 ;
        RECT 366.540 -131.485 366.775 -130.840 ;
        RECT 367.065 -130.965 367.235 -129.470 ;
        RECT 375.000 -129.690 375.170 -128.150 ;
        RECT 375.490 -129.690 375.660 -128.150 ;
        RECT 375.980 -129.690 376.150 -128.150 ;
        RECT 376.470 -129.690 376.640 -128.150 ;
        RECT 376.960 -129.690 377.130 -128.150 ;
        RECT 375.485 -129.950 375.660 -129.690 ;
        RECT 379.055 -129.860 379.360 -127.825 ;
        RECT 381.505 -128.645 381.855 -126.670 ;
        RECT 382.725 -127.940 382.895 -125.020 ;
        RECT 383.760 -125.060 383.970 -124.850 ;
        RECT 382.705 -128.235 382.915 -127.940 ;
        RECT 383.780 -127.970 383.950 -125.060 ;
        RECT 384.270 -127.960 384.440 -125.020 ;
        RECT 384.750 -125.070 384.960 -124.850 ;
        RECT 383.765 -128.235 383.975 -127.970 ;
        RECT 382.705 -128.415 383.975 -128.235 ;
        RECT 384.250 -128.230 384.460 -127.960 ;
        RECT 384.760 -128.060 384.930 -125.070 ;
        RECT 385.820 -127.990 385.990 -125.020 ;
        RECT 384.250 -128.425 384.955 -128.230 ;
        RECT 384.740 -128.485 384.955 -128.425 ;
        RECT 383.530 -128.645 384.305 -128.595 ;
        RECT 381.505 -128.825 384.305 -128.645 ;
        RECT 381.505 -128.835 381.855 -128.825 ;
        RECT 383.530 -128.870 384.305 -128.825 ;
        RECT 384.740 -128.760 385.645 -128.485 ;
        RECT 384.740 -129.110 384.955 -128.760 ;
        RECT 382.180 -129.180 382.955 -129.135 ;
        RECT 381.995 -129.350 382.955 -129.180 ;
        RECT 382.180 -129.410 382.955 -129.350 ;
        RECT 383.185 -129.310 384.955 -129.110 ;
        RECT 385.815 -129.210 386.030 -127.990 ;
        RECT 387.000 -128.335 387.350 -121.650 ;
        RECT 386.945 -128.695 387.470 -128.335 ;
        RECT 389.955 -129.210 390.465 -129.020 ;
        RECT 377.110 -129.950 379.360 -129.860 ;
        RECT 374.900 -130.165 379.360 -129.950 ;
        RECT 374.900 -130.255 377.145 -130.165 ;
        RECT 360.715 -132.050 368.100 -131.485 ;
        RECT 379.055 -131.640 379.360 -130.165 ;
        RECT 382.725 -131.050 382.895 -129.580 ;
        RECT 383.185 -129.660 383.410 -129.310 ;
        RECT 385.145 -129.410 391.155 -129.210 ;
        RECT 385.385 -129.425 391.155 -129.410 ;
        RECT 382.690 -131.640 382.925 -131.050 ;
        RECT 383.215 -131.120 383.385 -129.660 ;
        RECT 383.705 -131.045 383.875 -129.580 ;
        RECT 384.915 -130.995 385.085 -129.580 ;
        RECT 385.385 -129.625 385.605 -129.425 ;
        RECT 389.955 -129.575 390.465 -129.425 ;
        RECT 383.670 -131.640 383.905 -131.045 ;
        RECT 384.880 -131.640 385.115 -130.995 ;
        RECT 385.405 -131.120 385.575 -129.625 ;
        RECT 379.055 -132.205 386.440 -131.640 ;
        RECT 351.895 -136.550 353.125 -135.650 ;
        RECT 349.850 -138.635 351.760 -137.410 ;
        RECT 394.860 -137.425 396.330 -110.205 ;
        RECT 402.230 -110.320 405.790 -110.130 ;
        RECT 406.355 -110.215 409.430 -109.785 ;
        RECT 402.285 -115.225 402.665 -110.320 ;
        RECT 403.360 -110.325 405.790 -110.320 ;
        RECT 403.360 -110.330 403.715 -110.325 ;
        RECT 405.420 -110.355 405.790 -110.325 ;
        RECT 403.520 -112.080 403.690 -110.540 ;
        RECT 404.010 -112.080 404.180 -110.540 ;
        RECT 404.500 -112.080 404.670 -110.540 ;
        RECT 404.990 -112.080 405.160 -110.540 ;
        RECT 405.480 -112.080 405.650 -110.540 ;
        RECT 404.005 -112.340 404.180 -112.080 ;
        RECT 407.575 -112.250 407.880 -110.215 ;
        RECT 410.025 -111.035 410.375 -109.060 ;
        RECT 411.245 -110.330 411.415 -107.410 ;
        RECT 412.280 -107.450 412.490 -107.240 ;
        RECT 411.225 -110.625 411.435 -110.330 ;
        RECT 412.300 -110.360 412.470 -107.450 ;
        RECT 412.790 -110.350 412.960 -107.410 ;
        RECT 413.270 -107.460 413.480 -107.240 ;
        RECT 412.285 -110.625 412.495 -110.360 ;
        RECT 411.225 -110.805 412.495 -110.625 ;
        RECT 412.770 -110.620 412.980 -110.350 ;
        RECT 413.280 -110.450 413.450 -107.460 ;
        RECT 414.340 -110.380 414.510 -107.410 ;
        RECT 412.770 -110.815 413.475 -110.620 ;
        RECT 413.260 -110.875 413.475 -110.815 ;
        RECT 412.050 -111.035 412.825 -110.985 ;
        RECT 410.025 -111.215 412.825 -111.035 ;
        RECT 410.025 -111.225 410.375 -111.215 ;
        RECT 412.050 -111.260 412.825 -111.215 ;
        RECT 413.260 -111.150 414.165 -110.875 ;
        RECT 413.260 -111.500 413.475 -111.150 ;
        RECT 410.700 -111.570 411.475 -111.525 ;
        RECT 410.515 -111.740 411.475 -111.570 ;
        RECT 410.700 -111.800 411.475 -111.740 ;
        RECT 411.705 -111.700 413.475 -111.500 ;
        RECT 414.335 -111.600 414.550 -110.380 ;
        RECT 415.520 -110.725 415.870 -104.040 ;
        RECT 422.100 -106.520 423.705 -106.350 ;
        RECT 421.205 -109.200 421.375 -106.700 ;
        RECT 421.200 -109.430 421.375 -109.200 ;
        RECT 422.100 -109.430 422.300 -106.520 ;
        RECT 422.545 -106.720 422.720 -106.520 ;
        RECT 422.550 -109.240 422.720 -106.720 ;
        RECT 423.040 -109.205 423.210 -106.700 ;
        RECT 423.530 -106.715 423.705 -106.520 ;
        RECT 421.200 -109.630 422.300 -109.430 ;
        RECT 423.025 -109.805 423.215 -109.205 ;
        RECT 423.530 -109.240 423.700 -106.715 ;
        RECT 424.180 -109.620 424.350 -106.700 ;
        RECT 425.810 -109.270 425.980 -106.700 ;
        RECT 426.950 -108.150 427.120 -106.700 ;
        RECT 426.945 -108.615 427.130 -108.150 ;
        RECT 426.945 -108.800 427.630 -108.615 ;
        RECT 425.810 -109.440 426.605 -109.270 ;
        RECT 424.925 -109.620 425.615 -109.565 ;
        RECT 421.205 -109.995 423.215 -109.805 ;
        RECT 423.550 -109.790 425.615 -109.620 ;
        RECT 420.020 -110.050 420.710 -110.000 ;
        RECT 418.070 -110.220 420.710 -110.050 ;
        RECT 415.465 -111.085 415.990 -110.725 ;
        RECT 418.070 -111.600 418.285 -110.220 ;
        RECT 420.020 -110.270 420.710 -110.220 ;
        RECT 420.300 -110.725 420.990 -110.680 ;
        RECT 419.250 -110.895 420.990 -110.725 ;
        RECT 419.250 -111.530 419.610 -110.895 ;
        RECT 420.300 -110.950 420.990 -110.895 ;
        RECT 419.250 -111.575 419.670 -111.530 ;
        RECT 405.630 -112.340 407.880 -112.250 ;
        RECT 403.420 -112.555 407.880 -112.340 ;
        RECT 403.420 -112.645 405.665 -112.555 ;
        RECT 407.575 -114.030 407.880 -112.555 ;
        RECT 411.245 -113.440 411.415 -111.970 ;
        RECT 411.705 -112.050 411.930 -111.700 ;
        RECT 413.665 -111.800 418.285 -111.600 ;
        RECT 413.905 -111.815 418.285 -111.800 ;
        RECT 411.210 -114.030 411.445 -113.440 ;
        RECT 411.735 -113.510 411.905 -112.050 ;
        RECT 412.225 -113.435 412.395 -111.970 ;
        RECT 413.435 -113.385 413.605 -111.970 ;
        RECT 413.905 -112.015 414.125 -111.815 ;
        RECT 419.275 -111.925 419.670 -111.575 ;
        RECT 412.190 -114.030 412.425 -113.435 ;
        RECT 413.400 -114.030 413.635 -113.385 ;
        RECT 413.925 -113.510 414.095 -112.015 ;
        RECT 420.715 -113.135 420.885 -111.680 ;
        RECT 420.705 -113.690 420.890 -113.135 ;
        RECT 421.205 -113.220 421.375 -109.995 ;
        RECT 422.350 -110.345 422.540 -109.995 ;
        RECT 423.550 -110.185 423.720 -109.790 ;
        RECT 424.925 -109.835 425.615 -109.790 ;
        RECT 422.300 -111.035 422.570 -110.345 ;
        RECT 423.065 -110.355 423.720 -110.185 ;
        RECT 424.050 -110.270 424.740 -110.000 ;
        RECT 425.975 -110.345 426.245 -109.655 ;
        RECT 426.435 -109.660 426.605 -109.440 ;
        RECT 426.435 -109.930 427.265 -109.660 ;
        RECT 423.065 -113.220 423.235 -110.355 ;
        RECT 426.435 -110.505 426.605 -109.930 ;
        RECT 426.865 -110.505 427.135 -110.420 ;
        RECT 423.555 -110.700 424.350 -110.525 ;
        RECT 426.435 -110.530 427.135 -110.505 ;
        RECT 426.295 -110.675 427.135 -110.530 ;
        RECT 423.555 -113.220 423.725 -110.700 ;
        RECT 424.180 -113.220 424.350 -110.700 ;
        RECT 424.670 -113.135 424.840 -110.680 ;
        RECT 425.320 -113.130 425.490 -110.680 ;
        RECT 418.020 -113.710 421.075 -113.690 ;
        RECT 424.665 -113.710 424.850 -113.135 ;
        RECT 425.305 -113.710 425.490 -113.130 ;
        RECT 425.810 -113.220 425.980 -110.680 ;
        RECT 426.295 -110.700 426.605 -110.675 ;
        RECT 426.300 -113.220 426.470 -110.700 ;
        RECT 426.865 -110.715 427.135 -110.675 ;
        RECT 427.440 -111.265 427.630 -108.800 ;
        RECT 427.440 -111.455 428.900 -111.265 ;
        RECT 426.950 -113.125 427.120 -111.680 ;
        RECT 427.440 -111.705 427.630 -111.455 ;
        RECT 426.940 -113.710 427.125 -113.125 ;
        RECT 427.440 -113.220 427.610 -111.705 ;
        RECT 418.020 -114.030 427.690 -113.710 ;
        RECT 407.575 -114.255 427.690 -114.030 ;
        RECT 407.575 -114.595 418.585 -114.255 ;
        RECT 420.325 -114.515 427.690 -114.255 ;
        RECT 398.470 -115.960 402.875 -115.225 ;
        RECT 428.710 -115.930 428.900 -111.455 ;
        RECT 398.470 -116.340 418.835 -115.960 ;
        RECT 398.470 -116.355 402.875 -116.340 ;
        RECT 394.615 -138.615 396.615 -137.425 ;
        RECT 208.055 -140.645 209.255 -140.600 ;
        RECT 305.850 -140.765 307.570 -139.350 ;
        RECT 398.470 -139.365 399.600 -116.355 ;
        RECT 402.285 -117.250 402.665 -116.355 ;
        RECT 402.285 -117.630 402.995 -117.250 ;
        RECT 402.615 -119.575 402.995 -117.630 ;
        RECT 407.660 -117.460 410.985 -117.320 ;
        RECT 407.660 -117.750 412.835 -117.460 ;
        RECT 416.705 -117.745 417.165 -117.320 ;
        RECT 407.660 -118.155 408.090 -117.750 ;
        RECT 408.960 -117.935 409.135 -117.750 ;
        RECT 410.585 -117.765 412.835 -117.750 ;
        RECT 403.400 -118.585 408.090 -118.155 ;
        RECT 402.615 -120.035 403.290 -119.575 ;
        RECT 404.100 -119.865 404.270 -118.585 ;
        RECT 404.590 -119.865 404.760 -118.825 ;
        RECT 405.080 -119.865 405.250 -118.585 ;
        RECT 405.570 -119.695 405.740 -118.825 ;
        RECT 408.475 -119.475 408.645 -117.935 ;
        RECT 408.965 -119.475 409.135 -117.935 ;
        RECT 409.455 -119.475 409.625 -117.935 ;
        RECT 409.945 -119.475 410.115 -117.935 ;
        RECT 410.435 -119.475 410.605 -117.935 ;
        RECT 408.315 -119.690 408.670 -119.685 ;
        RECT 410.375 -119.690 410.745 -119.660 ;
        RECT 408.315 -119.695 410.745 -119.690 ;
        RECT 405.570 -119.865 410.745 -119.695 ;
        RECT 412.530 -119.800 412.835 -117.765 ;
        RECT 405.575 -119.885 410.745 -119.865 ;
        RECT 405.575 -119.895 408.320 -119.885 ;
        RECT 403.510 -120.035 403.875 -120.005 ;
        RECT 410.375 -120.015 410.745 -119.885 ;
        RECT 402.615 -120.120 403.875 -120.035 ;
        RECT 402.640 -120.240 403.875 -120.120 ;
        RECT 408.050 -120.175 408.725 -120.135 ;
        RECT 407.950 -120.185 408.725 -120.175 ;
        RECT 402.640 -120.325 403.290 -120.240 ;
        RECT 403.510 -120.305 403.875 -120.240 ;
        RECT 406.915 -120.365 408.725 -120.185 ;
        RECT 411.310 -120.230 415.235 -119.800 ;
        RECT 407.950 -120.375 408.725 -120.365 ;
        RECT 408.050 -120.405 408.725 -120.375 ;
        RECT 408.965 -120.290 411.060 -120.250 ;
        RECT 408.965 -120.440 411.115 -120.290 ;
        RECT 404.100 -121.515 404.270 -120.475 ;
        RECT 405.080 -121.515 405.250 -120.475 ;
        RECT 406.060 -121.515 406.230 -120.475 ;
        RECT 408.965 -122.160 409.135 -120.440 ;
        RECT 409.945 -122.160 410.115 -120.440 ;
        RECT 410.810 -121.185 411.115 -120.440 ;
        RECT 412.010 -121.010 412.180 -120.230 ;
        RECT 412.500 -121.010 412.670 -120.470 ;
        RECT 412.990 -121.010 413.160 -120.230 ;
        RECT 413.480 -121.010 413.650 -120.470 ;
        RECT 411.420 -121.185 411.785 -121.155 ;
        RECT 410.810 -121.250 411.785 -121.185 ;
        RECT 410.920 -121.390 411.785 -121.250 ;
        RECT 411.420 -121.455 411.785 -121.390 ;
        RECT 413.970 -121.305 415.830 -120.955 ;
        RECT 412.010 -122.165 412.180 -121.625 ;
        RECT 412.990 -122.165 413.160 -121.625 ;
        RECT 413.970 -122.165 414.140 -121.305 ;
        RECT 412.240 -124.505 413.440 -124.335 ;
        RECT 403.970 -126.840 404.140 -125.120 ;
        RECT 404.950 -126.840 405.120 -125.120 ;
        RECT 407.015 -125.655 407.185 -125.115 ;
        RECT 407.995 -125.655 408.165 -125.115 ;
        RECT 406.425 -125.890 406.790 -125.825 ;
        RECT 405.925 -126.030 406.790 -125.890 ;
        RECT 405.815 -126.095 406.790 -126.030 ;
        RECT 405.815 -126.840 406.120 -126.095 ;
        RECT 406.425 -126.125 406.790 -126.095 ;
        RECT 408.975 -125.975 409.145 -125.115 ;
        RECT 403.970 -126.990 406.120 -126.840 ;
        RECT 403.970 -127.030 406.065 -126.990 ;
        RECT 407.015 -127.050 407.185 -126.270 ;
        RECT 407.505 -126.810 407.675 -126.270 ;
        RECT 407.995 -127.050 408.165 -126.270 ;
        RECT 408.485 -126.810 408.655 -126.270 ;
        RECT 408.975 -126.325 410.365 -125.975 ;
        RECT 402.190 -127.395 403.325 -127.385 ;
        RECT 405.380 -127.395 405.750 -127.265 ;
        RECT 402.190 -127.585 405.750 -127.395 ;
        RECT 406.315 -127.480 409.390 -127.050 ;
        RECT 403.320 -127.590 405.750 -127.585 ;
        RECT 403.320 -127.595 403.675 -127.590 ;
        RECT 405.380 -127.620 405.750 -127.590 ;
        RECT 403.480 -129.345 403.650 -127.805 ;
        RECT 403.970 -129.345 404.140 -127.805 ;
        RECT 404.460 -129.345 404.630 -127.805 ;
        RECT 404.950 -129.345 405.120 -127.805 ;
        RECT 405.440 -129.345 405.610 -127.805 ;
        RECT 403.965 -129.605 404.140 -129.345 ;
        RECT 407.535 -129.515 407.840 -127.480 ;
        RECT 409.985 -128.300 410.335 -126.325 ;
        RECT 411.205 -127.595 411.375 -124.675 ;
        RECT 412.240 -124.715 412.450 -124.505 ;
        RECT 411.185 -127.890 411.395 -127.595 ;
        RECT 412.260 -127.625 412.430 -124.715 ;
        RECT 412.750 -127.615 412.920 -124.675 ;
        RECT 413.230 -124.725 413.440 -124.505 ;
        RECT 412.245 -127.890 412.455 -127.625 ;
        RECT 411.185 -128.070 412.455 -127.890 ;
        RECT 412.730 -127.885 412.940 -127.615 ;
        RECT 413.240 -127.715 413.410 -124.725 ;
        RECT 414.300 -127.645 414.470 -124.675 ;
        RECT 412.730 -128.080 413.435 -127.885 ;
        RECT 413.220 -128.140 413.435 -128.080 ;
        RECT 412.010 -128.300 412.785 -128.250 ;
        RECT 409.985 -128.480 412.785 -128.300 ;
        RECT 409.985 -128.490 410.335 -128.480 ;
        RECT 412.010 -128.525 412.785 -128.480 ;
        RECT 413.220 -128.415 414.125 -128.140 ;
        RECT 413.220 -128.765 413.435 -128.415 ;
        RECT 410.660 -128.835 411.435 -128.790 ;
        RECT 410.475 -129.005 411.435 -128.835 ;
        RECT 410.660 -129.065 411.435 -129.005 ;
        RECT 411.665 -128.965 413.435 -128.765 ;
        RECT 414.295 -128.865 414.510 -127.645 ;
        RECT 415.480 -127.990 415.830 -121.305 ;
        RECT 416.820 -127.620 417.035 -117.745 ;
        RECT 418.455 -119.860 418.835 -116.340 ;
        RECT 419.965 -116.120 428.900 -115.930 ;
        RECT 419.965 -118.010 420.155 -116.120 ;
        RECT 426.000 -117.615 429.325 -117.475 ;
        RECT 426.000 -117.905 431.175 -117.615 ;
        RECT 419.850 -118.280 420.215 -118.010 ;
        RECT 426.000 -118.310 426.430 -117.905 ;
        RECT 427.300 -118.090 427.475 -117.905 ;
        RECT 428.925 -117.920 431.175 -117.905 ;
        RECT 421.740 -118.740 426.430 -118.310 ;
        RECT 420.980 -119.860 421.630 -119.730 ;
        RECT 418.455 -120.190 421.630 -119.860 ;
        RECT 422.440 -120.020 422.610 -118.740 ;
        RECT 422.930 -120.020 423.100 -118.980 ;
        RECT 423.420 -120.020 423.590 -118.740 ;
        RECT 423.910 -119.850 424.080 -118.980 ;
        RECT 426.815 -119.630 426.985 -118.090 ;
        RECT 427.305 -119.630 427.475 -118.090 ;
        RECT 427.795 -119.630 427.965 -118.090 ;
        RECT 428.285 -119.630 428.455 -118.090 ;
        RECT 428.775 -119.630 428.945 -118.090 ;
        RECT 426.655 -119.845 427.010 -119.840 ;
        RECT 428.715 -119.845 429.085 -119.815 ;
        RECT 426.655 -119.850 429.085 -119.845 ;
        RECT 423.910 -120.020 429.085 -119.850 ;
        RECT 430.870 -119.955 431.175 -117.920 ;
        RECT 423.915 -120.040 429.085 -120.020 ;
        RECT 423.915 -120.050 426.660 -120.040 ;
        RECT 421.850 -120.190 422.215 -120.160 ;
        RECT 428.715 -120.170 429.085 -120.040 ;
        RECT 418.455 -120.240 422.215 -120.190 ;
        RECT 420.980 -120.395 422.215 -120.240 ;
        RECT 426.390 -120.330 427.065 -120.290 ;
        RECT 426.290 -120.340 427.065 -120.330 ;
        RECT 420.980 -120.480 421.630 -120.395 ;
        RECT 421.850 -120.460 422.215 -120.395 ;
        RECT 421.115 -120.730 421.495 -120.480 ;
        RECT 425.255 -120.520 427.065 -120.340 ;
        RECT 429.650 -120.385 433.575 -119.955 ;
        RECT 426.290 -120.530 427.065 -120.520 ;
        RECT 426.390 -120.560 427.065 -120.530 ;
        RECT 427.305 -120.445 429.400 -120.405 ;
        RECT 427.305 -120.595 429.455 -120.445 ;
        RECT 422.440 -121.670 422.610 -120.630 ;
        RECT 423.420 -121.670 423.590 -120.630 ;
        RECT 424.400 -121.670 424.570 -120.630 ;
        RECT 427.305 -122.315 427.475 -120.595 ;
        RECT 428.285 -122.315 428.455 -120.595 ;
        RECT 429.150 -121.340 429.455 -120.595 ;
        RECT 430.350 -121.165 430.520 -120.385 ;
        RECT 430.840 -121.165 431.010 -120.625 ;
        RECT 431.330 -121.165 431.500 -120.385 ;
        RECT 431.820 -121.165 431.990 -120.625 ;
        RECT 429.760 -121.340 430.125 -121.310 ;
        RECT 429.150 -121.405 430.125 -121.340 ;
        RECT 429.260 -121.545 430.125 -121.405 ;
        RECT 429.760 -121.610 430.125 -121.545 ;
        RECT 432.310 -121.460 434.170 -121.110 ;
        RECT 430.350 -122.320 430.520 -121.780 ;
        RECT 431.330 -122.320 431.500 -121.780 ;
        RECT 432.310 -122.320 432.480 -121.460 ;
        RECT 430.580 -124.660 431.780 -124.490 ;
        RECT 422.310 -126.995 422.480 -125.275 ;
        RECT 423.290 -126.995 423.460 -125.275 ;
        RECT 425.355 -125.810 425.525 -125.270 ;
        RECT 426.335 -125.810 426.505 -125.270 ;
        RECT 424.765 -126.045 425.130 -125.980 ;
        RECT 424.265 -126.185 425.130 -126.045 ;
        RECT 424.155 -126.250 425.130 -126.185 ;
        RECT 424.155 -126.995 424.460 -126.250 ;
        RECT 424.765 -126.280 425.130 -126.250 ;
        RECT 427.315 -126.130 427.485 -125.270 ;
        RECT 422.310 -127.145 424.460 -126.995 ;
        RECT 422.310 -127.185 424.405 -127.145 ;
        RECT 425.355 -127.205 425.525 -126.425 ;
        RECT 425.845 -126.965 426.015 -126.425 ;
        RECT 426.335 -127.205 426.505 -126.425 ;
        RECT 426.825 -126.965 426.995 -126.425 ;
        RECT 427.315 -126.480 428.705 -126.130 ;
        RECT 420.530 -127.550 421.665 -127.540 ;
        RECT 423.720 -127.550 424.090 -127.420 ;
        RECT 416.820 -127.835 418.245 -127.620 ;
        RECT 420.530 -127.740 424.090 -127.550 ;
        RECT 424.655 -127.635 427.730 -127.205 ;
        RECT 421.660 -127.745 424.090 -127.740 ;
        RECT 421.660 -127.750 422.015 -127.745 ;
        RECT 423.720 -127.775 424.090 -127.745 ;
        RECT 415.425 -128.350 415.950 -127.990 ;
        RECT 418.030 -128.865 418.245 -127.835 ;
        RECT 405.590 -129.605 407.840 -129.515 ;
        RECT 403.380 -129.820 407.840 -129.605 ;
        RECT 403.380 -129.910 405.625 -129.820 ;
        RECT 407.535 -131.295 407.840 -129.820 ;
        RECT 411.205 -130.705 411.375 -129.235 ;
        RECT 411.665 -129.315 411.890 -128.965 ;
        RECT 413.625 -129.065 418.245 -128.865 ;
        RECT 413.865 -129.080 418.245 -129.065 ;
        RECT 411.170 -131.295 411.405 -130.705 ;
        RECT 411.695 -130.775 411.865 -129.315 ;
        RECT 412.185 -130.700 412.355 -129.235 ;
        RECT 413.395 -130.650 413.565 -129.235 ;
        RECT 413.865 -129.280 414.085 -129.080 ;
        RECT 412.150 -131.295 412.385 -130.700 ;
        RECT 413.360 -131.295 413.595 -130.650 ;
        RECT 413.885 -130.775 414.055 -129.280 ;
        RECT 421.820 -129.500 421.990 -127.960 ;
        RECT 422.310 -129.500 422.480 -127.960 ;
        RECT 422.800 -129.500 422.970 -127.960 ;
        RECT 423.290 -129.500 423.460 -127.960 ;
        RECT 423.780 -129.500 423.950 -127.960 ;
        RECT 422.305 -129.760 422.480 -129.500 ;
        RECT 425.875 -129.670 426.180 -127.635 ;
        RECT 428.325 -128.455 428.675 -126.480 ;
        RECT 429.545 -127.750 429.715 -124.830 ;
        RECT 430.580 -124.870 430.790 -124.660 ;
        RECT 429.525 -128.045 429.735 -127.750 ;
        RECT 430.600 -127.780 430.770 -124.870 ;
        RECT 431.090 -127.770 431.260 -124.830 ;
        RECT 431.570 -124.880 431.780 -124.660 ;
        RECT 430.585 -128.045 430.795 -127.780 ;
        RECT 429.525 -128.225 430.795 -128.045 ;
        RECT 431.070 -128.040 431.280 -127.770 ;
        RECT 431.580 -127.870 431.750 -124.880 ;
        RECT 432.640 -127.800 432.810 -124.830 ;
        RECT 431.070 -128.235 431.775 -128.040 ;
        RECT 431.560 -128.295 431.775 -128.235 ;
        RECT 430.350 -128.455 431.125 -128.405 ;
        RECT 428.325 -128.635 431.125 -128.455 ;
        RECT 428.325 -128.645 428.675 -128.635 ;
        RECT 430.350 -128.680 431.125 -128.635 ;
        RECT 431.560 -128.570 432.465 -128.295 ;
        RECT 431.560 -128.920 431.775 -128.570 ;
        RECT 429.000 -128.990 429.775 -128.945 ;
        RECT 428.815 -129.160 429.775 -128.990 ;
        RECT 429.000 -129.220 429.775 -129.160 ;
        RECT 430.005 -129.120 431.775 -128.920 ;
        RECT 432.635 -129.020 432.850 -127.800 ;
        RECT 433.820 -128.145 434.170 -121.460 ;
        RECT 433.765 -128.505 434.290 -128.145 ;
        RECT 436.910 -129.020 438.705 -128.270 ;
        RECT 423.930 -129.760 426.180 -129.670 ;
        RECT 421.720 -129.975 426.180 -129.760 ;
        RECT 421.720 -130.065 423.965 -129.975 ;
        RECT 407.535 -131.860 414.920 -131.295 ;
        RECT 425.875 -131.450 426.180 -129.975 ;
        RECT 429.545 -130.860 429.715 -129.390 ;
        RECT 430.005 -129.470 430.230 -129.120 ;
        RECT 431.965 -129.220 438.705 -129.020 ;
        RECT 432.205 -129.235 438.705 -129.220 ;
        RECT 429.510 -131.450 429.745 -130.860 ;
        RECT 430.035 -130.930 430.205 -129.470 ;
        RECT 430.525 -130.855 430.695 -129.390 ;
        RECT 431.735 -130.805 431.905 -129.390 ;
        RECT 432.205 -129.435 432.425 -129.235 ;
        RECT 430.490 -131.450 430.725 -130.855 ;
        RECT 431.700 -131.450 431.935 -130.805 ;
        RECT 432.225 -130.930 432.395 -129.435 ;
        RECT 436.910 -129.985 438.705 -129.235 ;
        RECT 425.875 -132.015 433.260 -131.450 ;
        RECT 398.025 -140.745 399.960 -139.365 ;
        RECT -121.005 -148.995 -119.940 -148.835 ;
        RECT -123.785 -149.675 50.770 -148.995 ;
        RECT -121.005 -149.725 -119.940 -149.675 ;
        RECT -40.035 -150.975 84.685 -150.295 ;
        RECT -123.785 -152.160 52.055 -151.485 ;
        RECT -138.020 -185.870 -137.320 -185.020 ;
        RECT -135.145 -185.870 -134.545 -170.430 ;
        RECT -132.080 -170.585 -131.620 -170.455 ;
        RECT -134.120 -170.755 -131.620 -170.585 ;
        RECT -132.080 -171.175 -131.620 -170.755 ;
        RECT -134.120 -171.345 -131.620 -171.175 ;
        RECT -132.080 -171.765 -131.620 -171.345 ;
        RECT -134.120 -171.935 -131.620 -171.765 ;
        RECT -132.080 -172.355 -131.620 -171.935 ;
        RECT -134.120 -172.525 -131.620 -172.355 ;
        RECT -132.080 -172.945 -131.620 -172.525 ;
        RECT -134.120 -173.115 -131.620 -172.945 ;
        RECT -132.080 -173.535 -131.620 -173.115 ;
        RECT -134.120 -173.705 -131.620 -173.535 ;
        RECT -132.080 -174.125 -131.620 -173.705 ;
        RECT -134.120 -174.295 -131.620 -174.125 ;
        RECT -132.080 -174.715 -131.620 -174.295 ;
        RECT 41.205 -171.010 97.545 -169.345 ;
        RECT -134.120 -174.885 -131.620 -174.715 ;
        RECT -132.080 -175.305 -131.620 -174.885 ;
        RECT -64.480 -174.825 -61.340 -174.655 ;
        RECT -71.715 -174.940 -71.545 -174.920 ;
        RECT -134.120 -175.475 -131.620 -175.305 ;
        RECT -132.080 -175.895 -131.620 -175.475 ;
        RECT -134.120 -176.065 -131.620 -175.895 ;
        RECT -132.080 -176.485 -131.620 -176.065 ;
        RECT -71.745 -176.205 -71.515 -174.940 ;
        RECT -70.735 -175.880 -70.565 -174.920 ;
        RECT -69.755 -175.880 -69.585 -174.920 ;
        RECT -67.530 -174.940 -67.360 -174.920 ;
        RECT -68.635 -175.350 -68.350 -175.030 ;
        RECT -69.350 -175.595 -68.350 -175.350 ;
        RECT -70.765 -176.205 -70.535 -175.880 ;
        RECT -69.785 -176.205 -69.555 -175.880 ;
        RECT -71.745 -176.245 -69.555 -176.205 ;
        RECT -69.350 -176.245 -69.120 -175.595 ;
        RECT -68.635 -175.850 -68.350 -175.595 ;
        RECT -72.765 -176.430 -71.925 -176.280 ;
        RECT -134.120 -176.655 -131.620 -176.485 ;
        RECT -132.080 -177.075 -131.620 -176.655 ;
        RECT -134.120 -177.245 -131.620 -177.075 ;
        RECT -132.080 -177.665 -131.620 -177.245 ;
        RECT -134.120 -177.835 -131.620 -177.665 ;
        RECT -132.080 -178.255 -131.620 -177.835 ;
        RECT -134.120 -178.425 -131.620 -178.255 ;
        RECT -132.080 -178.845 -131.620 -178.425 ;
        RECT -72.800 -176.650 -71.925 -176.430 ;
        RECT -71.745 -176.435 -69.120 -176.245 ;
        RECT -67.560 -176.205 -67.330 -174.940 ;
        RECT -66.550 -175.880 -66.380 -174.920 ;
        RECT -65.570 -175.880 -65.400 -174.920 ;
        RECT -64.480 -175.050 -64.300 -174.825 ;
        RECT -66.580 -176.205 -66.350 -175.880 ;
        RECT -65.600 -176.205 -65.370 -175.880 ;
        RECT -67.560 -176.245 -65.370 -176.205 ;
        RECT -65.095 -176.125 -64.725 -175.285 ;
        RECT -64.475 -175.420 -64.305 -175.050 ;
        RECT -65.095 -176.245 -64.730 -176.125 ;
        RECT -68.580 -176.335 -67.740 -176.280 ;
        RECT -68.755 -176.340 -67.740 -176.335 ;
        RECT -72.800 -178.510 -72.560 -176.650 ;
        RECT -72.205 -177.615 -72.035 -176.820 ;
        RECT -71.745 -176.900 -71.515 -176.435 ;
        RECT -71.715 -177.360 -71.545 -176.900 ;
        RECT -71.225 -177.615 -71.055 -176.820 ;
        RECT -70.765 -176.900 -70.535 -176.435 ;
        RECT -69.785 -176.595 -69.120 -176.435 ;
        RECT -70.735 -177.360 -70.565 -176.900 ;
        RECT -70.245 -177.615 -70.075 -176.820 ;
        RECT -69.785 -176.900 -69.555 -176.595 ;
        RECT -68.940 -176.650 -67.740 -176.340 ;
        RECT -67.560 -176.435 -64.730 -176.245 ;
        RECT -69.755 -177.360 -69.585 -176.900 ;
        RECT -68.940 -177.370 -68.640 -176.650 ;
        RECT -68.020 -177.615 -67.850 -176.820 ;
        RECT -67.560 -176.900 -67.330 -176.435 ;
        RECT -67.530 -177.360 -67.360 -176.900 ;
        RECT -67.040 -177.615 -66.870 -176.820 ;
        RECT -66.580 -176.900 -66.350 -176.435 ;
        RECT -65.600 -176.595 -64.730 -176.435 ;
        RECT -64.505 -176.155 -64.270 -175.420 ;
        RECT -63.985 -175.455 -63.815 -174.995 ;
        RECT -63.500 -175.100 -63.290 -174.825 ;
        RECT -63.990 -175.715 -63.810 -175.455 ;
        RECT -63.495 -175.535 -63.325 -175.100 ;
        RECT -63.005 -175.445 -62.835 -174.995 ;
        RECT -62.530 -175.105 -62.320 -174.825 ;
        RECT -63.005 -175.535 -62.820 -175.445 ;
        RECT -62.515 -175.535 -62.345 -175.105 ;
        RECT -62.025 -175.445 -61.855 -174.995 ;
        RECT -61.550 -175.080 -61.340 -174.825 ;
        RECT -50.980 -174.825 -47.840 -174.655 ;
        RECT -58.215 -174.940 -58.045 -174.920 ;
        RECT -63.000 -175.715 -62.820 -175.535 ;
        RECT -62.030 -175.715 -61.850 -175.445 ;
        RECT -61.535 -175.535 -61.365 -175.080 ;
        RECT -61.045 -175.495 -60.875 -174.995 ;
        RECT -61.060 -175.715 -60.850 -175.495 ;
        RECT -63.990 -175.885 -60.850 -175.715 ;
        RECT -64.505 -176.525 -63.645 -176.155 ;
        RECT -61.725 -176.420 -60.850 -175.885 ;
        RECT -58.245 -176.205 -58.015 -174.940 ;
        RECT -57.235 -175.880 -57.065 -174.920 ;
        RECT -56.255 -175.880 -56.085 -174.920 ;
        RECT -54.030 -174.940 -53.860 -174.920 ;
        RECT -55.135 -175.290 -54.850 -175.030 ;
        RECT -55.875 -175.600 -54.850 -175.290 ;
        RECT -57.265 -176.205 -57.035 -175.880 ;
        RECT -56.285 -176.205 -56.055 -175.880 ;
        RECT -58.245 -176.245 -56.055 -176.205 ;
        RECT -55.875 -176.245 -55.565 -175.600 ;
        RECT -55.135 -175.850 -54.850 -175.600 ;
        RECT -59.265 -176.315 -58.425 -176.280 ;
        RECT -66.550 -177.360 -66.380 -176.900 ;
        RECT -66.060 -177.615 -65.890 -176.820 ;
        RECT -65.600 -176.900 -65.370 -176.595 ;
        RECT -65.570 -177.360 -65.400 -176.900 ;
        RECT -64.505 -177.200 -64.270 -176.525 ;
        RECT -61.725 -176.720 -60.395 -176.420 ;
        RECT -59.375 -176.615 -58.425 -176.315 ;
        RECT -59.265 -176.650 -58.425 -176.615 ;
        RECT -58.245 -176.435 -55.565 -176.245 ;
        RECT -54.060 -176.205 -53.830 -174.940 ;
        RECT -53.050 -175.880 -52.880 -174.920 ;
        RECT -52.070 -175.880 -51.900 -174.920 ;
        RECT -50.980 -175.050 -50.800 -174.825 ;
        RECT -53.080 -176.205 -52.850 -175.880 ;
        RECT -52.100 -176.205 -51.870 -175.880 ;
        RECT -54.060 -176.245 -51.870 -176.205 ;
        RECT -51.595 -176.125 -51.225 -175.285 ;
        RECT -50.975 -175.420 -50.805 -175.050 ;
        RECT -51.595 -176.245 -51.230 -176.125 ;
        RECT -55.080 -176.335 -54.240 -176.280 ;
        RECT -64.005 -176.890 -60.850 -176.720 ;
        RECT -64.005 -177.095 -63.800 -176.890 ;
        RECT -64.475 -177.550 -64.305 -177.200 ;
        RECT -72.250 -177.955 -65.395 -177.615 ;
        RECT -64.500 -177.840 -64.280 -177.550 ;
        RECT -63.985 -177.610 -63.815 -177.095 ;
        RECT -63.495 -177.495 -63.325 -177.070 ;
        RECT -63.015 -177.135 -62.810 -176.890 ;
        RECT -63.520 -177.840 -63.300 -177.495 ;
        RECT -63.005 -177.610 -62.835 -177.135 ;
        RECT -62.515 -177.495 -62.345 -177.070 ;
        RECT -62.045 -177.135 -61.840 -176.890 ;
        RECT -61.060 -176.925 -60.850 -176.890 ;
        RECT -62.540 -177.840 -62.320 -177.495 ;
        RECT -62.025 -177.610 -61.855 -177.135 ;
        RECT -61.535 -177.550 -61.365 -177.070 ;
        RECT -61.060 -177.140 -60.855 -176.925 ;
        RECT -61.555 -177.840 -61.335 -177.550 ;
        RECT -61.045 -177.610 -60.875 -177.140 ;
        RECT -58.705 -177.615 -58.535 -176.820 ;
        RECT -58.245 -176.900 -58.015 -176.435 ;
        RECT -58.215 -177.360 -58.045 -176.900 ;
        RECT -57.725 -177.615 -57.555 -176.820 ;
        RECT -57.265 -176.900 -57.035 -176.435 ;
        RECT -56.285 -176.595 -55.565 -176.435 ;
        RECT -57.235 -177.360 -57.065 -176.900 ;
        RECT -56.745 -177.615 -56.575 -176.820 ;
        RECT -56.285 -176.900 -56.055 -176.595 ;
        RECT -55.380 -176.650 -54.240 -176.335 ;
        RECT -54.060 -176.435 -51.230 -176.245 ;
        RECT -56.255 -177.360 -56.085 -176.900 ;
        RECT -55.380 -177.445 -55.080 -176.650 ;
        RECT -54.520 -177.615 -54.350 -176.820 ;
        RECT -54.060 -176.900 -53.830 -176.435 ;
        RECT -54.030 -177.360 -53.860 -176.900 ;
        RECT -53.540 -177.615 -53.370 -176.820 ;
        RECT -53.080 -176.900 -52.850 -176.435 ;
        RECT -52.100 -176.595 -51.230 -176.435 ;
        RECT -51.005 -176.155 -50.770 -175.420 ;
        RECT -50.485 -175.455 -50.315 -174.995 ;
        RECT -50.000 -175.100 -49.790 -174.825 ;
        RECT -50.490 -175.715 -50.310 -175.455 ;
        RECT -49.995 -175.535 -49.825 -175.100 ;
        RECT -49.505 -175.445 -49.335 -174.995 ;
        RECT -49.030 -175.105 -48.820 -174.825 ;
        RECT -49.505 -175.535 -49.320 -175.445 ;
        RECT -49.015 -175.535 -48.845 -175.105 ;
        RECT -48.525 -175.445 -48.355 -174.995 ;
        RECT -48.050 -175.080 -47.840 -174.825 ;
        RECT -39.855 -174.800 -38.655 -174.630 ;
        RECT -49.500 -175.715 -49.320 -175.535 ;
        RECT -48.530 -175.715 -48.350 -175.445 ;
        RECT -48.035 -175.535 -47.865 -175.080 ;
        RECT -47.545 -175.495 -47.375 -174.995 ;
        RECT -47.560 -175.715 -47.350 -175.495 ;
        RECT -50.490 -175.885 -47.350 -175.715 ;
        RECT -51.005 -176.525 -50.145 -176.155 ;
        RECT -48.225 -176.430 -47.350 -175.885 ;
        RECT -53.050 -177.360 -52.880 -176.900 ;
        RECT -52.560 -177.615 -52.390 -176.820 ;
        RECT -52.100 -176.900 -51.870 -176.595 ;
        RECT -52.070 -177.360 -51.900 -176.900 ;
        RECT -51.005 -177.200 -50.770 -176.525 ;
        RECT -48.225 -176.720 -46.975 -176.430 ;
        RECT -50.505 -176.730 -46.975 -176.720 ;
        RECT -50.505 -176.890 -47.350 -176.730 ;
        RECT -50.505 -177.095 -50.300 -176.890 ;
        RECT -50.975 -177.550 -50.805 -177.200 ;
        RECT -71.010 -178.155 -70.455 -177.955 ;
        RECT -71.065 -178.195 -70.380 -178.155 ;
        RECT -66.955 -178.195 -66.400 -177.955 ;
        RECT -64.500 -178.010 -61.335 -177.840 ;
        RECT -58.750 -177.625 -56.080 -177.615 ;
        RECT -54.565 -177.625 -51.895 -177.615 ;
        RECT -58.750 -177.955 -51.895 -177.625 ;
        RECT -51.000 -177.840 -50.780 -177.550 ;
        RECT -50.485 -177.610 -50.315 -177.095 ;
        RECT -49.995 -177.495 -49.825 -177.070 ;
        RECT -49.515 -177.135 -49.310 -176.890 ;
        RECT -50.020 -177.840 -49.800 -177.495 ;
        RECT -49.505 -177.610 -49.335 -177.135 ;
        RECT -49.015 -177.495 -48.845 -177.070 ;
        RECT -48.545 -177.135 -48.340 -176.890 ;
        RECT -47.560 -176.925 -47.350 -176.890 ;
        RECT -49.040 -177.840 -48.820 -177.495 ;
        RECT -48.525 -177.610 -48.355 -177.135 ;
        RECT -48.035 -177.550 -47.865 -177.070 ;
        RECT -47.560 -177.140 -47.355 -176.925 ;
        RECT -48.055 -177.840 -47.835 -177.550 ;
        RECT -47.545 -177.610 -47.375 -177.140 ;
        RECT -57.965 -178.185 -57.410 -177.955 ;
        RECT -57.050 -177.965 -54.450 -177.955 ;
        RECT -58.080 -178.195 -57.395 -178.185 ;
        RECT -53.575 -178.195 -53.020 -177.955 ;
        RECT -51.000 -178.010 -47.835 -177.840 ;
        RECT -40.885 -177.940 -40.715 -174.970 ;
        RECT -39.855 -175.020 -39.645 -174.800 ;
        RECT -44.890 -178.195 -44.230 -178.185 ;
        RECT -71.150 -178.390 -44.225 -178.195 ;
        RECT -71.065 -178.455 -70.380 -178.390 ;
        RECT -58.080 -178.485 -57.395 -178.390 ;
        RECT -44.890 -178.485 -44.230 -178.390 ;
        RECT -134.120 -179.015 -131.620 -178.845 ;
        RECT -132.080 -179.435 -131.620 -179.015 ;
        RECT -134.120 -179.605 -131.620 -179.435 ;
        RECT -132.080 -180.025 -131.620 -179.605 ;
        RECT -134.120 -180.195 -131.620 -180.025 ;
        RECT -132.080 -180.615 -131.620 -180.195 ;
        RECT -109.710 -180.075 -109.540 -178.855 ;
        RECT -108.730 -180.075 -108.560 -178.855 ;
        RECT -107.750 -180.075 -107.580 -178.855 ;
        RECT -109.710 -180.260 -106.935 -180.075 ;
        RECT -134.120 -180.785 -131.620 -180.615 ;
        RECT -132.080 -181.205 -131.620 -180.785 ;
        RECT -134.120 -181.375 -131.620 -181.205 ;
        RECT -132.080 -181.795 -131.620 -181.375 ;
        RECT -107.120 -180.950 -106.935 -180.260 ;
        RECT -104.910 -180.950 -104.235 -180.900 ;
        RECT -107.120 -181.135 -104.235 -180.950 ;
        RECT -107.120 -181.405 -106.935 -181.135 ;
        RECT -104.910 -181.170 -104.235 -181.135 ;
        RECT -134.120 -181.965 -131.620 -181.795 ;
        RECT -132.080 -182.385 -131.620 -181.965 ;
        RECT -134.120 -182.555 -131.620 -182.385 ;
        RECT -132.080 -182.975 -131.620 -182.555 ;
        RECT -134.120 -183.145 -131.620 -182.975 ;
        RECT -132.080 -183.565 -131.620 -183.145 ;
        RECT -110.200 -181.575 -107.985 -181.405 ;
        RECT -107.120 -181.575 -105.955 -181.405 ;
        RECT -110.200 -183.430 -110.030 -181.575 ;
        RECT -109.220 -181.580 -107.985 -181.575 ;
        RECT -134.120 -183.735 -131.620 -183.565 ;
        RECT -132.080 -184.155 -131.620 -183.735 ;
        RECT -134.120 -184.325 -131.620 -184.155 ;
        RECT -132.080 -184.745 -131.620 -184.325 ;
        RECT -109.710 -184.375 -109.540 -181.890 ;
        RECT -109.220 -183.430 -109.050 -181.580 ;
        RECT -108.160 -181.895 -107.985 -181.580 ;
        RECT -108.650 -183.390 -108.480 -181.895 ;
        RECT -108.650 -183.910 -108.475 -183.390 ;
        RECT -108.160 -183.435 -107.990 -181.895 ;
        RECT -107.670 -183.380 -107.500 -181.895 ;
        RECT -107.670 -183.910 -107.495 -183.380 ;
        RECT -107.105 -183.435 -106.935 -181.575 ;
        RECT -108.650 -183.925 -107.495 -183.910 ;
        RECT -106.615 -183.925 -106.445 -181.895 ;
        RECT -106.125 -183.435 -105.955 -181.575 ;
        RECT -108.650 -184.095 -106.445 -183.925 ;
        RECT -104.550 -183.930 -104.380 -182.395 ;
        RECT -104.060 -183.435 -103.890 -178.855 ;
        RECT -101.780 -181.260 -101.095 -181.175 ;
        RECT -99.715 -181.185 -99.545 -179.465 ;
        RECT -98.735 -181.185 -98.565 -179.465 ;
        RECT -96.670 -180.000 -96.500 -179.460 ;
        RECT -95.690 -180.000 -95.520 -179.460 ;
        RECT -97.260 -180.235 -96.895 -180.170 ;
        RECT -97.760 -180.375 -96.895 -180.235 ;
        RECT -97.870 -180.440 -96.895 -180.375 ;
        RECT -97.870 -181.185 -97.565 -180.440 ;
        RECT -97.260 -180.470 -96.895 -180.440 ;
        RECT -94.710 -180.320 -94.540 -179.460 ;
        RECT -87.970 -179.640 -80.585 -179.075 ;
        RECT -72.805 -179.195 -72.505 -178.510 ;
        RECT -60.255 -178.655 -59.570 -178.600 ;
        RECT -55.525 -178.655 -54.865 -178.605 ;
        RECT -71.150 -178.850 -42.500 -178.655 ;
        RECT -60.255 -178.900 -59.570 -178.850 ;
        RECT -55.525 -178.905 -54.865 -178.850 ;
        RECT -69.120 -179.085 -68.460 -179.045 ;
        RECT -46.505 -179.085 -45.845 -179.035 ;
        RECT -94.710 -180.325 -92.690 -180.320 ;
        RECT -94.710 -180.615 -92.370 -180.325 ;
        RECT -100.630 -181.250 -99.955 -181.220 ;
        RECT -100.730 -181.260 -99.955 -181.250 ;
        RECT -101.780 -181.440 -99.955 -181.260 ;
        RECT -99.715 -181.335 -97.565 -181.185 ;
        RECT -99.715 -181.375 -97.620 -181.335 ;
        RECT -96.670 -181.395 -96.500 -180.615 ;
        RECT -96.180 -181.155 -96.010 -180.615 ;
        RECT -95.690 -181.395 -95.520 -180.615 ;
        RECT -95.200 -181.155 -95.030 -180.615 ;
        RECT -94.710 -180.670 -92.690 -180.615 ;
        RECT -92.125 -181.115 -89.880 -181.025 ;
        RECT -87.970 -181.115 -87.665 -179.640 ;
        RECT -84.335 -180.230 -84.100 -179.640 ;
        RECT -94.505 -181.395 -87.665 -181.115 ;
        RECT -101.780 -181.465 -101.095 -181.440 ;
        RECT -100.730 -181.450 -99.955 -181.440 ;
        RECT -100.630 -181.490 -99.955 -181.450 ;
        RECT -97.370 -181.420 -87.665 -181.395 ;
        RECT -97.370 -181.825 -94.200 -181.420 ;
        RECT -91.540 -181.590 -91.365 -181.420 ;
        RECT -100.205 -183.690 -100.035 -182.150 ;
        RECT -99.715 -183.690 -99.545 -182.150 ;
        RECT -99.225 -183.690 -99.055 -182.150 ;
        RECT -98.735 -183.690 -98.565 -182.150 ;
        RECT -98.245 -183.690 -98.075 -182.150 ;
        RECT -99.720 -183.930 -99.545 -183.690 ;
        RECT -96.150 -183.860 -95.845 -181.825 ;
        RECT -94.505 -181.835 -94.200 -181.825 ;
        RECT -92.025 -183.130 -91.855 -181.590 ;
        RECT -91.535 -183.130 -91.365 -181.590 ;
        RECT -91.045 -183.130 -90.875 -181.590 ;
        RECT -90.555 -183.130 -90.385 -181.590 ;
        RECT -90.065 -183.130 -89.895 -181.590 ;
        RECT -92.185 -183.345 -91.830 -183.340 ;
        RECT -90.125 -183.345 -89.755 -183.315 ;
        RECT -92.185 -183.350 -89.755 -183.345 ;
        RECT -93.315 -183.540 -89.755 -183.350 ;
        RECT -87.970 -183.455 -87.665 -181.420 ;
        RECT -84.300 -181.700 -84.130 -180.230 ;
        RECT -83.810 -181.620 -83.640 -180.160 ;
        RECT -83.355 -180.235 -83.120 -179.640 ;
        RECT -84.845 -181.930 -84.070 -181.870 ;
        RECT -85.030 -182.100 -84.070 -181.930 ;
        RECT -84.845 -182.145 -84.070 -182.100 ;
        RECT -83.840 -181.970 -83.615 -181.620 ;
        RECT -83.320 -181.700 -83.150 -180.235 ;
        RECT -82.145 -180.285 -81.910 -179.640 ;
        RECT -82.110 -181.700 -81.940 -180.285 ;
        RECT -81.620 -181.655 -81.450 -180.160 ;
        RECT -72.800 -180.985 -72.560 -179.195 ;
        RECT -71.150 -179.280 -45.845 -179.085 ;
        RECT -42.695 -179.160 -42.500 -178.850 ;
        RECT -40.925 -179.160 -40.710 -177.940 ;
        RECT -39.825 -178.010 -39.655 -175.020 ;
        RECT -39.335 -177.910 -39.165 -174.970 ;
        RECT -38.865 -175.010 -38.655 -174.800 ;
        RECT -39.355 -178.180 -39.145 -177.910 ;
        RECT -38.845 -177.920 -38.675 -175.010 ;
        RECT -37.790 -177.890 -37.620 -174.970 ;
        RECT -33.735 -175.430 -30.095 -175.260 ;
        RECT -33.735 -176.990 -33.565 -175.430 ;
        RECT -33.245 -177.170 -33.075 -175.950 ;
        RECT -32.755 -176.990 -32.585 -175.430 ;
        RECT -32.155 -175.775 -30.445 -175.605 ;
        RECT -32.155 -176.990 -31.985 -175.775 ;
        RECT -31.665 -177.170 -31.495 -175.950 ;
        RECT -31.175 -176.990 -31.005 -175.775 ;
        RECT -34.290 -177.340 -30.920 -177.170 ;
        RECT -39.850 -178.375 -39.145 -178.180 ;
        RECT -38.870 -178.185 -38.660 -177.920 ;
        RECT -37.810 -178.185 -37.600 -177.890 ;
        RECT -38.870 -178.365 -37.600 -178.185 ;
        RECT -39.850 -178.435 -39.635 -178.375 ;
        RECT -40.540 -178.710 -39.635 -178.435 ;
        RECT -39.850 -179.060 -39.635 -178.710 ;
        RECT -39.200 -178.595 -38.425 -178.545 ;
        RECT -36.500 -178.595 -35.840 -178.240 ;
        RECT -39.200 -178.775 -35.840 -178.595 ;
        RECT -39.200 -178.820 -38.425 -178.775 ;
        RECT -69.120 -179.345 -68.460 -179.280 ;
        RECT -46.505 -179.335 -45.845 -179.280 ;
        RECT -42.715 -179.360 -40.040 -179.160 ;
        RECT -39.850 -179.260 -38.080 -179.060 ;
        RECT -42.715 -179.375 -40.280 -179.360 ;
        RECT -72.210 -179.855 -69.540 -179.515 ;
        RECT -67.555 -179.630 -64.390 -179.460 ;
        RECT -72.205 -180.570 -72.035 -180.110 ;
        RECT -72.235 -180.875 -72.005 -180.570 ;
        RECT -71.715 -180.650 -71.545 -179.855 ;
        RECT -71.225 -180.570 -71.055 -180.110 ;
        RECT -72.385 -180.985 -72.005 -180.875 ;
        RECT -72.800 -181.035 -72.005 -180.985 ;
        RECT -71.255 -181.035 -71.025 -180.570 ;
        RECT -70.735 -180.650 -70.565 -179.855 ;
        RECT -70.245 -180.570 -70.075 -180.110 ;
        RECT -70.275 -181.035 -70.045 -180.570 ;
        RECT -69.755 -180.650 -69.585 -179.855 ;
        RECT -68.015 -180.330 -67.845 -179.860 ;
        RECT -67.555 -179.920 -67.335 -179.630 ;
        RECT -68.035 -180.545 -67.830 -180.330 ;
        RECT -67.525 -180.400 -67.355 -179.920 ;
        RECT -67.035 -180.335 -66.865 -179.860 ;
        RECT -66.570 -179.975 -66.350 -179.630 ;
        RECT -68.040 -180.580 -67.830 -180.545 ;
        RECT -67.050 -180.580 -66.845 -180.335 ;
        RECT -66.545 -180.400 -66.375 -179.975 ;
        RECT -66.055 -180.335 -65.885 -179.860 ;
        RECT -65.590 -179.975 -65.370 -179.630 ;
        RECT -66.080 -180.580 -65.875 -180.335 ;
        RECT -65.565 -180.400 -65.395 -179.975 ;
        RECT -65.075 -180.375 -64.905 -179.860 ;
        RECT -64.610 -179.920 -64.390 -179.630 ;
        RECT -63.495 -179.855 -56.040 -179.515 ;
        RECT -54.055 -179.630 -50.890 -179.460 ;
        RECT -64.585 -180.270 -64.415 -179.920 ;
        RECT -65.090 -180.580 -64.885 -180.375 ;
        RECT -68.040 -180.750 -64.885 -180.580 ;
        RECT -72.800 -181.170 -70.045 -181.035 ;
        RECT -72.795 -181.180 -70.045 -181.170 ;
        RECT -72.385 -181.225 -70.045 -181.180 ;
        RECT -69.865 -180.895 -69.025 -180.820 ;
        RECT -68.040 -180.895 -67.165 -180.750 ;
        RECT -69.865 -181.160 -67.165 -180.895 ;
        RECT -64.620 -180.945 -64.385 -180.270 ;
        RECT -63.490 -180.570 -63.320 -180.110 ;
        RECT -63.520 -180.875 -63.290 -180.570 ;
        RECT -63.000 -180.650 -62.830 -179.855 ;
        RECT -62.510 -180.570 -62.340 -180.110 ;
        RECT -69.865 -181.190 -69.025 -181.160 ;
        RECT -72.235 -181.265 -70.045 -181.225 ;
        RECT -72.235 -181.590 -72.005 -181.265 ;
        RECT -71.255 -181.590 -71.025 -181.265 ;
        RECT -81.640 -181.855 -81.420 -181.655 ;
        RECT -81.640 -181.870 -75.940 -181.855 ;
        RECT -83.840 -182.170 -82.070 -181.970 ;
        RECT -81.880 -182.070 -75.940 -181.870 ;
        RECT -85.520 -182.455 -85.170 -182.445 ;
        RECT -83.495 -182.455 -82.720 -182.410 ;
        RECT -85.520 -182.635 -82.720 -182.455 ;
        RECT -93.315 -183.550 -92.180 -183.540 ;
        RECT -90.125 -183.670 -89.755 -183.540 ;
        RECT -98.095 -183.930 -95.845 -183.860 ;
        RECT -89.190 -183.885 -86.115 -183.455 ;
        RECT -105.475 -184.375 -95.695 -183.930 ;
        RECT -134.120 -184.915 -131.620 -184.745 ;
        RECT -132.080 -185.335 -131.620 -184.915 ;
        RECT -134.120 -185.505 -131.620 -185.335 ;
        RECT -138.020 -186.755 -134.545 -185.870 ;
        RECT -132.080 -185.925 -131.620 -185.505 ;
        RECT -113.370 -185.495 -113.065 -184.605 ;
        RECT -110.200 -184.690 -95.695 -184.375 ;
        RECT -91.535 -183.945 -89.440 -183.905 ;
        RECT -91.535 -184.095 -89.385 -183.945 ;
        RECT -110.200 -184.700 -103.830 -184.690 ;
        RECT -101.930 -185.495 -101.665 -185.015 ;
        RECT -113.370 -185.675 -101.665 -185.495 ;
        RECT -113.370 -185.685 -113.065 -185.675 ;
        RECT -91.535 -185.815 -91.365 -184.095 ;
        RECT -90.555 -185.815 -90.385 -184.095 ;
        RECT -89.690 -184.840 -89.385 -184.095 ;
        RECT -88.490 -184.665 -88.320 -183.885 ;
        RECT -88.000 -184.665 -87.830 -184.125 ;
        RECT -87.510 -184.665 -87.340 -183.885 ;
        RECT -87.020 -184.665 -86.850 -184.125 ;
        RECT -85.520 -184.610 -85.170 -182.635 ;
        RECT -83.495 -182.685 -82.720 -182.635 ;
        RECT -82.285 -182.520 -82.070 -182.170 ;
        RECT -82.285 -182.795 -81.380 -182.520 ;
        RECT -82.285 -182.855 -82.070 -182.795 ;
        RECT -84.320 -183.045 -83.050 -182.865 ;
        RECT -84.320 -183.340 -84.110 -183.045 ;
        RECT -83.260 -183.310 -83.050 -183.045 ;
        RECT -82.775 -183.050 -82.070 -182.855 ;
        RECT -89.080 -184.840 -88.715 -184.810 ;
        RECT -89.690 -184.905 -88.715 -184.840 ;
        RECT -89.580 -185.045 -88.715 -184.905 ;
        RECT -89.080 -185.110 -88.715 -185.045 ;
        RECT -86.530 -184.960 -85.140 -184.610 ;
        RECT -88.490 -185.820 -88.320 -185.280 ;
        RECT -87.510 -185.820 -87.340 -185.280 ;
        RECT -86.530 -185.820 -86.360 -184.960 ;
        RECT -134.120 -186.095 -131.620 -185.925 ;
        RECT -132.080 -186.515 -131.620 -186.095 ;
        RECT -84.300 -186.260 -84.130 -183.340 ;
        RECT -83.245 -186.220 -83.075 -183.310 ;
        RECT -82.775 -183.320 -82.565 -183.050 ;
        RECT -134.120 -186.685 -131.620 -186.515 ;
        RECT -83.265 -186.430 -83.055 -186.220 ;
        RECT -82.755 -186.260 -82.585 -183.320 ;
        RECT -82.265 -186.210 -82.095 -183.220 ;
        RECT -81.210 -183.290 -80.995 -182.070 ;
        RECT -80.080 -182.945 -79.555 -182.585 ;
        RECT -82.275 -186.430 -82.065 -186.210 ;
        RECT -81.205 -186.260 -81.035 -183.290 ;
        RECT -83.265 -186.600 -82.065 -186.430 ;
        RECT -138.020 -188.425 -137.320 -186.755 ;
        RECT -135.145 -188.285 -134.545 -186.755 ;
        RECT -132.080 -187.105 -131.620 -186.685 ;
        RECT -134.120 -187.275 -131.620 -187.105 ;
        RECT -132.080 -187.695 -131.620 -187.275 ;
        RECT -134.120 -187.865 -131.620 -187.695 ;
        RECT -132.080 -188.285 -131.760 -187.865 ;
        RECT -135.145 -188.425 -131.760 -188.285 ;
        RECT -138.020 -188.455 -131.760 -188.425 ;
        RECT -138.020 -189.310 -134.545 -188.455 ;
        RECT -132.080 -188.605 -131.760 -188.455 ;
        RECT -131.590 -188.845 -130.810 -188.485 ;
        RECT -138.020 -191.500 -137.320 -189.310 ;
        RECT -135.145 -189.465 -134.545 -189.310 ;
        RECT -135.145 -189.635 -132.080 -189.465 ;
        RECT -135.145 -190.645 -134.545 -189.635 ;
        RECT -131.250 -190.215 -131.080 -188.845 ;
        RECT -131.250 -190.385 -128.040 -190.215 ;
        RECT -135.145 -190.815 -132.080 -190.645 ;
        RECT -112.075 -190.805 -111.775 -189.810 ;
        RECT -109.425 -190.730 -109.255 -189.010 ;
        RECT -108.445 -190.730 -108.275 -189.010 ;
        RECT -106.380 -189.545 -106.210 -189.005 ;
        RECT -105.400 -189.545 -105.230 -189.005 ;
        RECT -106.970 -189.780 -106.605 -189.715 ;
        RECT -107.470 -189.920 -106.605 -189.780 ;
        RECT -107.580 -189.985 -106.605 -189.920 ;
        RECT -107.580 -190.730 -107.275 -189.985 ;
        RECT -106.970 -190.015 -106.605 -189.985 ;
        RECT -104.420 -189.865 -104.250 -189.005 ;
        RECT -100.560 -189.755 -100.390 -188.535 ;
        RECT -99.580 -189.755 -99.410 -188.535 ;
        RECT -98.600 -189.755 -98.430 -188.535 ;
        RECT -101.435 -189.810 -100.760 -189.770 ;
        RECT -103.235 -189.865 -100.760 -189.810 ;
        RECT -104.420 -189.985 -100.760 -189.865 ;
        RECT -100.560 -189.940 -97.785 -189.755 ;
        RECT -110.340 -190.795 -109.665 -190.765 ;
        RECT -110.440 -190.805 -109.665 -190.795 ;
        RECT -135.145 -191.500 -134.545 -190.815 ;
        RECT -112.075 -190.985 -109.665 -190.805 ;
        RECT -109.425 -190.880 -107.275 -190.730 ;
        RECT -109.425 -190.920 -107.330 -190.880 ;
        RECT -106.380 -190.940 -106.210 -190.160 ;
        RECT -105.890 -190.700 -105.720 -190.160 ;
        RECT -105.400 -190.940 -105.230 -190.160 ;
        RECT -104.910 -190.700 -104.740 -190.160 ;
        RECT -104.420 -190.215 -103.030 -189.985 ;
        RECT -101.530 -189.995 -100.760 -189.985 ;
        RECT -101.435 -190.040 -100.760 -189.995 ;
        RECT -102.010 -190.225 -101.720 -190.185 ;
        RECT -99.755 -190.225 -99.080 -190.180 ;
        RECT -102.140 -190.415 -99.080 -190.225 ;
        RECT -112.075 -190.995 -111.775 -190.985 ;
        RECT -110.440 -190.995 -109.665 -190.985 ;
        RECT -110.340 -191.035 -109.665 -190.995 ;
        RECT -112.705 -191.285 -110.070 -191.275 ;
        RECT -108.015 -191.285 -107.645 -191.155 ;
        RECT -138.020 -191.825 -134.545 -191.500 ;
        RECT -130.080 -191.565 -128.040 -191.395 ;
        RECT -112.705 -191.475 -107.645 -191.285 ;
        RECT -107.080 -191.370 -104.005 -190.940 ;
        RECT -138.020 -191.995 -132.080 -191.825 ;
        RECT -138.020 -192.385 -134.545 -191.995 ;
        RECT -112.705 -192.000 -112.505 -191.475 ;
        RECT -110.075 -191.480 -107.645 -191.475 ;
        RECT -110.075 -191.485 -109.720 -191.480 ;
        RECT -108.015 -191.510 -107.645 -191.480 ;
        RECT -138.020 -195.460 -137.320 -192.385 ;
        RECT -135.145 -193.005 -134.545 -192.385 ;
        RECT -130.080 -192.745 -128.040 -192.575 ;
        RECT -135.145 -193.175 -132.080 -193.005 ;
        RECT -135.145 -194.185 -134.545 -193.175 ;
        RECT -112.790 -193.185 -112.490 -192.000 ;
        RECT -109.915 -193.235 -109.745 -191.695 ;
        RECT -109.425 -193.235 -109.255 -191.695 ;
        RECT -108.935 -193.235 -108.765 -191.695 ;
        RECT -108.445 -193.235 -108.275 -191.695 ;
        RECT -107.955 -193.235 -107.785 -191.695 ;
        RECT -109.430 -193.495 -109.255 -193.235 ;
        RECT -105.860 -193.405 -105.555 -191.370 ;
        RECT -103.565 -192.010 -103.275 -191.325 ;
        RECT -102.495 -191.340 -102.205 -190.840 ;
        RECT -102.010 -190.870 -101.720 -190.415 ;
        RECT -99.755 -190.450 -99.080 -190.415 ;
        RECT -98.815 -190.635 -98.140 -190.570 ;
        RECT -101.520 -190.805 -98.140 -190.635 ;
        RECT -101.520 -191.340 -101.350 -190.805 ;
        RECT -98.815 -190.840 -98.140 -190.805 ;
        RECT -97.970 -190.630 -97.785 -189.940 ;
        RECT -95.760 -190.630 -95.085 -190.580 ;
        RECT -97.970 -190.815 -95.085 -190.630 ;
        RECT -97.970 -191.085 -97.785 -190.815 ;
        RECT -95.760 -190.850 -95.085 -190.815 ;
        RECT -94.910 -190.940 -94.740 -188.535 ;
        RECT -91.405 -190.460 -91.235 -189.420 ;
        RECT -90.425 -190.460 -90.255 -189.420 ;
        RECT -89.445 -190.460 -89.275 -189.420 ;
        RECT -86.540 -190.495 -86.370 -188.775 ;
        RECT -85.560 -190.495 -85.390 -188.775 ;
        RECT -83.495 -189.310 -83.325 -188.770 ;
        RECT -82.515 -189.310 -82.345 -188.770 ;
        RECT -84.085 -189.545 -83.720 -189.480 ;
        RECT -84.585 -189.685 -83.720 -189.545 ;
        RECT -84.695 -189.750 -83.720 -189.685 ;
        RECT -84.695 -190.495 -84.390 -189.750 ;
        RECT -84.085 -189.780 -83.720 -189.750 ;
        RECT -81.535 -189.630 -81.365 -188.770 ;
        RECT -80.025 -189.630 -79.675 -182.945 ;
        RECT -87.455 -190.560 -86.780 -190.530 ;
        RECT -87.555 -190.570 -86.780 -190.560 ;
        RECT -92.865 -190.695 -92.215 -190.610 ;
        RECT -91.995 -190.695 -91.630 -190.630 ;
        RECT -92.865 -190.900 -91.630 -190.695 ;
        RECT -88.590 -190.750 -86.780 -190.570 ;
        RECT -86.540 -190.645 -84.390 -190.495 ;
        RECT -86.540 -190.685 -84.445 -190.645 ;
        RECT -83.495 -190.705 -83.325 -189.925 ;
        RECT -83.005 -190.465 -82.835 -189.925 ;
        RECT -82.515 -190.705 -82.345 -189.925 ;
        RECT -82.025 -190.465 -81.855 -189.925 ;
        RECT -81.535 -189.980 -79.675 -189.630 ;
        RECT -87.555 -190.760 -86.780 -190.750 ;
        RECT -87.455 -190.800 -86.780 -190.760 ;
        RECT -92.865 -190.940 -92.215 -190.900 ;
        RECT -91.995 -190.930 -91.630 -190.900 ;
        RECT -102.495 -191.510 -101.350 -191.340 ;
        RECT -101.050 -191.255 -98.835 -191.085 ;
        RECT -97.970 -191.255 -96.805 -191.085 ;
        RECT -102.495 -191.525 -102.205 -191.510 ;
        RECT -101.050 -193.110 -100.880 -191.255 ;
        RECT -100.070 -191.260 -98.835 -191.255 ;
        RECT -102.685 -193.405 -102.110 -193.400 ;
        RECT -107.805 -193.495 -101.960 -193.405 ;
        RECT -130.080 -193.925 -128.040 -193.755 ;
        RECT -110.015 -193.800 -101.960 -193.495 ;
        RECT -107.810 -193.980 -101.960 -193.800 ;
        RECT -102.685 -194.070 -101.960 -193.980 ;
        RECT -100.560 -194.055 -100.390 -191.570 ;
        RECT -100.070 -193.110 -99.900 -191.260 ;
        RECT -99.010 -191.575 -98.835 -191.260 ;
        RECT -99.500 -193.070 -99.330 -191.575 ;
        RECT -99.500 -193.590 -99.325 -193.070 ;
        RECT -99.010 -193.115 -98.840 -191.575 ;
        RECT -98.520 -193.060 -98.350 -191.575 ;
        RECT -98.520 -193.590 -98.345 -193.060 ;
        RECT -97.955 -193.115 -97.785 -191.255 ;
        RECT -99.500 -193.605 -98.345 -193.590 ;
        RECT -97.465 -193.605 -97.295 -191.575 ;
        RECT -96.975 -193.115 -96.805 -191.255 ;
        RECT -94.910 -191.110 -92.215 -190.940 ;
        RECT -89.930 -191.050 -87.185 -191.040 ;
        RECT -85.130 -191.050 -84.760 -190.920 ;
        RECT -89.930 -191.070 -84.760 -191.050 ;
        RECT -99.500 -193.775 -97.295 -193.605 ;
        RECT -95.400 -193.920 -95.230 -192.075 ;
        RECT -94.910 -193.115 -94.740 -191.110 ;
        RECT -92.865 -191.360 -92.215 -191.110 ;
        RECT -91.405 -192.350 -91.235 -191.070 ;
        RECT -90.915 -192.110 -90.745 -191.070 ;
        RECT -90.425 -192.350 -90.255 -191.070 ;
        RECT -89.935 -191.240 -84.760 -191.070 ;
        RECT -84.195 -191.135 -80.270 -190.705 ;
        RECT -89.935 -192.110 -89.765 -191.240 ;
        RECT -87.190 -191.245 -84.760 -191.240 ;
        RECT -87.190 -191.250 -86.835 -191.245 ;
        RECT -85.130 -191.275 -84.760 -191.245 ;
        RECT -92.105 -192.780 -87.415 -192.350 ;
        RECT -87.845 -193.185 -87.415 -192.780 ;
        RECT -87.030 -193.000 -86.860 -191.460 ;
        RECT -86.540 -193.000 -86.370 -191.460 ;
        RECT -86.050 -193.000 -85.880 -191.460 ;
        RECT -85.560 -193.000 -85.390 -191.460 ;
        RECT -85.070 -193.000 -84.900 -191.460 ;
        RECT -86.545 -193.185 -86.370 -193.000 ;
        RECT -82.975 -193.170 -82.670 -191.135 ;
        RECT -84.920 -193.185 -82.670 -193.170 ;
        RECT -87.845 -193.475 -82.670 -193.185 ;
        RECT -87.845 -193.615 -84.520 -193.475 ;
        RECT -87.665 -193.920 -86.615 -193.615 ;
        RECT -96.405 -194.055 -86.615 -193.920 ;
        RECT -101.050 -194.070 -86.615 -194.055 ;
        RECT -135.145 -194.355 -132.080 -194.185 ;
        RECT -135.145 -195.365 -134.545 -194.355 ;
        RECT -102.685 -194.465 -86.615 -194.070 ;
        RECT -122.250 -194.695 -86.615 -194.465 ;
        RECT -82.005 -193.865 -80.665 -193.615 ;
        RECT -76.855 -193.865 -75.940 -182.070 ;
        RECT -72.205 -182.550 -72.035 -181.590 ;
        RECT -71.225 -182.550 -71.055 -181.590 ;
        RECT -70.275 -182.530 -70.045 -181.265 ;
        RECT -68.040 -181.585 -67.165 -181.160 ;
        RECT -65.245 -181.315 -64.385 -180.945 ;
        RECT -68.040 -181.755 -64.900 -181.585 ;
        RECT -68.040 -181.975 -67.830 -181.755 ;
        RECT -68.015 -182.475 -67.845 -181.975 ;
        RECT -67.525 -182.390 -67.355 -181.935 ;
        RECT -67.040 -182.025 -66.860 -181.755 ;
        RECT -66.070 -181.935 -65.890 -181.755 ;
        RECT -70.245 -182.550 -70.075 -182.530 ;
        RECT -67.550 -182.645 -67.340 -182.390 ;
        RECT -67.035 -182.475 -66.865 -182.025 ;
        RECT -66.545 -182.365 -66.375 -181.935 ;
        RECT -66.070 -182.025 -65.885 -181.935 ;
        RECT -66.570 -182.645 -66.360 -182.365 ;
        RECT -66.055 -182.475 -65.885 -182.025 ;
        RECT -65.565 -182.370 -65.395 -181.935 ;
        RECT -65.080 -182.015 -64.900 -181.755 ;
        RECT -65.600 -182.645 -65.390 -182.370 ;
        RECT -65.075 -182.475 -64.905 -182.015 ;
        RECT -64.620 -182.050 -64.385 -181.315 ;
        RECT -64.160 -181.035 -63.290 -180.875 ;
        RECT -62.540 -181.035 -62.310 -180.570 ;
        RECT -62.020 -180.650 -61.850 -179.855 ;
        RECT -61.530 -180.570 -61.360 -180.110 ;
        RECT -61.560 -181.035 -61.330 -180.570 ;
        RECT -61.040 -180.650 -60.870 -179.855 ;
        RECT -64.160 -181.225 -61.330 -181.035 ;
        RECT -61.150 -180.845 -60.310 -180.820 ;
        RECT -60.010 -180.845 -59.710 -180.480 ;
        RECT -61.150 -181.135 -59.710 -180.845 ;
        RECT -59.435 -180.930 -59.135 -180.355 ;
        RECT -58.705 -180.570 -58.535 -180.110 ;
        RECT -58.735 -180.875 -58.505 -180.570 ;
        RECT -58.215 -180.650 -58.045 -179.855 ;
        RECT -57.725 -180.570 -57.555 -180.110 ;
        RECT -58.885 -180.930 -58.505 -180.875 ;
        RECT -61.150 -181.190 -60.310 -181.135 ;
        RECT -60.010 -181.140 -59.710 -181.135 ;
        RECT -59.460 -181.035 -58.505 -180.930 ;
        RECT -57.755 -181.035 -57.525 -180.570 ;
        RECT -57.235 -180.650 -57.065 -179.855 ;
        RECT -56.745 -180.570 -56.575 -180.110 ;
        RECT -56.775 -181.035 -56.545 -180.570 ;
        RECT -56.255 -180.650 -56.085 -179.855 ;
        RECT -54.530 -180.330 -54.300 -179.720 ;
        RECT -54.055 -179.920 -53.835 -179.630 ;
        RECT -54.535 -180.380 -54.300 -180.330 ;
        RECT -54.535 -180.545 -54.330 -180.380 ;
        RECT -54.025 -180.400 -53.855 -179.920 ;
        RECT -53.535 -180.335 -53.365 -179.860 ;
        RECT -53.070 -179.975 -52.850 -179.630 ;
        RECT -54.540 -180.580 -54.330 -180.545 ;
        RECT -53.550 -180.580 -53.345 -180.335 ;
        RECT -53.045 -180.400 -52.875 -179.975 ;
        RECT -52.555 -180.335 -52.385 -179.860 ;
        RECT -52.090 -179.975 -51.870 -179.630 ;
        RECT -52.580 -180.580 -52.375 -180.335 ;
        RECT -52.065 -180.400 -51.895 -179.975 ;
        RECT -51.575 -180.375 -51.405 -179.860 ;
        RECT -51.110 -179.920 -50.890 -179.630 ;
        RECT -49.995 -179.855 -42.915 -179.515 ;
        RECT -51.085 -180.270 -50.915 -179.920 ;
        RECT -51.590 -180.580 -51.385 -180.375 ;
        RECT -54.540 -180.750 -51.385 -180.580 ;
        RECT -59.460 -181.155 -56.545 -181.035 ;
        RECT -64.160 -181.345 -63.795 -181.225 ;
        RECT -64.585 -182.420 -64.415 -182.050 ;
        RECT -64.165 -182.185 -63.795 -181.345 ;
        RECT -63.520 -181.265 -61.330 -181.225 ;
        RECT -63.520 -181.590 -63.290 -181.265 ;
        RECT -62.540 -181.590 -62.310 -181.265 ;
        RECT -64.590 -182.645 -64.410 -182.420 ;
        RECT -63.490 -182.550 -63.320 -181.590 ;
        RECT -62.510 -182.550 -62.340 -181.590 ;
        RECT -61.560 -182.530 -61.330 -181.265 ;
        RECT -60.540 -181.825 -60.255 -181.620 ;
        RECT -59.460 -181.825 -59.235 -181.155 ;
        RECT -58.885 -181.225 -56.545 -181.155 ;
        RECT -56.365 -180.860 -55.525 -180.820 ;
        RECT -54.540 -180.860 -53.665 -180.750 ;
        RECT -56.365 -181.145 -53.665 -180.860 ;
        RECT -51.120 -180.945 -50.885 -180.270 ;
        RECT -49.990 -180.570 -49.820 -180.110 ;
        RECT -50.020 -180.875 -49.790 -180.570 ;
        RECT -49.500 -180.650 -49.330 -179.855 ;
        RECT -49.010 -180.570 -48.840 -180.110 ;
        RECT -56.365 -181.190 -55.525 -181.145 ;
        RECT -58.735 -181.265 -56.545 -181.225 ;
        RECT -58.735 -181.590 -58.505 -181.265 ;
        RECT -57.755 -181.590 -57.525 -181.265 ;
        RECT -60.540 -182.050 -59.235 -181.825 ;
        RECT -60.540 -182.440 -60.255 -182.050 ;
        RECT -61.530 -182.550 -61.360 -182.530 ;
        RECT -58.705 -182.550 -58.535 -181.590 ;
        RECT -57.725 -182.550 -57.555 -181.590 ;
        RECT -56.775 -182.530 -56.545 -181.265 ;
        RECT -54.540 -181.585 -53.665 -181.145 ;
        RECT -51.745 -181.315 -50.885 -180.945 ;
        RECT -54.540 -181.755 -51.400 -181.585 ;
        RECT -54.540 -181.975 -54.330 -181.755 ;
        RECT -54.515 -182.475 -54.345 -181.975 ;
        RECT -54.025 -182.390 -53.855 -181.935 ;
        RECT -53.540 -182.025 -53.360 -181.755 ;
        RECT -52.570 -181.935 -52.390 -181.755 ;
        RECT -56.745 -182.550 -56.575 -182.530 ;
        RECT -67.550 -182.815 -64.410 -182.645 ;
        RECT -54.050 -182.645 -53.840 -182.390 ;
        RECT -53.535 -182.475 -53.365 -182.025 ;
        RECT -53.045 -182.365 -52.875 -181.935 ;
        RECT -52.570 -182.025 -52.385 -181.935 ;
        RECT -53.070 -182.645 -52.860 -182.365 ;
        RECT -52.555 -182.475 -52.385 -182.025 ;
        RECT -52.065 -182.370 -51.895 -181.935 ;
        RECT -51.580 -182.015 -51.400 -181.755 ;
        RECT -52.100 -182.645 -51.890 -182.370 ;
        RECT -51.575 -182.475 -51.405 -182.015 ;
        RECT -51.120 -182.050 -50.885 -181.315 ;
        RECT -50.660 -181.035 -49.790 -180.875 ;
        RECT -49.040 -181.035 -48.810 -180.570 ;
        RECT -48.520 -180.650 -48.350 -179.855 ;
        RECT -48.030 -180.570 -47.860 -180.110 ;
        RECT -48.060 -181.035 -47.830 -180.570 ;
        RECT -47.540 -180.650 -47.370 -179.855 ;
        RECT -50.660 -181.225 -47.830 -181.035 ;
        RECT -47.650 -180.845 -46.810 -180.820 ;
        RECT -47.650 -180.905 -46.635 -180.845 ;
        RECT -46.350 -180.905 -46.050 -180.475 ;
        RECT -45.580 -180.570 -45.410 -180.110 ;
        RECT -45.610 -180.875 -45.380 -180.570 ;
        RECT -45.090 -180.650 -44.920 -179.855 ;
        RECT -44.600 -180.570 -44.430 -180.110 ;
        RECT -45.760 -180.905 -45.380 -180.875 ;
        RECT -47.650 -181.035 -45.380 -180.905 ;
        RECT -44.630 -181.035 -44.400 -180.570 ;
        RECT -44.110 -180.650 -43.940 -179.855 ;
        RECT -43.620 -180.570 -43.450 -180.110 ;
        RECT -43.650 -181.035 -43.420 -180.570 ;
        RECT -43.130 -180.650 -42.960 -179.855 ;
        RECT -42.695 -180.820 -42.500 -179.375 ;
        RECT -40.500 -179.575 -40.280 -179.375 ;
        RECT -47.650 -181.115 -43.420 -181.035 ;
        RECT -47.650 -181.135 -46.635 -181.115 ;
        RECT -46.350 -181.135 -46.050 -181.115 ;
        RECT -47.650 -181.190 -46.810 -181.135 ;
        RECT -45.760 -181.225 -43.420 -181.115 ;
        RECT -43.240 -181.190 -42.400 -180.820 ;
        RECT -40.470 -181.070 -40.300 -179.575 ;
        RECT -39.980 -180.945 -39.810 -179.530 ;
        RECT -50.660 -181.345 -50.295 -181.225 ;
        RECT -51.085 -182.420 -50.915 -182.050 ;
        RECT -50.665 -182.185 -50.295 -181.345 ;
        RECT -50.020 -181.265 -47.830 -181.225 ;
        RECT -50.020 -181.590 -49.790 -181.265 ;
        RECT -49.040 -181.590 -48.810 -181.265 ;
        RECT -51.090 -182.645 -50.910 -182.420 ;
        RECT -49.990 -182.550 -49.820 -181.590 ;
        RECT -49.010 -182.550 -48.840 -181.590 ;
        RECT -48.060 -182.530 -47.830 -181.265 ;
        RECT -45.610 -181.265 -43.420 -181.225 ;
        RECT -45.610 -181.590 -45.380 -181.265 ;
        RECT -44.630 -181.590 -44.400 -181.265 ;
        RECT -47.040 -182.440 -46.755 -181.620 ;
        RECT -48.030 -182.550 -47.860 -182.530 ;
        RECT -45.580 -182.550 -45.410 -181.590 ;
        RECT -44.600 -182.550 -44.430 -181.590 ;
        RECT -43.650 -182.530 -43.420 -181.265 ;
        RECT -42.130 -181.595 -40.740 -181.590 ;
        RECT -40.010 -181.595 -39.775 -180.945 ;
        RECT -38.770 -180.995 -38.600 -179.530 ;
        RECT -38.305 -179.610 -38.080 -179.260 ;
        RECT -37.850 -179.130 -37.075 -179.085 ;
        RECT -37.850 -179.300 -35.040 -179.130 ;
        RECT -37.850 -179.360 -37.075 -179.300 ;
        RECT -38.800 -181.595 -38.565 -180.995 ;
        RECT -38.280 -181.070 -38.110 -179.610 ;
        RECT -37.790 -181.000 -37.620 -179.530 ;
        RECT -37.820 -181.595 -37.585 -181.000 ;
        RECT -42.130 -182.005 -37.175 -181.595 ;
        RECT -43.620 -182.550 -43.450 -182.530 ;
        RECT -54.050 -182.815 -50.910 -182.645 ;
        RECT -63.025 -184.520 -55.640 -183.955 ;
        RECT -67.180 -185.995 -64.935 -185.905 ;
        RECT -63.025 -185.995 -62.720 -184.520 ;
        RECT -59.390 -185.110 -59.155 -184.520 ;
        RECT -67.180 -186.210 -62.720 -185.995 ;
        RECT -66.595 -186.470 -66.420 -186.210 ;
        RECT -64.970 -186.300 -62.720 -186.210 ;
        RECT -67.080 -188.010 -66.910 -186.470 ;
        RECT -66.590 -188.010 -66.420 -186.470 ;
        RECT -66.100 -188.010 -65.930 -186.470 ;
        RECT -65.610 -188.010 -65.440 -186.470 ;
        RECT -65.120 -188.010 -64.950 -186.470 ;
        RECT -63.025 -188.335 -62.720 -186.300 ;
        RECT -59.355 -186.580 -59.185 -185.110 ;
        RECT -58.865 -186.500 -58.695 -185.040 ;
        RECT -58.410 -185.115 -58.175 -184.520 ;
        RECT -59.900 -186.810 -59.125 -186.750 ;
        RECT -60.085 -186.980 -59.125 -186.810 ;
        RECT -59.900 -187.025 -59.125 -186.980 ;
        RECT -58.895 -186.850 -58.670 -186.500 ;
        RECT -58.375 -186.580 -58.205 -185.115 ;
        RECT -57.200 -185.165 -56.965 -184.520 ;
        RECT -57.165 -186.580 -56.995 -185.165 ;
        RECT -56.675 -186.535 -56.505 -185.040 ;
        RECT -56.695 -186.735 -56.475 -186.535 ;
        RECT -56.695 -186.750 -41.295 -186.735 ;
        RECT -58.895 -187.050 -57.125 -186.850 ;
        RECT -56.935 -186.950 -41.295 -186.750 ;
        RECT -60.575 -187.335 -60.225 -187.325 ;
        RECT -58.550 -187.335 -57.775 -187.290 ;
        RECT -60.575 -187.515 -57.775 -187.335 ;
        RECT -69.805 -188.720 -68.875 -188.435 ;
        RECT -67.505 -188.710 -66.830 -188.670 ;
        RECT -67.605 -188.720 -66.830 -188.710 ;
        RECT -69.805 -188.900 -66.830 -188.720 ;
        RECT -64.245 -188.765 -61.170 -188.335 ;
        RECT -69.805 -189.205 -68.875 -188.900 ;
        RECT -67.605 -188.910 -66.830 -188.900 ;
        RECT -67.505 -188.940 -66.830 -188.910 ;
        RECT -66.590 -188.825 -64.495 -188.785 ;
        RECT -66.590 -188.975 -64.440 -188.825 ;
        RECT -66.590 -190.695 -66.420 -188.975 ;
        RECT -65.610 -190.695 -65.440 -188.975 ;
        RECT -64.745 -189.720 -64.440 -188.975 ;
        RECT -63.545 -189.545 -63.375 -188.765 ;
        RECT -63.055 -189.545 -62.885 -189.005 ;
        RECT -62.565 -189.545 -62.395 -188.765 ;
        RECT -62.075 -189.545 -61.905 -189.005 ;
        RECT -60.575 -189.490 -60.225 -187.515 ;
        RECT -58.550 -187.565 -57.775 -187.515 ;
        RECT -57.340 -187.400 -57.125 -187.050 ;
        RECT -57.340 -187.675 -56.435 -187.400 ;
        RECT -57.340 -187.735 -57.125 -187.675 ;
        RECT -59.375 -187.925 -58.105 -187.745 ;
        RECT -59.375 -188.220 -59.165 -187.925 ;
        RECT -58.315 -188.190 -58.105 -187.925 ;
        RECT -57.830 -187.930 -57.125 -187.735 ;
        RECT -64.135 -189.720 -63.770 -189.690 ;
        RECT -64.745 -189.785 -63.770 -189.720 ;
        RECT -64.635 -189.925 -63.770 -189.785 ;
        RECT -64.135 -189.990 -63.770 -189.925 ;
        RECT -61.585 -189.840 -60.195 -189.490 ;
        RECT -63.545 -190.700 -63.375 -190.160 ;
        RECT -62.565 -190.700 -62.395 -190.160 ;
        RECT -61.585 -190.700 -61.415 -189.840 ;
        RECT -59.355 -191.140 -59.185 -188.220 ;
        RECT -58.300 -191.100 -58.130 -188.190 ;
        RECT -57.830 -188.200 -57.620 -187.930 ;
        RECT -58.320 -191.310 -58.110 -191.100 ;
        RECT -57.810 -191.140 -57.640 -188.200 ;
        RECT -57.320 -191.090 -57.150 -188.100 ;
        RECT -56.265 -188.170 -56.050 -186.950 ;
        RECT -42.175 -187.345 -41.295 -186.950 ;
        RECT -55.135 -187.825 -54.610 -187.465 ;
        RECT -57.330 -191.310 -57.120 -191.090 ;
        RECT -56.260 -191.140 -56.090 -188.170 ;
        RECT -58.320 -191.480 -57.120 -191.310 ;
        RECT -130.080 -195.105 -128.040 -194.935 ;
        RECT -122.250 -195.040 -102.110 -194.695 ;
        RECT -82.005 -194.780 -75.940 -193.865 ;
        RECT -82.005 -194.940 -80.665 -194.780 ;
        RECT -135.145 -195.460 -132.080 -195.365 ;
        RECT -138.020 -195.535 -132.080 -195.460 ;
        RECT -138.020 -196.345 -134.545 -195.535 ;
        RECT -130.080 -196.285 -128.040 -196.115 ;
        RECT -138.020 -199.865 -137.320 -196.345 ;
        RECT -135.145 -196.545 -134.545 -196.345 ;
        RECT -135.145 -196.715 -132.080 -196.545 ;
        RECT -135.145 -197.725 -134.545 -196.715 ;
        RECT -130.080 -197.465 -128.040 -197.295 ;
        RECT -135.145 -197.895 -132.080 -197.725 ;
        RECT -135.145 -198.905 -134.545 -197.895 ;
        RECT -131.420 -198.285 -130.640 -197.925 ;
        RECT -134.120 -198.485 -132.080 -198.315 ;
        RECT -135.145 -199.075 -132.080 -198.905 ;
        RECT -135.145 -199.865 -134.545 -199.075 ;
        RECT -134.120 -199.665 -132.080 -199.495 ;
        RECT -138.020 -200.085 -134.545 -199.865 ;
        RECT -138.020 -200.255 -132.080 -200.085 ;
        RECT -138.020 -200.750 -134.545 -200.255 ;
        RECT -131.180 -200.305 -131.010 -198.285 ;
        RECT -130.080 -198.645 -128.040 -198.475 ;
        RECT -131.180 -200.475 -128.040 -200.305 ;
        RECT -138.020 -203.975 -137.320 -200.750 ;
        RECT -135.145 -201.265 -134.545 -200.750 ;
        RECT -134.120 -200.845 -132.080 -200.675 ;
        RECT -135.145 -201.435 -132.080 -201.265 ;
        RECT -135.145 -202.445 -134.545 -201.435 ;
        RECT -130.080 -201.655 -128.040 -201.485 ;
        RECT -134.120 -202.025 -132.080 -201.855 ;
        RECT -135.145 -202.615 -132.080 -202.445 ;
        RECT -135.145 -203.625 -134.545 -202.615 ;
        RECT -134.120 -203.205 -132.080 -203.035 ;
        RECT -131.485 -203.090 -130.785 -202.580 ;
        RECT -130.080 -202.835 -128.040 -202.665 ;
        RECT -135.145 -203.795 -132.080 -203.625 ;
        RECT -135.145 -203.975 -134.545 -203.795 ;
        RECT -138.020 -204.805 -134.545 -203.975 ;
        RECT -134.120 -204.385 -132.080 -204.215 ;
        RECT -131.195 -204.805 -131.025 -203.090 ;
        RECT -130.080 -204.015 -128.040 -203.845 ;
        RECT -138.020 -204.860 -132.080 -204.805 ;
        RECT -138.020 -205.920 -137.320 -204.860 ;
        RECT -135.145 -204.975 -132.080 -204.860 ;
        RECT -131.195 -204.975 -130.410 -204.805 ;
        RECT -135.145 -205.985 -134.545 -204.975 ;
        RECT -134.120 -205.565 -132.080 -205.395 ;
        RECT -131.760 -205.970 -130.875 -205.590 ;
        RECT -130.580 -205.675 -130.410 -204.975 ;
        RECT -130.580 -205.845 -128.040 -205.675 ;
        RECT -135.145 -206.155 -132.080 -205.985 ;
        RECT -135.145 -206.365 -134.545 -206.155 ;
        RECT -131.480 -207.005 -131.175 -205.970 ;
        RECT -131.940 -207.100 -131.010 -207.005 ;
        RECT -130.080 -207.025 -128.040 -206.855 ;
        RECT -131.940 -220.870 -130.975 -207.100 ;
        RECT -129.885 -214.360 -128.195 -213.945 ;
        RECT -122.250 -214.360 -121.675 -195.040 ;
        RECT -66.460 -195.340 -66.290 -194.300 ;
        RECT -65.480 -195.340 -65.310 -194.300 ;
        RECT -64.500 -195.340 -64.330 -194.300 ;
        RECT -61.595 -195.375 -61.425 -193.655 ;
        RECT -60.615 -195.375 -60.445 -193.655 ;
        RECT -58.550 -194.190 -58.380 -193.650 ;
        RECT -57.570 -194.190 -57.400 -193.650 ;
        RECT -59.140 -194.425 -58.775 -194.360 ;
        RECT -59.640 -194.565 -58.775 -194.425 ;
        RECT -59.750 -194.630 -58.775 -194.565 ;
        RECT -59.750 -195.375 -59.445 -194.630 ;
        RECT -59.140 -194.660 -58.775 -194.630 ;
        RECT -56.590 -194.510 -56.420 -193.650 ;
        RECT -55.080 -194.510 -54.730 -187.825 ;
        RECT -35.210 -190.595 -35.040 -179.300 ;
        RECT -34.290 -185.040 -34.120 -177.340 ;
        RECT -33.740 -178.010 -33.045 -177.740 ;
        RECT -31.090 -177.915 -30.920 -177.340 ;
        RECT -30.615 -177.535 -30.445 -175.775 ;
        RECT -30.265 -177.165 -30.095 -175.430 ;
        RECT -21.235 -175.430 -17.595 -175.260 ;
        RECT -29.365 -177.165 -29.195 -175.950 ;
        RECT -30.265 -177.335 -29.195 -177.165 ;
        RECT -28.385 -177.535 -28.215 -175.950 ;
        RECT -26.835 -176.915 -26.665 -175.950 ;
        RECT -25.290 -176.905 -25.120 -175.950 ;
        RECT -30.615 -177.705 -28.215 -177.535 ;
        RECT -27.950 -177.790 -27.255 -177.520 ;
        RECT -31.090 -178.085 -30.360 -177.915 ;
        RECT -33.745 -178.600 -32.090 -178.415 ;
        RECT -31.830 -178.530 -31.135 -178.260 ;
        RECT -30.530 -178.395 -30.360 -178.085 ;
        RECT -29.995 -178.160 -29.300 -177.890 ;
        RECT -30.530 -178.565 -27.725 -178.395 ;
        RECT -33.745 -179.015 -33.560 -178.600 ;
        RECT -32.275 -178.720 -32.090 -178.600 ;
        RECT -32.275 -178.905 -31.495 -178.720 ;
        RECT -33.735 -179.960 -33.565 -179.015 ;
        RECT -33.755 -180.575 -33.560 -179.960 ;
        RECT -33.245 -180.205 -33.075 -178.980 ;
        RECT -31.680 -179.010 -31.495 -178.905 ;
        RECT -31.665 -180.020 -31.495 -179.010 ;
        RECT -31.185 -179.025 -29.685 -178.830 ;
        RECT -31.175 -180.020 -31.005 -179.025 ;
        RECT -29.855 -180.020 -29.685 -179.025 ;
        RECT -29.365 -180.020 -29.195 -178.565 ;
        RECT -28.385 -179.935 -28.215 -178.980 ;
        RECT -28.385 -180.205 -28.205 -179.935 ;
        RECT -27.895 -180.020 -27.725 -178.565 ;
        RECT -26.860 -178.610 -26.645 -176.915 ;
        RECT -25.310 -177.890 -25.095 -176.905 ;
        RECT -21.235 -176.990 -21.065 -175.430 ;
        RECT -20.745 -177.170 -20.575 -175.950 ;
        RECT -20.255 -176.990 -20.085 -175.430 ;
        RECT -19.655 -175.775 -17.945 -175.605 ;
        RECT -19.655 -176.990 -19.485 -175.775 ;
        RECT -19.165 -177.170 -18.995 -175.950 ;
        RECT -18.675 -176.990 -18.505 -175.775 ;
        RECT -22.075 -177.340 -18.420 -177.170 ;
        RECT -24.875 -177.820 -24.180 -177.550 ;
        RECT -25.810 -178.120 -25.095 -177.890 ;
        RECT -26.440 -178.560 -25.745 -178.290 ;
        RECT -27.340 -178.840 -26.645 -178.610 ;
        RECT -26.860 -179.065 -26.645 -178.840 ;
        RECT -26.835 -180.020 -26.665 -179.065 ;
        RECT -26.345 -179.985 -26.175 -178.980 ;
        RECT -25.310 -179.075 -25.095 -178.120 ;
        RECT -33.245 -180.385 -28.205 -180.205 ;
        RECT -26.370 -180.405 -26.155 -179.985 ;
        RECT -25.290 -180.020 -25.120 -179.075 ;
        RECT -24.800 -179.975 -24.630 -178.980 ;
        RECT -22.075 -179.155 -21.905 -177.340 ;
        RECT -21.240 -178.010 -20.545 -177.740 ;
        RECT -18.590 -177.915 -18.420 -177.340 ;
        RECT -18.115 -177.535 -17.945 -175.775 ;
        RECT -17.765 -177.165 -17.595 -175.430 ;
        RECT -8.735 -175.430 -5.095 -175.260 ;
        RECT -16.865 -177.165 -16.695 -175.950 ;
        RECT -17.765 -177.335 -16.695 -177.165 ;
        RECT -15.885 -177.535 -15.715 -175.950 ;
        RECT -14.335 -176.915 -14.165 -175.950 ;
        RECT -12.790 -176.905 -12.620 -175.950 ;
        RECT -18.115 -177.705 -15.715 -177.535 ;
        RECT -15.450 -177.790 -14.755 -177.520 ;
        RECT -18.590 -178.085 -17.860 -177.915 ;
        RECT -21.245 -178.600 -19.590 -178.415 ;
        RECT -19.330 -178.530 -18.635 -178.260 ;
        RECT -18.030 -178.395 -17.860 -178.085 ;
        RECT -17.495 -178.160 -16.800 -177.890 ;
        RECT -18.030 -178.565 -15.225 -178.395 ;
        RECT -21.245 -179.015 -21.060 -178.600 ;
        RECT -19.775 -178.720 -19.590 -178.600 ;
        RECT -19.775 -178.905 -18.995 -178.720 ;
        RECT -22.105 -179.835 -21.875 -179.155 ;
        RECT -21.235 -179.960 -21.065 -179.015 ;
        RECT -24.825 -180.400 -24.610 -179.975 ;
        RECT -21.255 -180.400 -21.060 -179.960 ;
        RECT -20.745 -180.205 -20.575 -178.980 ;
        RECT -19.180 -179.010 -18.995 -178.905 ;
        RECT -19.165 -180.020 -18.995 -179.010 ;
        RECT -18.685 -179.025 -17.185 -178.830 ;
        RECT -18.675 -180.020 -18.505 -179.025 ;
        RECT -17.355 -180.020 -17.185 -179.025 ;
        RECT -16.865 -180.020 -16.695 -178.565 ;
        RECT -15.885 -179.935 -15.715 -178.980 ;
        RECT -15.885 -180.205 -15.705 -179.935 ;
        RECT -15.395 -180.020 -15.225 -178.565 ;
        RECT -14.360 -178.610 -14.145 -176.915 ;
        RECT -12.810 -177.890 -12.595 -176.905 ;
        RECT -8.735 -176.990 -8.565 -175.430 ;
        RECT -8.245 -177.170 -8.075 -175.950 ;
        RECT -7.755 -176.990 -7.585 -175.430 ;
        RECT -7.155 -175.775 -5.445 -175.605 ;
        RECT -7.155 -176.990 -6.985 -175.775 ;
        RECT -6.665 -177.170 -6.495 -175.950 ;
        RECT -6.175 -176.990 -6.005 -175.775 ;
        RECT -9.335 -177.340 -5.920 -177.170 ;
        RECT -12.375 -177.820 -11.680 -177.550 ;
        RECT -13.310 -178.120 -12.595 -177.890 ;
        RECT -13.940 -178.560 -13.245 -178.290 ;
        RECT -14.840 -178.840 -14.145 -178.610 ;
        RECT -14.360 -179.065 -14.145 -178.840 ;
        RECT -14.335 -180.020 -14.165 -179.065 ;
        RECT -13.845 -179.985 -13.675 -178.980 ;
        RECT -12.810 -179.075 -12.595 -178.120 ;
        RECT -20.745 -180.385 -15.705 -180.205 ;
        RECT -25.195 -180.405 -21.060 -180.400 ;
        RECT -13.870 -180.405 -13.655 -179.985 ;
        RECT -12.790 -180.020 -12.620 -179.075 ;
        RECT -12.300 -179.975 -12.130 -178.980 ;
        RECT -9.335 -179.175 -9.165 -177.340 ;
        RECT -8.740 -178.010 -8.045 -177.740 ;
        RECT -6.090 -177.915 -5.920 -177.340 ;
        RECT -5.615 -177.535 -5.445 -175.775 ;
        RECT -5.265 -177.165 -5.095 -175.430 ;
        RECT 3.765 -175.430 7.405 -175.260 ;
        RECT -4.365 -177.165 -4.195 -175.950 ;
        RECT -5.265 -177.335 -4.195 -177.165 ;
        RECT -3.385 -177.535 -3.215 -175.950 ;
        RECT -1.835 -176.915 -1.665 -175.950 ;
        RECT -0.290 -176.905 -0.120 -175.950 ;
        RECT -5.615 -177.705 -3.215 -177.535 ;
        RECT -2.950 -177.790 -2.255 -177.520 ;
        RECT -6.090 -178.085 -5.360 -177.915 ;
        RECT -8.745 -178.600 -7.090 -178.415 ;
        RECT -6.830 -178.530 -6.135 -178.260 ;
        RECT -5.530 -178.395 -5.360 -178.085 ;
        RECT -4.995 -178.160 -4.300 -177.890 ;
        RECT -5.530 -178.565 -2.725 -178.395 ;
        RECT -8.745 -179.015 -8.560 -178.600 ;
        RECT -7.275 -178.720 -7.090 -178.600 ;
        RECT -7.275 -178.905 -6.495 -178.720 ;
        RECT -9.365 -179.855 -9.135 -179.175 ;
        RECT -8.735 -179.960 -8.565 -179.015 ;
        RECT -12.325 -180.405 -12.110 -179.975 ;
        RECT -27.750 -180.575 -21.060 -180.405 ;
        RECT -15.250 -180.575 -12.090 -180.405 ;
        RECT -8.755 -180.575 -8.560 -179.960 ;
        RECT -8.245 -180.205 -8.075 -178.980 ;
        RECT -6.680 -179.010 -6.495 -178.905 ;
        RECT -6.665 -180.020 -6.495 -179.010 ;
        RECT -6.185 -179.025 -4.685 -178.830 ;
        RECT -6.175 -180.020 -6.005 -179.025 ;
        RECT -4.855 -180.020 -4.685 -179.025 ;
        RECT -4.365 -180.020 -4.195 -178.565 ;
        RECT -3.385 -179.935 -3.215 -178.980 ;
        RECT -3.385 -180.205 -3.205 -179.935 ;
        RECT -2.895 -180.020 -2.725 -178.565 ;
        RECT -1.860 -178.610 -1.645 -176.915 ;
        RECT -0.310 -177.890 -0.095 -176.905 ;
        RECT 3.765 -176.990 3.935 -175.430 ;
        RECT 3.065 -177.170 3.235 -177.165 ;
        RECT 4.255 -177.170 4.425 -175.950 ;
        RECT 4.745 -176.990 4.915 -175.430 ;
        RECT 5.345 -175.775 7.055 -175.605 ;
        RECT 5.345 -176.990 5.515 -175.775 ;
        RECT 5.835 -177.170 6.005 -175.950 ;
        RECT 6.325 -176.990 6.495 -175.775 ;
        RECT 3.065 -177.340 6.580 -177.170 ;
        RECT 0.125 -177.820 0.820 -177.550 ;
        RECT -0.810 -178.120 -0.095 -177.890 ;
        RECT -1.440 -178.560 -0.745 -178.290 ;
        RECT -2.340 -178.840 -1.645 -178.610 ;
        RECT -1.860 -179.065 -1.645 -178.840 ;
        RECT -1.835 -180.020 -1.665 -179.065 ;
        RECT -1.345 -179.985 -1.175 -178.980 ;
        RECT -0.310 -179.075 -0.095 -178.120 ;
        RECT -8.245 -180.385 -3.205 -180.205 ;
        RECT -1.370 -180.405 -1.155 -179.985 ;
        RECT -0.290 -180.020 -0.120 -179.075 ;
        RECT 0.200 -179.975 0.370 -178.980 ;
        RECT 3.065 -179.175 3.235 -177.340 ;
        RECT 3.760 -178.010 4.455 -177.740 ;
        RECT 6.410 -177.915 6.580 -177.340 ;
        RECT 6.885 -177.535 7.055 -175.775 ;
        RECT 7.235 -177.165 7.405 -175.430 ;
        RECT 16.265 -175.430 19.905 -175.260 ;
        RECT 8.135 -177.165 8.305 -175.950 ;
        RECT 7.235 -177.335 8.305 -177.165 ;
        RECT 9.115 -177.535 9.285 -175.950 ;
        RECT 10.665 -176.915 10.835 -175.950 ;
        RECT 12.210 -176.905 12.380 -175.950 ;
        RECT 6.885 -177.705 9.285 -177.535 ;
        RECT 9.550 -177.790 10.245 -177.520 ;
        RECT 6.410 -178.085 7.140 -177.915 ;
        RECT 3.755 -178.600 5.410 -178.415 ;
        RECT 5.670 -178.530 6.365 -178.260 ;
        RECT 6.970 -178.395 7.140 -178.085 ;
        RECT 7.505 -178.160 8.200 -177.890 ;
        RECT 6.970 -178.565 9.775 -178.395 ;
        RECT 3.755 -179.015 3.940 -178.600 ;
        RECT 5.225 -178.720 5.410 -178.600 ;
        RECT 5.225 -178.905 6.005 -178.720 ;
        RECT 3.035 -179.855 3.265 -179.175 ;
        RECT 3.765 -179.960 3.935 -179.015 ;
        RECT 0.175 -180.405 0.390 -179.975 ;
        RECT -2.750 -180.575 0.410 -180.405 ;
        RECT 3.745 -180.575 3.940 -179.960 ;
        RECT 4.255 -180.205 4.425 -178.980 ;
        RECT 5.820 -179.010 6.005 -178.905 ;
        RECT 5.835 -180.020 6.005 -179.010 ;
        RECT 6.315 -179.025 7.815 -178.830 ;
        RECT 6.325 -180.020 6.495 -179.025 ;
        RECT 7.645 -180.020 7.815 -179.025 ;
        RECT 8.135 -180.020 8.305 -178.565 ;
        RECT 9.115 -179.935 9.285 -178.980 ;
        RECT 9.115 -180.205 9.295 -179.935 ;
        RECT 9.605 -180.020 9.775 -178.565 ;
        RECT 10.640 -178.610 10.855 -176.915 ;
        RECT 12.190 -177.890 12.405 -176.905 ;
        RECT 16.265 -176.990 16.435 -175.430 ;
        RECT 16.755 -177.170 16.925 -175.950 ;
        RECT 17.245 -176.990 17.415 -175.430 ;
        RECT 17.845 -175.775 19.555 -175.605 ;
        RECT 17.845 -176.990 18.015 -175.775 ;
        RECT 18.335 -177.170 18.505 -175.950 ;
        RECT 18.825 -176.990 18.995 -175.775 ;
        RECT 15.145 -177.340 19.080 -177.170 ;
        RECT 12.625 -177.820 13.320 -177.550 ;
        RECT 11.690 -178.120 12.405 -177.890 ;
        RECT 11.060 -178.560 11.755 -178.290 ;
        RECT 10.160 -178.840 10.855 -178.610 ;
        RECT 10.640 -179.065 10.855 -178.840 ;
        RECT 10.665 -180.020 10.835 -179.065 ;
        RECT 11.155 -179.985 11.325 -178.980 ;
        RECT 12.190 -179.075 12.405 -178.120 ;
        RECT 4.255 -180.385 9.295 -180.205 ;
        RECT 11.130 -180.405 11.345 -179.985 ;
        RECT 12.210 -180.020 12.380 -179.075 ;
        RECT 12.700 -179.975 12.870 -178.980 ;
        RECT 15.145 -179.170 15.315 -177.340 ;
        RECT 16.260 -178.010 16.955 -177.740 ;
        RECT 18.910 -177.915 19.080 -177.340 ;
        RECT 19.385 -177.535 19.555 -175.775 ;
        RECT 19.735 -177.165 19.905 -175.430 ;
        RECT 31.265 -175.430 34.905 -175.260 ;
        RECT 20.635 -177.165 20.805 -175.950 ;
        RECT 19.735 -177.335 20.805 -177.165 ;
        RECT 21.615 -177.535 21.785 -175.950 ;
        RECT 23.165 -176.915 23.335 -175.950 ;
        RECT 24.710 -176.905 24.880 -175.950 ;
        RECT 19.385 -177.705 21.785 -177.535 ;
        RECT 22.050 -177.790 22.745 -177.520 ;
        RECT 18.910 -178.085 19.640 -177.915 ;
        RECT 19.470 -178.395 19.640 -178.085 ;
        RECT 20.005 -178.160 20.700 -177.890 ;
        RECT 16.255 -178.600 17.910 -178.415 ;
        RECT 19.470 -178.565 22.275 -178.395 ;
        RECT 16.255 -179.015 16.440 -178.600 ;
        RECT 17.725 -178.720 17.910 -178.600 ;
        RECT 17.725 -178.905 18.505 -178.720 ;
        RECT 15.145 -179.175 15.320 -179.170 ;
        RECT 15.120 -179.855 15.350 -179.175 ;
        RECT 16.265 -179.960 16.435 -179.015 ;
        RECT 12.675 -180.405 12.890 -179.975 ;
        RECT 9.750 -180.575 12.910 -180.405 ;
        RECT 16.245 -180.575 16.440 -179.960 ;
        RECT 16.755 -180.205 16.925 -178.980 ;
        RECT 18.320 -179.010 18.505 -178.905 ;
        RECT 18.335 -180.020 18.505 -179.010 ;
        RECT 18.815 -179.025 20.315 -178.830 ;
        RECT 18.825 -180.020 18.995 -179.025 ;
        RECT 20.145 -180.020 20.315 -179.025 ;
        RECT 20.635 -180.020 20.805 -178.565 ;
        RECT 21.615 -179.935 21.785 -178.980 ;
        RECT 21.615 -180.205 21.795 -179.935 ;
        RECT 22.105 -180.020 22.275 -178.565 ;
        RECT 23.140 -178.610 23.355 -176.915 ;
        RECT 24.690 -177.890 24.905 -176.905 ;
        RECT 31.265 -176.990 31.435 -175.430 ;
        RECT 31.755 -177.170 31.925 -175.950 ;
        RECT 32.245 -176.990 32.415 -175.430 ;
        RECT 32.845 -175.775 34.555 -175.605 ;
        RECT 32.845 -176.990 33.015 -175.775 ;
        RECT 33.335 -177.170 33.505 -175.950 ;
        RECT 33.825 -176.990 33.995 -175.775 ;
        RECT 29.675 -177.340 34.080 -177.170 ;
        RECT 25.125 -177.820 25.820 -177.550 ;
        RECT 24.190 -178.120 24.905 -177.890 ;
        RECT 22.660 -178.840 23.355 -178.610 ;
        RECT 23.140 -179.065 23.355 -178.840 ;
        RECT 23.165 -180.020 23.335 -179.065 ;
        RECT 23.655 -179.985 23.825 -178.980 ;
        RECT 24.690 -179.075 24.905 -178.120 ;
        RECT 16.755 -180.385 21.795 -180.205 ;
        RECT 23.630 -180.405 23.845 -179.985 ;
        RECT 24.710 -180.020 24.880 -179.075 ;
        RECT 25.200 -179.975 25.370 -178.980 ;
        RECT 29.675 -179.175 29.845 -177.340 ;
        RECT 31.260 -178.010 31.955 -177.740 ;
        RECT 33.910 -177.915 34.080 -177.340 ;
        RECT 34.385 -177.535 34.555 -175.775 ;
        RECT 34.735 -177.165 34.905 -175.430 ;
        RECT 35.635 -177.165 35.805 -175.950 ;
        RECT 34.735 -177.335 35.805 -177.165 ;
        RECT 36.615 -177.535 36.785 -175.950 ;
        RECT 38.165 -176.915 38.335 -175.950 ;
        RECT 39.710 -176.905 39.880 -175.950 ;
        RECT 34.385 -177.705 36.785 -177.535 ;
        RECT 37.050 -177.790 37.745 -177.520 ;
        RECT 33.910 -178.085 34.640 -177.915 ;
        RECT 34.470 -178.395 34.640 -178.085 ;
        RECT 35.005 -178.160 35.700 -177.890 ;
        RECT 31.255 -178.600 32.910 -178.415 ;
        RECT 34.470 -178.565 37.275 -178.395 ;
        RECT 31.255 -179.015 31.440 -178.600 ;
        RECT 32.725 -178.720 32.910 -178.600 ;
        RECT 32.725 -178.905 33.505 -178.720 ;
        RECT 29.645 -179.855 29.875 -179.175 ;
        RECT 31.265 -179.960 31.435 -179.015 ;
        RECT 25.175 -180.405 25.390 -179.975 ;
        RECT 22.250 -180.575 25.410 -180.405 ;
        RECT 31.245 -180.575 31.440 -179.960 ;
        RECT 31.755 -180.205 31.925 -178.980 ;
        RECT 33.320 -179.010 33.505 -178.905 ;
        RECT 33.335 -180.020 33.505 -179.010 ;
        RECT 33.815 -179.025 35.315 -178.830 ;
        RECT 33.825 -180.020 33.995 -179.025 ;
        RECT 35.145 -180.020 35.315 -179.025 ;
        RECT 35.635 -180.020 35.805 -178.565 ;
        RECT 36.615 -179.935 36.785 -178.980 ;
        RECT 36.615 -180.205 36.795 -179.935 ;
        RECT 37.105 -180.020 37.275 -178.565 ;
        RECT 38.140 -178.610 38.355 -176.915 ;
        RECT 39.690 -177.890 39.905 -176.905 ;
        RECT 40.125 -177.820 40.820 -177.550 ;
        RECT 39.190 -178.120 39.905 -177.890 ;
        RECT 37.660 -178.840 38.355 -178.610 ;
        RECT 38.140 -179.065 38.355 -178.840 ;
        RECT 38.165 -180.020 38.335 -179.065 ;
        RECT 38.655 -179.985 38.825 -178.980 ;
        RECT 39.690 -179.075 39.905 -178.120 ;
        RECT 31.755 -180.385 36.795 -180.205 ;
        RECT 38.630 -180.315 38.845 -179.985 ;
        RECT 39.710 -180.020 39.880 -179.075 ;
        RECT 40.200 -179.975 40.370 -178.980 ;
        RECT 40.175 -180.315 40.390 -179.975 ;
        RECT 41.205 -180.315 42.510 -171.010 ;
        RECT 84.280 -172.630 85.265 -171.725 ;
        RECT 82.560 -175.005 83.965 -173.960 ;
        RECT 43.630 -176.020 44.630 -175.850 ;
        RECT 80.760 -176.020 82.570 -175.790 ;
        RECT 43.630 -176.880 82.570 -176.020 ;
        RECT 43.630 -177.705 44.630 -176.880 ;
        RECT 80.760 -177.145 82.570 -176.880 ;
        RECT 37.170 -180.575 42.510 -180.315 ;
        RECT 79.560 -180.510 81.020 -180.505 ;
        RECT -33.755 -180.835 42.510 -180.575 ;
        RECT -33.755 -180.840 -24.590 -180.835 ;
        RECT -21.255 -180.840 42.510 -180.835 ;
        RECT -31.595 -180.940 -28.925 -180.840 ;
        RECT -27.750 -180.885 -24.590 -180.840 ;
        RECT -15.250 -180.885 -12.090 -180.840 ;
        RECT -2.750 -180.885 0.410 -180.840 ;
        RECT 9.750 -180.885 12.910 -180.840 ;
        RECT 22.250 -180.885 25.410 -180.840 ;
        RECT -31.550 -181.735 -31.380 -180.940 ;
        RECT -31.060 -181.655 -30.890 -181.195 ;
        RECT -31.090 -182.120 -30.860 -181.655 ;
        RECT -30.570 -181.735 -30.400 -180.940 ;
        RECT -30.080 -181.655 -29.910 -181.195 ;
        RECT -30.110 -182.120 -29.880 -181.655 ;
        RECT -29.590 -181.735 -29.420 -180.940 ;
        RECT 37.170 -180.950 42.510 -180.840 ;
        RECT -29.100 -181.655 -28.930 -181.195 ;
        RECT -8.540 -181.265 -7.860 -181.035 ;
        RECT 3.945 -181.115 4.625 -181.100 ;
        RECT -8.105 -181.505 -7.860 -181.265 ;
        RECT 3.780 -181.285 14.635 -181.115 ;
        RECT 3.945 -181.330 4.625 -181.285 ;
        RECT -29.130 -181.960 -28.900 -181.655 ;
        RECT -24.015 -181.960 -23.785 -181.630 ;
        RECT -8.105 -181.685 14.155 -181.505 ;
        RECT -29.130 -182.120 -23.785 -181.960 ;
        RECT -31.090 -182.310 -23.785 -182.120 ;
        RECT 13.975 -182.245 14.155 -181.685 ;
        RECT 14.465 -181.905 14.635 -181.285 ;
        RECT 29.385 -181.365 30.065 -181.335 ;
        RECT 14.860 -181.460 15.540 -181.415 ;
        RECT 14.860 -181.630 28.865 -181.460 ;
        RECT 29.385 -181.535 30.745 -181.365 ;
        RECT 29.385 -181.565 30.065 -181.535 ;
        RECT 14.860 -181.645 15.540 -181.630 ;
        RECT 28.695 -181.825 28.865 -181.630 ;
        RECT 14.465 -182.075 21.975 -181.905 ;
        RECT 28.695 -181.995 30.395 -181.825 ;
        RECT -31.090 -182.350 -28.900 -182.310 ;
        RECT -31.090 -183.615 -30.860 -182.350 ;
        RECT -30.110 -182.675 -29.880 -182.350 ;
        RECT -29.130 -182.675 -28.900 -182.350 ;
        RECT 13.975 -182.425 21.580 -182.245 ;
        RECT -31.060 -183.635 -30.890 -183.615 ;
        RECT -30.080 -183.635 -29.910 -182.675 ;
        RECT -29.100 -183.635 -28.930 -182.675 ;
        RECT -22.105 -183.365 -21.875 -182.685 ;
        RECT -22.090 -184.630 -21.890 -183.365 ;
        RECT -22.090 -184.860 -21.410 -184.630 ;
        RECT 13.155 -184.850 13.835 -184.620 ;
        RECT -34.490 -185.270 -33.810 -185.040 ;
        RECT 12.635 -185.270 13.410 -185.040 ;
        RECT -28.180 -187.015 -25.040 -186.845 ;
        RECT -32.835 -188.070 -32.665 -187.110 ;
        RECT -31.855 -188.070 -31.685 -187.110 ;
        RECT -30.875 -187.130 -30.705 -187.110 ;
        RECT -32.865 -188.395 -32.635 -188.070 ;
        RECT -31.885 -188.395 -31.655 -188.070 ;
        RECT -30.905 -188.395 -30.675 -187.130 ;
        RECT -28.645 -187.685 -28.475 -187.185 ;
        RECT -28.180 -187.270 -27.970 -187.015 ;
        RECT -32.865 -188.435 -30.675 -188.395 ;
        RECT -33.015 -188.480 -30.675 -188.435 ;
        RECT -28.670 -187.905 -28.460 -187.685 ;
        RECT -28.155 -187.725 -27.985 -187.270 ;
        RECT -27.665 -187.635 -27.495 -187.185 ;
        RECT -27.200 -187.295 -26.990 -187.015 ;
        RECT -27.670 -187.905 -27.490 -187.635 ;
        RECT -27.175 -187.725 -27.005 -187.295 ;
        RECT -26.685 -187.635 -26.515 -187.185 ;
        RECT -26.230 -187.290 -26.020 -187.015 ;
        RECT -26.700 -187.725 -26.515 -187.635 ;
        RECT -26.195 -187.725 -26.025 -187.290 ;
        RECT -25.705 -187.645 -25.535 -187.185 ;
        RECT -25.220 -187.240 -25.040 -187.015 ;
        RECT -14.680 -187.015 -11.540 -186.845 ;
        RECT -25.215 -187.610 -25.045 -187.240 ;
        RECT -26.700 -187.905 -26.520 -187.725 ;
        RECT -25.710 -187.905 -25.530 -187.645 ;
        RECT -28.670 -188.075 -25.530 -187.905 ;
        RECT -33.425 -188.490 -30.675 -188.480 ;
        RECT -33.430 -188.625 -30.675 -188.490 ;
        RECT -33.430 -188.675 -32.635 -188.625 ;
        RECT -33.430 -190.465 -33.190 -188.675 ;
        RECT -33.015 -188.785 -32.635 -188.675 ;
        RECT -32.865 -189.090 -32.635 -188.785 ;
        RECT -32.835 -189.550 -32.665 -189.090 ;
        RECT -32.345 -189.805 -32.175 -189.010 ;
        RECT -31.885 -189.090 -31.655 -188.625 ;
        RECT -31.855 -189.550 -31.685 -189.090 ;
        RECT -31.365 -189.805 -31.195 -189.010 ;
        RECT -30.905 -189.090 -30.675 -188.625 ;
        RECT -30.495 -188.500 -29.655 -188.470 ;
        RECT -28.670 -188.500 -27.795 -188.075 ;
        RECT -25.250 -188.345 -25.015 -187.610 ;
        RECT -24.795 -188.315 -24.425 -187.475 ;
        RECT -24.120 -188.070 -23.950 -187.110 ;
        RECT -23.140 -188.070 -22.970 -187.110 ;
        RECT -22.160 -187.130 -21.990 -187.110 ;
        RECT -30.495 -188.765 -27.795 -188.500 ;
        RECT -25.875 -188.715 -25.015 -188.345 ;
        RECT -30.495 -188.840 -29.655 -188.765 ;
        RECT -28.670 -188.910 -27.795 -188.765 ;
        RECT -30.875 -189.550 -30.705 -189.090 ;
        RECT -30.385 -189.805 -30.215 -189.010 ;
        RECT -28.670 -189.080 -25.515 -188.910 ;
        RECT -28.670 -189.115 -28.460 -189.080 ;
        RECT -28.665 -189.330 -28.460 -189.115 ;
        RECT -28.645 -189.800 -28.475 -189.330 ;
        RECT -28.155 -189.740 -27.985 -189.260 ;
        RECT -27.680 -189.325 -27.475 -189.080 ;
        RECT -32.840 -190.145 -30.170 -189.805 ;
        RECT -28.185 -190.030 -27.965 -189.740 ;
        RECT -27.665 -189.800 -27.495 -189.325 ;
        RECT -27.175 -189.685 -27.005 -189.260 ;
        RECT -26.710 -189.325 -26.505 -189.080 ;
        RECT -27.200 -190.030 -26.980 -189.685 ;
        RECT -26.685 -189.800 -26.515 -189.325 ;
        RECT -26.195 -189.685 -26.025 -189.260 ;
        RECT -25.720 -189.285 -25.515 -189.080 ;
        RECT -26.220 -190.030 -26.000 -189.685 ;
        RECT -25.705 -189.800 -25.535 -189.285 ;
        RECT -25.250 -189.390 -25.015 -188.715 ;
        RECT -24.790 -188.435 -24.425 -188.315 ;
        RECT -24.150 -188.395 -23.920 -188.070 ;
        RECT -23.170 -188.395 -22.940 -188.070 ;
        RECT -22.190 -188.395 -21.960 -187.130 ;
        RECT -21.170 -187.610 -20.885 -187.220 ;
        RECT -21.170 -187.835 -19.865 -187.610 ;
        RECT -21.170 -188.040 -20.885 -187.835 ;
        RECT -24.150 -188.435 -21.960 -188.395 ;
        RECT -24.790 -188.625 -21.960 -188.435 ;
        RECT -24.790 -188.785 -23.920 -188.625 ;
        RECT -24.150 -189.090 -23.920 -188.785 ;
        RECT -25.215 -189.740 -25.045 -189.390 ;
        RECT -24.120 -189.550 -23.950 -189.090 ;
        RECT -25.240 -190.030 -25.020 -189.740 ;
        RECT -23.630 -189.805 -23.460 -189.010 ;
        RECT -23.170 -189.090 -22.940 -188.625 ;
        RECT -23.140 -189.550 -22.970 -189.090 ;
        RECT -22.650 -189.805 -22.480 -189.010 ;
        RECT -22.190 -189.090 -21.960 -188.625 ;
        RECT -21.780 -188.525 -20.940 -188.470 ;
        RECT -20.090 -188.505 -19.865 -187.835 ;
        RECT -19.335 -188.070 -19.165 -187.110 ;
        RECT -18.355 -188.070 -18.185 -187.110 ;
        RECT -17.375 -187.130 -17.205 -187.110 ;
        RECT -19.365 -188.395 -19.135 -188.070 ;
        RECT -18.385 -188.395 -18.155 -188.070 ;
        RECT -17.405 -188.395 -17.175 -187.130 ;
        RECT -15.145 -187.685 -14.975 -187.185 ;
        RECT -14.680 -187.270 -14.470 -187.015 ;
        RECT -19.365 -188.435 -17.175 -188.395 ;
        RECT -19.515 -188.505 -17.175 -188.435 ;
        RECT -15.170 -187.905 -14.960 -187.685 ;
        RECT -14.655 -187.725 -14.485 -187.270 ;
        RECT -14.165 -187.635 -13.995 -187.185 ;
        RECT -13.700 -187.295 -13.490 -187.015 ;
        RECT -14.170 -187.905 -13.990 -187.635 ;
        RECT -13.675 -187.725 -13.505 -187.295 ;
        RECT -13.185 -187.635 -13.015 -187.185 ;
        RECT -12.730 -187.290 -12.520 -187.015 ;
        RECT -13.200 -187.725 -13.015 -187.635 ;
        RECT -12.695 -187.725 -12.525 -187.290 ;
        RECT -12.205 -187.645 -12.035 -187.185 ;
        RECT -11.720 -187.240 -11.540 -187.015 ;
        RECT -11.715 -187.610 -11.545 -187.240 ;
        RECT -13.200 -187.905 -13.020 -187.725 ;
        RECT -12.210 -187.905 -12.030 -187.645 ;
        RECT -15.170 -188.075 -12.030 -187.905 ;
        RECT -20.640 -188.525 -20.340 -188.520 ;
        RECT -21.780 -188.815 -20.340 -188.525 ;
        RECT -20.090 -188.625 -17.175 -188.505 ;
        RECT -20.090 -188.730 -19.135 -188.625 ;
        RECT -21.780 -188.840 -20.940 -188.815 ;
        RECT -22.160 -189.550 -21.990 -189.090 ;
        RECT -21.670 -189.805 -21.500 -189.010 ;
        RECT -20.640 -189.180 -20.340 -188.815 ;
        RECT -20.065 -189.305 -19.765 -188.730 ;
        RECT -19.515 -188.785 -19.135 -188.730 ;
        RECT -19.365 -189.090 -19.135 -188.785 ;
        RECT -19.335 -189.550 -19.165 -189.090 ;
        RECT -18.845 -189.805 -18.675 -189.010 ;
        RECT -18.385 -189.090 -18.155 -188.625 ;
        RECT -18.355 -189.550 -18.185 -189.090 ;
        RECT -17.865 -189.805 -17.695 -189.010 ;
        RECT -17.405 -189.090 -17.175 -188.625 ;
        RECT -16.995 -188.515 -16.155 -188.470 ;
        RECT -15.170 -188.515 -14.295 -188.075 ;
        RECT -11.750 -188.345 -11.515 -187.610 ;
        RECT -11.295 -188.315 -10.925 -187.475 ;
        RECT -10.620 -188.070 -10.450 -187.110 ;
        RECT -9.640 -188.070 -9.470 -187.110 ;
        RECT -8.660 -187.130 -8.490 -187.110 ;
        RECT -16.995 -188.800 -14.295 -188.515 ;
        RECT -12.375 -188.715 -11.515 -188.345 ;
        RECT -16.995 -188.840 -16.155 -188.800 ;
        RECT -15.170 -188.910 -14.295 -188.800 ;
        RECT -17.375 -189.550 -17.205 -189.090 ;
        RECT -16.885 -189.805 -16.715 -189.010 ;
        RECT -15.170 -189.080 -12.015 -188.910 ;
        RECT -15.170 -189.115 -14.960 -189.080 ;
        RECT -15.165 -189.280 -14.960 -189.115 ;
        RECT -15.165 -189.330 -14.930 -189.280 ;
        RECT -28.185 -190.200 -25.020 -190.030 ;
        RECT -24.125 -190.145 -16.670 -189.805 ;
        RECT -15.160 -189.940 -14.930 -189.330 ;
        RECT -14.655 -189.740 -14.485 -189.260 ;
        RECT -14.180 -189.325 -13.975 -189.080 ;
        RECT -14.685 -190.030 -14.465 -189.740 ;
        RECT -14.165 -189.800 -13.995 -189.325 ;
        RECT -13.675 -189.685 -13.505 -189.260 ;
        RECT -13.210 -189.325 -13.005 -189.080 ;
        RECT -13.700 -190.030 -13.480 -189.685 ;
        RECT -13.185 -189.800 -13.015 -189.325 ;
        RECT -12.695 -189.685 -12.525 -189.260 ;
        RECT -12.220 -189.285 -12.015 -189.080 ;
        RECT -12.720 -190.030 -12.500 -189.685 ;
        RECT -12.205 -189.800 -12.035 -189.285 ;
        RECT -11.750 -189.390 -11.515 -188.715 ;
        RECT -11.290 -188.435 -10.925 -188.315 ;
        RECT -10.650 -188.395 -10.420 -188.070 ;
        RECT -9.670 -188.395 -9.440 -188.070 ;
        RECT -8.690 -188.395 -8.460 -187.130 ;
        RECT -7.670 -188.040 -7.385 -187.220 ;
        RECT -6.210 -188.070 -6.040 -187.110 ;
        RECT -5.230 -188.070 -5.060 -187.110 ;
        RECT -4.250 -187.130 -4.080 -187.110 ;
        RECT -10.650 -188.435 -8.460 -188.395 ;
        RECT -6.240 -188.395 -6.010 -188.070 ;
        RECT -5.260 -188.395 -5.030 -188.070 ;
        RECT -4.280 -188.395 -4.050 -187.130 ;
        RECT -6.240 -188.435 -4.050 -188.395 ;
        RECT -11.290 -188.625 -8.460 -188.435 ;
        RECT -11.290 -188.785 -10.420 -188.625 ;
        RECT -10.650 -189.090 -10.420 -188.785 ;
        RECT -11.715 -189.740 -11.545 -189.390 ;
        RECT -10.620 -189.550 -10.450 -189.090 ;
        RECT -11.740 -190.030 -11.520 -189.740 ;
        RECT -10.130 -189.805 -9.960 -189.010 ;
        RECT -9.670 -189.090 -9.440 -188.625 ;
        RECT -9.640 -189.550 -9.470 -189.090 ;
        RECT -9.150 -189.805 -8.980 -189.010 ;
        RECT -8.690 -189.090 -8.460 -188.625 ;
        RECT -6.980 -188.545 -6.680 -188.525 ;
        RECT -6.390 -188.545 -4.050 -188.435 ;
        RECT -6.980 -188.625 -4.050 -188.545 ;
        RECT -6.980 -188.755 -6.010 -188.625 ;
        RECT -8.660 -189.550 -8.490 -189.090 ;
        RECT -8.170 -189.805 -8.000 -189.010 ;
        RECT -6.980 -189.185 -6.680 -188.755 ;
        RECT -6.390 -188.785 -6.010 -188.755 ;
        RECT -6.240 -189.090 -6.010 -188.785 ;
        RECT -6.210 -189.550 -6.040 -189.090 ;
        RECT -5.720 -189.805 -5.550 -189.010 ;
        RECT -5.260 -189.090 -5.030 -188.625 ;
        RECT -5.230 -189.550 -5.060 -189.090 ;
        RECT -4.740 -189.805 -4.570 -189.010 ;
        RECT -4.280 -189.090 -4.050 -188.625 ;
        RECT -4.250 -189.550 -4.080 -189.090 ;
        RECT -3.760 -189.805 -3.590 -189.010 ;
        RECT -1.560 -189.245 -1.390 -187.195 ;
        RECT 2.130 -188.415 2.300 -187.195 ;
        RECT 3.110 -188.415 3.280 -187.195 ;
        RECT 4.090 -188.415 4.260 -187.195 ;
        RECT 1.485 -188.600 4.260 -188.415 ;
        RECT 5.190 -188.430 5.420 -188.010 ;
        RECT 7.105 -188.120 7.275 -187.260 ;
        RECT 8.085 -187.800 8.255 -187.260 ;
        RECT 9.065 -187.800 9.235 -187.260 ;
        RECT -2.315 -189.510 -1.390 -189.245 ;
        RECT -1.215 -189.290 -0.540 -189.240 ;
        RECT 1.485 -189.290 1.670 -188.600 ;
        RECT 4.460 -188.700 5.420 -188.430 ;
        RECT 6.420 -188.470 7.275 -188.120 ;
        RECT 9.460 -188.035 9.825 -187.970 ;
        RECT 9.460 -188.175 10.325 -188.035 ;
        RECT 9.460 -188.240 10.435 -188.175 ;
        RECT 9.460 -188.270 9.825 -188.240 ;
        RECT 2.780 -188.885 3.455 -188.840 ;
        RECT 5.595 -188.885 6.275 -188.880 ;
        RECT 2.780 -189.075 6.275 -188.885 ;
        RECT 2.780 -189.110 3.455 -189.075 ;
        RECT 5.595 -189.110 6.275 -189.075 ;
        RECT -1.215 -189.475 1.670 -189.290 ;
        RECT -1.215 -189.510 -0.540 -189.475 ;
        RECT -14.685 -190.200 -11.520 -190.030 ;
        RECT -10.625 -190.145 -3.545 -189.805 ;
        RECT -35.210 -190.910 -34.290 -190.595 ;
        RECT -35.105 -190.915 -34.290 -190.910 ;
        RECT -33.435 -191.150 -33.135 -190.465 ;
        RECT -20.885 -190.810 -20.200 -190.760 ;
        RECT -16.155 -190.810 -15.495 -190.755 ;
        RECT -6.085 -190.810 -5.425 -190.760 ;
        RECT -31.780 -191.005 -5.425 -190.810 ;
        RECT -20.885 -191.060 -20.200 -191.005 ;
        RECT -16.155 -191.055 -15.495 -191.005 ;
        RECT -6.085 -191.060 -5.425 -191.005 ;
        RECT -33.430 -193.010 -33.190 -191.150 ;
        RECT -31.695 -191.270 -31.010 -191.205 ;
        RECT -18.710 -191.270 -18.025 -191.175 ;
        RECT -4.870 -191.270 -4.210 -191.175 ;
        RECT -31.780 -191.465 -4.205 -191.270 ;
        RECT -31.695 -191.505 -31.010 -191.465 ;
        RECT -31.640 -191.705 -31.085 -191.505 ;
        RECT -27.585 -191.705 -27.030 -191.465 ;
        RECT -18.710 -191.475 -18.025 -191.465 ;
        RECT -32.880 -192.045 -26.025 -191.705 ;
        RECT -25.130 -191.820 -21.965 -191.650 ;
        RECT -18.595 -191.705 -18.040 -191.475 ;
        RECT -17.680 -191.705 -15.080 -191.695 ;
        RECT -14.205 -191.705 -13.650 -191.465 ;
        RECT -32.835 -192.840 -32.665 -192.045 ;
        RECT -32.345 -192.760 -32.175 -192.300 ;
        RECT -33.430 -193.230 -32.555 -193.010 ;
        RECT -33.395 -193.380 -32.555 -193.230 ;
        RECT -32.375 -193.225 -32.145 -192.760 ;
        RECT -31.855 -192.840 -31.685 -192.045 ;
        RECT -31.365 -192.760 -31.195 -192.300 ;
        RECT -31.395 -193.225 -31.165 -192.760 ;
        RECT -30.875 -192.840 -30.705 -192.045 ;
        RECT -30.385 -192.760 -30.215 -192.300 ;
        RECT -30.415 -193.065 -30.185 -192.760 ;
        RECT -28.650 -192.840 -28.480 -192.045 ;
        RECT -28.160 -192.760 -27.990 -192.300 ;
        RECT -30.415 -193.225 -29.750 -193.065 ;
        RECT -62.510 -195.440 -61.835 -195.410 ;
        RECT -62.610 -195.450 -61.835 -195.440 ;
        RECT -93.935 -196.650 -76.245 -195.620 ;
        RECT -63.645 -195.630 -61.835 -195.450 ;
        RECT -61.595 -195.525 -59.445 -195.375 ;
        RECT -61.595 -195.565 -59.500 -195.525 ;
        RECT -58.550 -195.585 -58.380 -194.805 ;
        RECT -58.060 -195.345 -57.890 -194.805 ;
        RECT -57.570 -195.585 -57.400 -194.805 ;
        RECT -57.080 -195.345 -56.910 -194.805 ;
        RECT -56.590 -194.860 -54.730 -194.510 ;
        RECT -32.375 -193.415 -29.750 -193.225 ;
        RECT -32.375 -193.455 -30.185 -193.415 ;
        RECT -32.375 -194.720 -32.145 -193.455 ;
        RECT -31.395 -193.780 -31.165 -193.455 ;
        RECT -30.415 -193.780 -30.185 -193.455 ;
        RECT -32.345 -194.740 -32.175 -194.720 ;
        RECT -31.365 -194.740 -31.195 -193.780 ;
        RECT -30.385 -194.740 -30.215 -193.780 ;
        RECT -29.980 -194.065 -29.750 -193.415 ;
        RECT -28.190 -193.225 -27.960 -192.760 ;
        RECT -27.670 -192.840 -27.500 -192.045 ;
        RECT -27.180 -192.760 -27.010 -192.300 ;
        RECT -27.210 -193.225 -26.980 -192.760 ;
        RECT -26.690 -192.840 -26.520 -192.045 ;
        RECT -25.130 -192.110 -24.910 -191.820 ;
        RECT -26.200 -192.760 -26.030 -192.300 ;
        RECT -25.105 -192.460 -24.935 -192.110 ;
        RECT -26.230 -193.065 -26.000 -192.760 ;
        RECT -26.230 -193.225 -25.360 -193.065 ;
        RECT -28.190 -193.415 -25.360 -193.225 ;
        RECT -28.190 -193.455 -26.000 -193.415 ;
        RECT -29.265 -194.065 -28.980 -193.810 ;
        RECT -29.980 -194.310 -28.980 -194.065 ;
        RECT -29.265 -194.630 -28.980 -194.310 ;
        RECT -28.190 -194.720 -27.960 -193.455 ;
        RECT -27.210 -193.780 -26.980 -193.455 ;
        RECT -26.230 -193.780 -26.000 -193.455 ;
        RECT -25.725 -193.535 -25.360 -193.415 ;
        RECT -25.135 -193.135 -24.900 -192.460 ;
        RECT -24.615 -192.565 -24.445 -192.050 ;
        RECT -24.150 -192.165 -23.930 -191.820 ;
        RECT -24.635 -192.770 -24.430 -192.565 ;
        RECT -24.125 -192.590 -23.955 -192.165 ;
        RECT -23.635 -192.525 -23.465 -192.050 ;
        RECT -23.170 -192.165 -22.950 -191.820 ;
        RECT -23.645 -192.770 -23.440 -192.525 ;
        RECT -23.145 -192.590 -22.975 -192.165 ;
        RECT -22.655 -192.525 -22.485 -192.050 ;
        RECT -22.185 -192.110 -21.965 -191.820 ;
        RECT -19.380 -192.035 -12.525 -191.705 ;
        RECT -19.380 -192.045 -16.710 -192.035 ;
        RECT -15.195 -192.045 -12.525 -192.035 ;
        RECT -11.630 -191.820 -8.465 -191.650 ;
        RECT -22.675 -192.770 -22.470 -192.525 ;
        RECT -22.165 -192.590 -21.995 -192.110 ;
        RECT -21.675 -192.520 -21.505 -192.050 ;
        RECT -21.690 -192.735 -21.485 -192.520 ;
        RECT -21.690 -192.770 -21.480 -192.735 ;
        RECT -24.635 -192.940 -21.480 -192.770 ;
        RECT -19.335 -192.840 -19.165 -192.045 ;
        RECT -18.845 -192.760 -18.675 -192.300 ;
        RECT -25.135 -193.505 -24.275 -193.135 ;
        RECT -22.355 -193.240 -21.025 -192.940 ;
        RECT -19.895 -193.045 -19.055 -193.010 ;
        RECT -28.160 -194.740 -27.990 -194.720 ;
        RECT -27.180 -194.740 -27.010 -193.780 ;
        RECT -26.200 -194.740 -26.030 -193.780 ;
        RECT -25.725 -194.375 -25.355 -193.535 ;
        RECT -25.135 -194.240 -24.900 -193.505 ;
        RECT -22.355 -193.775 -21.480 -193.240 ;
        RECT -20.005 -193.345 -19.055 -193.045 ;
        RECT -19.895 -193.380 -19.055 -193.345 ;
        RECT -18.875 -193.225 -18.645 -192.760 ;
        RECT -18.355 -192.840 -18.185 -192.045 ;
        RECT -17.865 -192.760 -17.695 -192.300 ;
        RECT -17.895 -193.225 -17.665 -192.760 ;
        RECT -17.375 -192.840 -17.205 -192.045 ;
        RECT -16.885 -192.760 -16.715 -192.300 ;
        RECT -16.915 -193.065 -16.685 -192.760 ;
        RECT -16.010 -193.010 -15.710 -192.215 ;
        RECT -15.150 -192.840 -14.980 -192.045 ;
        RECT -14.660 -192.760 -14.490 -192.300 ;
        RECT -16.915 -193.225 -16.195 -193.065 ;
        RECT -24.620 -193.945 -21.480 -193.775 ;
        RECT -24.620 -194.205 -24.440 -193.945 ;
        RECT -23.630 -194.125 -23.450 -193.945 ;
        RECT -25.105 -194.610 -24.935 -194.240 ;
        RECT -25.110 -194.835 -24.930 -194.610 ;
        RECT -24.615 -194.665 -24.445 -194.205 ;
        RECT -24.125 -194.560 -23.955 -194.125 ;
        RECT -23.635 -194.215 -23.450 -194.125 ;
        RECT -24.130 -194.835 -23.920 -194.560 ;
        RECT -23.635 -194.665 -23.465 -194.215 ;
        RECT -23.145 -194.555 -22.975 -194.125 ;
        RECT -22.660 -194.215 -22.480 -193.945 ;
        RECT -23.160 -194.835 -22.950 -194.555 ;
        RECT -22.655 -194.665 -22.485 -194.215 ;
        RECT -22.165 -194.580 -21.995 -194.125 ;
        RECT -21.690 -194.165 -21.480 -193.945 ;
        RECT -18.875 -193.415 -16.195 -193.225 ;
        RECT -16.010 -193.325 -14.870 -193.010 ;
        RECT -15.710 -193.380 -14.870 -193.325 ;
        RECT -14.690 -193.225 -14.460 -192.760 ;
        RECT -14.170 -192.840 -14.000 -192.045 ;
        RECT -13.680 -192.760 -13.510 -192.300 ;
        RECT -13.710 -193.225 -13.480 -192.760 ;
        RECT -13.190 -192.840 -13.020 -192.045 ;
        RECT -11.630 -192.110 -11.410 -191.820 ;
        RECT -12.700 -192.760 -12.530 -192.300 ;
        RECT -11.605 -192.460 -11.435 -192.110 ;
        RECT -12.730 -193.065 -12.500 -192.760 ;
        RECT -12.730 -193.225 -11.860 -193.065 ;
        RECT -18.875 -193.455 -16.685 -193.415 ;
        RECT -22.180 -194.835 -21.970 -194.580 ;
        RECT -21.675 -194.665 -21.505 -194.165 ;
        RECT -18.875 -194.720 -18.645 -193.455 ;
        RECT -17.895 -193.780 -17.665 -193.455 ;
        RECT -16.915 -193.780 -16.685 -193.455 ;
        RECT -18.845 -194.740 -18.675 -194.720 ;
        RECT -17.865 -194.740 -17.695 -193.780 ;
        RECT -16.885 -194.740 -16.715 -193.780 ;
        RECT -16.505 -194.060 -16.195 -193.415 ;
        RECT -14.690 -193.415 -11.860 -193.225 ;
        RECT -14.690 -193.455 -12.500 -193.415 ;
        RECT -15.765 -194.060 -15.480 -193.810 ;
        RECT -16.505 -194.370 -15.480 -194.060 ;
        RECT -15.765 -194.630 -15.480 -194.370 ;
        RECT -14.690 -194.720 -14.460 -193.455 ;
        RECT -13.710 -193.780 -13.480 -193.455 ;
        RECT -12.730 -193.780 -12.500 -193.455 ;
        RECT -12.225 -193.535 -11.860 -193.415 ;
        RECT -11.635 -193.135 -11.400 -192.460 ;
        RECT -11.115 -192.565 -10.945 -192.050 ;
        RECT -10.650 -192.165 -10.430 -191.820 ;
        RECT -11.135 -192.770 -10.930 -192.565 ;
        RECT -10.625 -192.590 -10.455 -192.165 ;
        RECT -10.135 -192.525 -9.965 -192.050 ;
        RECT -9.670 -192.165 -9.450 -191.820 ;
        RECT -10.145 -192.770 -9.940 -192.525 ;
        RECT -9.645 -192.590 -9.475 -192.165 ;
        RECT -9.155 -192.525 -8.985 -192.050 ;
        RECT -8.685 -192.110 -8.465 -191.820 ;
        RECT -9.175 -192.770 -8.970 -192.525 ;
        RECT -8.665 -192.590 -8.495 -192.110 ;
        RECT -8.175 -192.520 -8.005 -192.050 ;
        RECT -8.190 -192.735 -7.985 -192.520 ;
        RECT -8.190 -192.770 -7.980 -192.735 ;
        RECT -11.135 -192.930 -7.980 -192.770 ;
        RECT -11.135 -192.940 -7.605 -192.930 ;
        RECT -11.635 -193.505 -10.775 -193.135 ;
        RECT -8.855 -193.230 -7.605 -192.940 ;
        RECT -14.660 -194.740 -14.490 -194.720 ;
        RECT -13.680 -194.740 -13.510 -193.780 ;
        RECT -12.700 -194.740 -12.530 -193.780 ;
        RECT -12.225 -194.375 -11.855 -193.535 ;
        RECT -11.635 -194.240 -11.400 -193.505 ;
        RECT -8.855 -193.775 -7.980 -193.230 ;
        RECT -11.120 -193.945 -7.980 -193.775 ;
        RECT -11.120 -194.205 -10.940 -193.945 ;
        RECT -10.130 -194.125 -9.950 -193.945 ;
        RECT -11.605 -194.610 -11.435 -194.240 ;
        RECT -25.110 -195.005 -21.970 -194.835 ;
        RECT -11.610 -194.835 -11.430 -194.610 ;
        RECT -11.115 -194.665 -10.945 -194.205 ;
        RECT -10.625 -194.560 -10.455 -194.125 ;
        RECT -10.135 -194.215 -9.950 -194.125 ;
        RECT -10.630 -194.835 -10.420 -194.560 ;
        RECT -10.135 -194.665 -9.965 -194.215 ;
        RECT -9.645 -194.555 -9.475 -194.125 ;
        RECT -9.160 -194.215 -8.980 -193.945 ;
        RECT -9.660 -194.835 -9.450 -194.555 ;
        RECT -9.155 -194.665 -8.985 -194.215 ;
        RECT -8.665 -194.580 -8.495 -194.125 ;
        RECT -8.190 -194.165 -7.980 -193.945 ;
        RECT -8.680 -194.835 -8.470 -194.580 ;
        RECT -8.175 -194.665 -8.005 -194.165 ;
        RECT -6.785 -194.365 -5.295 -191.465 ;
        RECT -4.870 -191.475 -4.210 -191.465 ;
        RECT -1.560 -191.775 -1.390 -189.510 ;
        RECT 1.485 -189.745 1.670 -189.475 ;
        RECT 1.840 -189.295 2.515 -189.230 ;
        RECT 6.450 -189.295 6.620 -188.470 ;
        RECT 7.595 -188.955 7.765 -188.415 ;
        RECT 8.085 -189.195 8.255 -188.415 ;
        RECT 8.575 -188.955 8.745 -188.415 ;
        RECT 9.065 -189.195 9.235 -188.415 ;
        RECT 10.130 -188.985 10.435 -188.240 ;
        RECT 11.130 -188.985 11.300 -187.265 ;
        RECT 12.110 -188.985 12.280 -187.265 ;
        RECT 10.130 -189.135 12.280 -188.985 ;
        RECT 13.230 -189.020 13.410 -185.270 ;
        RECT 10.185 -189.175 12.280 -189.135 ;
        RECT 12.520 -189.060 13.410 -189.020 ;
        RECT 1.840 -189.465 6.620 -189.295 ;
        RECT 1.840 -189.500 2.515 -189.465 ;
        RECT 6.860 -189.625 9.935 -189.195 ;
        RECT 12.520 -189.240 13.455 -189.060 ;
        RECT 12.520 -189.260 13.345 -189.240 ;
        RECT 12.520 -189.290 13.195 -189.260 ;
        RECT 10.500 -189.540 10.870 -189.410 ;
        RECT 13.635 -189.530 13.835 -184.850 ;
        RECT 15.130 -188.130 15.300 -187.270 ;
        RECT 16.110 -187.810 16.280 -187.270 ;
        RECT 17.090 -187.810 17.260 -187.270 ;
        RECT 12.925 -189.540 13.835 -189.530 ;
        RECT 0.505 -189.915 1.670 -189.745 ;
        RECT 2.535 -189.915 4.750 -189.745 ;
        RECT -1.070 -192.715 -0.900 -190.735 ;
        RECT 0.505 -191.775 0.675 -189.915 ;
        RECT 0.995 -192.265 1.165 -190.235 ;
        RECT 1.485 -191.775 1.655 -189.915 ;
        RECT 2.535 -189.920 3.770 -189.915 ;
        RECT 2.535 -190.235 2.710 -189.920 ;
        RECT 2.050 -191.720 2.220 -190.235 ;
        RECT 2.045 -192.250 2.220 -191.720 ;
        RECT 2.540 -191.775 2.710 -190.235 ;
        RECT 3.030 -191.730 3.200 -190.235 ;
        RECT 3.025 -192.250 3.200 -191.730 ;
        RECT 3.600 -191.770 3.770 -189.920 ;
        RECT 2.045 -192.265 3.200 -192.250 ;
        RECT 0.995 -192.435 3.200 -192.265 ;
        RECT 4.090 -192.715 4.260 -190.230 ;
        RECT 4.580 -191.770 4.750 -189.915 ;
        RECT 8.410 -191.660 8.715 -189.625 ;
        RECT 10.500 -189.730 13.835 -189.540 ;
        RECT 14.310 -188.480 15.300 -188.130 ;
        RECT 17.485 -188.045 17.850 -187.980 ;
        RECT 17.485 -188.185 18.350 -188.045 ;
        RECT 17.485 -188.250 18.460 -188.185 ;
        RECT 17.485 -188.280 17.850 -188.250 ;
        RECT 10.500 -189.735 12.930 -189.730 ;
        RECT 10.500 -189.765 10.870 -189.735 ;
        RECT 12.575 -189.740 12.930 -189.735 ;
        RECT 10.640 -191.490 10.810 -189.950 ;
        RECT 11.130 -191.490 11.300 -189.950 ;
        RECT 11.620 -191.490 11.790 -189.950 ;
        RECT 12.110 -191.490 12.280 -189.950 ;
        RECT 12.600 -191.490 12.770 -189.950 ;
        RECT 8.410 -191.750 10.660 -191.660 ;
        RECT 12.110 -191.750 12.285 -191.490 ;
        RECT 8.410 -191.965 12.870 -191.750 ;
        RECT -1.620 -193.040 4.750 -192.715 ;
        RECT -1.555 -194.365 -0.905 -193.040 ;
        RECT -0.025 -194.365 0.625 -193.040 ;
        RECT 1.560 -194.365 2.210 -193.040 ;
        RECT 3.790 -194.365 4.440 -193.040 ;
        RECT 8.410 -194.365 9.165 -191.965 ;
        RECT 10.295 -192.055 12.870 -191.965 ;
        RECT 10.295 -194.365 10.915 -192.055 ;
        RECT 11.945 -194.365 12.565 -192.055 ;
        RECT 14.310 -192.155 14.660 -188.480 ;
        RECT 15.620 -188.965 15.790 -188.425 ;
        RECT 16.110 -189.205 16.280 -188.425 ;
        RECT 16.600 -188.965 16.770 -188.425 ;
        RECT 17.090 -189.205 17.260 -188.425 ;
        RECT 18.155 -188.995 18.460 -188.250 ;
        RECT 19.155 -188.995 19.325 -187.275 ;
        RECT 20.135 -188.995 20.305 -187.275 ;
        RECT 18.155 -189.145 20.305 -188.995 ;
        RECT 18.210 -189.185 20.305 -189.145 ;
        RECT 20.545 -189.060 21.220 -189.030 ;
        RECT 21.400 -189.060 21.580 -182.425 ;
        RECT 14.885 -189.635 17.960 -189.205 ;
        RECT 20.545 -189.250 21.580 -189.060 ;
        RECT 20.545 -189.260 21.480 -189.250 ;
        RECT 20.545 -189.300 21.220 -189.260 ;
        RECT 18.525 -189.550 18.895 -189.420 ;
        RECT 21.775 -189.540 21.975 -182.075 ;
        RECT 20.950 -189.550 21.975 -189.540 ;
        RECT 13.980 -192.385 14.660 -192.155 ;
        RECT 16.435 -191.670 16.740 -189.635 ;
        RECT 18.525 -189.740 21.975 -189.550 ;
        RECT 18.525 -189.745 20.955 -189.740 ;
        RECT 18.525 -189.775 18.895 -189.745 ;
        RECT 20.600 -189.750 20.955 -189.745 ;
        RECT 18.665 -191.500 18.835 -189.960 ;
        RECT 19.155 -191.500 19.325 -189.960 ;
        RECT 19.645 -191.500 19.815 -189.960 ;
        RECT 20.135 -191.500 20.305 -189.960 ;
        RECT 20.625 -191.500 20.795 -189.960 ;
        RECT 23.250 -190.150 23.420 -187.150 ;
        RECT 26.940 -188.370 27.110 -187.150 ;
        RECT 27.920 -188.370 28.090 -187.150 ;
        RECT 28.900 -188.370 29.070 -187.150 ;
        RECT 26.295 -188.555 29.070 -188.370 ;
        RECT 29.270 -188.425 29.945 -188.385 ;
        RECT 23.595 -189.245 24.270 -189.195 ;
        RECT 26.295 -189.245 26.480 -188.555 ;
        RECT 29.265 -188.610 30.040 -188.425 ;
        RECT 29.265 -188.655 29.945 -188.610 ;
        RECT 27.590 -188.840 28.265 -188.795 ;
        RECT 30.225 -188.840 30.395 -181.995 ;
        RECT 27.590 -189.030 30.395 -188.840 ;
        RECT 27.590 -189.065 28.265 -189.030 ;
        RECT 23.595 -189.430 26.480 -189.245 ;
        RECT 23.595 -189.465 24.270 -189.430 ;
        RECT 26.295 -189.700 26.480 -189.430 ;
        RECT 26.650 -189.250 27.325 -189.185 ;
        RECT 30.575 -189.250 30.745 -181.535 ;
        RECT 31.315 -186.685 34.955 -186.515 ;
        RECT 31.315 -188.245 31.485 -186.685 ;
        RECT 31.805 -188.425 31.975 -187.205 ;
        RECT 32.295 -188.245 32.465 -186.685 ;
        RECT 32.895 -187.030 34.605 -186.860 ;
        RECT 32.895 -188.245 33.065 -187.030 ;
        RECT 33.385 -188.425 33.555 -187.205 ;
        RECT 33.875 -188.245 34.045 -187.030 ;
        RECT 31.060 -188.595 34.130 -188.425 ;
        RECT 26.650 -189.420 30.745 -189.250 ;
        RECT 31.310 -189.265 32.005 -188.995 ;
        RECT 33.960 -189.170 34.130 -188.595 ;
        RECT 34.435 -188.790 34.605 -187.030 ;
        RECT 34.785 -188.420 34.955 -186.685 ;
        RECT 35.685 -188.420 35.855 -187.205 ;
        RECT 34.785 -188.590 35.855 -188.420 ;
        RECT 36.665 -188.790 36.835 -187.205 ;
        RECT 38.215 -188.170 38.385 -187.205 ;
        RECT 39.760 -188.160 39.930 -187.205 ;
        RECT 34.435 -188.960 36.835 -188.790 ;
        RECT 37.100 -189.045 37.795 -188.775 ;
        RECT 33.960 -189.340 34.690 -189.170 ;
        RECT 26.650 -189.455 27.325 -189.420 ;
        RECT 34.520 -189.650 34.690 -189.340 ;
        RECT 35.055 -189.415 35.750 -189.145 ;
        RECT 22.170 -190.440 23.420 -190.150 ;
        RECT 16.435 -191.760 18.685 -191.670 ;
        RECT 20.135 -191.760 20.310 -191.500 ;
        RECT 16.435 -191.975 20.895 -191.760 ;
        RECT 16.435 -194.365 17.190 -191.975 ;
        RECT 18.645 -192.065 20.895 -191.975 ;
        RECT 18.645 -194.365 19.400 -192.065 ;
        RECT 20.110 -194.365 20.865 -192.065 ;
        RECT 22.170 -192.715 22.495 -190.440 ;
        RECT 23.250 -191.730 23.420 -190.440 ;
        RECT 25.315 -189.870 26.480 -189.700 ;
        RECT 27.345 -189.870 29.560 -189.700 ;
        RECT 23.740 -192.670 23.910 -190.690 ;
        RECT 25.315 -191.730 25.485 -189.870 ;
        RECT 25.805 -192.220 25.975 -190.190 ;
        RECT 26.295 -191.730 26.465 -189.870 ;
        RECT 27.345 -189.875 28.580 -189.870 ;
        RECT 27.345 -190.190 27.520 -189.875 ;
        RECT 26.860 -191.675 27.030 -190.190 ;
        RECT 26.855 -192.205 27.030 -191.675 ;
        RECT 27.350 -191.730 27.520 -190.190 ;
        RECT 27.840 -191.685 28.010 -190.190 ;
        RECT 27.835 -192.205 28.010 -191.685 ;
        RECT 28.410 -191.725 28.580 -189.875 ;
        RECT 26.855 -192.220 28.010 -192.205 ;
        RECT 25.805 -192.390 28.010 -192.220 ;
        RECT 28.900 -192.670 29.070 -190.185 ;
        RECT 29.390 -191.725 29.560 -189.870 ;
        RECT 31.305 -189.855 32.960 -189.670 ;
        RECT 34.520 -189.820 37.325 -189.650 ;
        RECT 31.305 -190.270 31.490 -189.855 ;
        RECT 32.775 -189.975 32.960 -189.855 ;
        RECT 32.775 -190.160 33.555 -189.975 ;
        RECT 31.315 -191.215 31.485 -190.270 ;
        RECT 31.295 -191.830 31.490 -191.215 ;
        RECT 31.805 -191.460 31.975 -190.235 ;
        RECT 33.370 -190.265 33.555 -190.160 ;
        RECT 33.385 -191.275 33.555 -190.265 ;
        RECT 33.865 -190.280 35.365 -190.085 ;
        RECT 33.875 -191.275 34.045 -190.280 ;
        RECT 35.195 -191.275 35.365 -190.280 ;
        RECT 35.685 -191.275 35.855 -189.820 ;
        RECT 36.665 -191.190 36.835 -190.235 ;
        RECT 36.665 -191.460 36.845 -191.190 ;
        RECT 37.155 -191.275 37.325 -189.820 ;
        RECT 38.190 -189.865 38.405 -188.170 ;
        RECT 39.740 -189.145 39.955 -188.160 ;
        RECT 40.175 -189.075 40.870 -188.805 ;
        RECT 39.240 -189.375 39.955 -189.145 ;
        RECT 37.710 -190.095 38.405 -189.865 ;
        RECT 38.190 -190.320 38.405 -190.095 ;
        RECT 38.215 -191.275 38.385 -190.320 ;
        RECT 38.705 -191.240 38.875 -190.235 ;
        RECT 39.740 -190.330 39.955 -189.375 ;
        RECT 31.805 -191.640 36.845 -191.460 ;
        RECT 38.680 -191.660 38.895 -191.240 ;
        RECT 39.760 -191.275 39.930 -190.330 ;
        RECT 40.250 -191.230 40.420 -190.235 ;
        RECT 40.225 -191.660 40.440 -191.230 ;
        RECT 37.300 -191.830 40.460 -191.660 ;
        RECT 31.295 -192.095 40.460 -191.830 ;
        RECT 21.820 -192.945 22.500 -192.715 ;
        RECT 23.190 -192.995 29.560 -192.670 ;
        RECT 23.310 -194.365 24.040 -192.995 ;
        RECT 25.535 -194.365 26.265 -192.995 ;
        RECT 26.865 -194.365 27.595 -192.995 ;
        RECT 28.665 -194.365 29.395 -192.995 ;
        RECT 31.485 -194.365 32.470 -192.095 ;
        RECT 34.150 -194.365 35.135 -192.095 ;
        RECT 36.715 -192.140 40.460 -192.095 ;
        RECT 36.715 -194.365 37.700 -192.140 ;
        RECT 39.230 -194.365 40.215 -192.140 ;
        RECT 41.205 -194.365 42.510 -180.950 ;
        RECT 44.690 -181.205 81.020 -180.510 ;
        RECT 79.395 -185.605 80.730 -185.425 ;
        RECT 52.670 -186.780 80.730 -185.605 ;
        RECT 79.395 -186.915 80.730 -186.780 ;
        RECT 44.830 -188.575 45.920 -188.535 ;
        RECT 80.710 -188.575 81.475 -188.380 ;
        RECT 44.830 -188.950 81.475 -188.575 ;
        RECT 44.830 -188.980 45.920 -188.950 ;
        RECT 80.710 -189.135 81.475 -188.950 ;
        RECT 49.740 -189.680 49.990 -189.650 ;
        RECT 77.300 -189.680 77.790 -189.610 ;
        RECT 49.695 -190.295 77.790 -189.680 ;
        RECT 49.740 -190.315 49.990 -190.295 ;
        RECT 77.300 -190.430 77.790 -190.295 ;
        RECT 81.885 -191.705 82.525 -177.145 ;
        RECT 83.150 -191.260 83.810 -175.005 ;
        RECT 84.360 -188.380 84.805 -172.630 ;
        RECT 94.820 -178.700 97.545 -171.010 ;
        RECT 91.905 -181.230 421.770 -178.700 ;
        RECT 84.360 -189.135 84.845 -188.380 ;
        RECT 94.820 -188.550 97.545 -181.230 ;
        RECT 143.550 -183.535 144.965 -181.230 ;
        RECT 142.330 -183.675 145.655 -183.535 ;
        RECT 170.390 -183.610 172.175 -183.275 ;
        RECT 176.280 -183.610 178.065 -183.445 ;
        RECT 185.545 -183.590 186.960 -181.230 ;
        RECT 142.330 -183.965 147.505 -183.675 ;
        RECT 142.330 -184.370 142.760 -183.965 ;
        RECT 143.630 -184.150 143.805 -183.965 ;
        RECT 145.255 -183.980 147.505 -183.965 ;
        RECT 138.070 -184.800 142.760 -184.370 ;
        RECT 137.310 -186.250 137.960 -185.790 ;
        RECT 138.770 -186.080 138.940 -184.800 ;
        RECT 139.260 -186.080 139.430 -185.040 ;
        RECT 139.750 -186.080 139.920 -184.800 ;
        RECT 140.240 -185.910 140.410 -185.040 ;
        RECT 143.145 -185.690 143.315 -184.150 ;
        RECT 143.635 -185.690 143.805 -184.150 ;
        RECT 144.125 -185.690 144.295 -184.150 ;
        RECT 144.615 -185.690 144.785 -184.150 ;
        RECT 145.105 -185.690 145.275 -184.150 ;
        RECT 142.985 -185.905 143.340 -185.900 ;
        RECT 145.045 -185.905 145.415 -185.875 ;
        RECT 142.985 -185.910 145.415 -185.905 ;
        RECT 140.240 -186.080 145.415 -185.910 ;
        RECT 147.200 -186.015 147.505 -183.980 ;
        RECT 170.390 -184.555 178.065 -183.610 ;
        RECT 184.530 -183.730 187.855 -183.590 ;
        RECT 184.530 -184.020 189.705 -183.730 ;
        RECT 230.105 -183.785 231.520 -181.230 ;
        RECT 276.200 -183.615 277.615 -181.230 ;
        RECT 302.945 -183.455 304.825 -182.980 ;
        RECT 320.175 -183.285 321.710 -181.230 ;
        RECT 310.950 -183.455 312.200 -183.320 ;
        RECT 184.530 -184.425 184.960 -184.020 ;
        RECT 185.830 -184.205 186.005 -184.020 ;
        RECT 187.455 -184.035 189.705 -184.020 ;
        RECT 170.390 -184.610 172.175 -184.555 ;
        RECT 176.280 -184.780 178.065 -184.555 ;
        RECT 180.270 -184.855 184.960 -184.425 ;
        RECT 140.245 -186.100 145.415 -186.080 ;
        RECT 140.245 -186.110 142.990 -186.100 ;
        RECT 138.180 -186.250 138.545 -186.220 ;
        RECT 145.045 -186.230 145.415 -186.100 ;
        RECT 137.310 -186.455 138.545 -186.250 ;
        RECT 145.980 -186.445 149.905 -186.015 ;
        RECT 179.510 -186.305 180.160 -185.845 ;
        RECT 180.970 -186.135 181.140 -184.855 ;
        RECT 181.460 -186.135 181.630 -185.095 ;
        RECT 181.950 -186.135 182.120 -184.855 ;
        RECT 182.440 -185.965 182.610 -185.095 ;
        RECT 185.345 -185.745 185.515 -184.205 ;
        RECT 185.835 -185.745 186.005 -184.205 ;
        RECT 186.325 -185.745 186.495 -184.205 ;
        RECT 186.815 -185.745 186.985 -184.205 ;
        RECT 187.305 -185.745 187.475 -184.205 ;
        RECT 185.185 -185.960 185.540 -185.955 ;
        RECT 187.245 -185.960 187.615 -185.930 ;
        RECT 185.185 -185.965 187.615 -185.960 ;
        RECT 182.440 -186.135 187.615 -185.965 ;
        RECT 189.400 -186.070 189.705 -184.035 ;
        RECT 213.170 -184.055 214.495 -183.900 ;
        RECT 220.800 -184.055 222.285 -183.890 ;
        RECT 213.170 -184.890 222.285 -184.055 ;
        RECT 228.845 -183.925 232.170 -183.785 ;
        RECT 228.845 -184.215 234.020 -183.925 ;
        RECT 228.845 -184.620 229.275 -184.215 ;
        RECT 230.145 -184.400 230.320 -184.215 ;
        RECT 231.770 -184.230 234.020 -184.215 ;
        RECT 213.170 -185.225 214.495 -184.890 ;
        RECT 220.800 -185.000 222.285 -184.890 ;
        RECT 224.585 -185.050 229.275 -184.620 ;
        RECT 182.445 -186.155 187.615 -186.135 ;
        RECT 182.445 -186.165 185.190 -186.155 ;
        RECT 180.380 -186.305 180.745 -186.275 ;
        RECT 187.245 -186.285 187.615 -186.155 ;
        RECT 137.310 -186.540 137.960 -186.455 ;
        RECT 138.180 -186.520 138.545 -186.455 ;
        RECT 143.635 -186.505 145.730 -186.465 ;
        RECT 143.635 -186.655 145.785 -186.505 ;
        RECT 138.770 -187.730 138.940 -186.690 ;
        RECT 139.750 -187.730 139.920 -186.690 ;
        RECT 140.730 -187.730 140.900 -186.690 ;
        RECT 101.870 -188.360 105.010 -188.190 ;
        RECT 90.330 -189.080 99.180 -188.550 ;
        RECT 101.405 -189.030 101.575 -188.530 ;
        RECT 101.870 -188.615 102.080 -188.360 ;
        RECT 84.360 -190.800 84.805 -189.135 ;
        RECT 90.850 -189.810 91.090 -189.080 ;
        RECT 90.875 -190.665 91.045 -189.810 ;
        RECT 91.365 -190.580 91.535 -189.625 ;
        RECT 91.820 -189.825 92.060 -189.080 ;
        RECT 89.945 -190.800 90.670 -190.765 ;
        RECT 84.360 -191.005 90.670 -190.800 ;
        RECT 89.945 -191.045 90.670 -191.005 ;
        RECT 91.345 -190.835 91.555 -190.580 ;
        RECT 91.855 -190.665 92.025 -189.825 ;
        RECT 92.345 -190.580 92.515 -189.625 ;
        RECT 92.325 -190.835 92.535 -190.580 ;
        RECT 91.345 -191.045 95.275 -190.835 ;
        RECT 94.580 -191.135 95.275 -191.045 ;
        RECT 91.590 -191.260 92.315 -191.240 ;
        RECT 83.150 -191.465 92.315 -191.260 ;
        RECT 91.590 -191.520 92.315 -191.465 ;
        RECT 93.190 -191.680 93.915 -191.400 ;
        RECT 93.190 -191.705 93.490 -191.680 ;
        RECT 81.885 -191.910 93.490 -191.705 ;
        RECT 94.580 -192.045 94.790 -191.135 ;
        RECT 90.855 -192.275 93.100 -192.090 ;
        RECT 90.855 -192.530 91.060 -192.275 ;
        RECT 91.910 -192.495 92.120 -192.275 ;
        RECT -11.610 -195.005 -8.470 -194.835 ;
        RECT -62.610 -195.640 -61.835 -195.630 ;
        RECT -62.510 -195.680 -61.835 -195.640 ;
        RECT -64.985 -195.930 -62.240 -195.920 ;
        RECT -60.185 -195.930 -59.815 -195.800 ;
        RECT -64.985 -195.950 -59.815 -195.930 ;
        RECT -77.285 -196.660 -76.245 -196.650 ;
        RECT -66.460 -197.230 -66.290 -195.950 ;
        RECT -65.970 -196.990 -65.800 -195.950 ;
        RECT -65.480 -197.230 -65.310 -195.950 ;
        RECT -64.990 -196.120 -59.815 -195.950 ;
        RECT -59.250 -196.015 -55.325 -195.585 ;
        RECT -6.785 -195.670 42.510 -194.365 ;
        RECT 90.875 -195.485 91.045 -192.530 ;
        RECT 91.935 -195.485 92.105 -192.495 ;
        RECT 92.425 -195.455 92.595 -192.445 ;
        RECT 92.890 -192.500 93.100 -192.275 ;
        RECT 93.950 -192.255 94.790 -192.045 ;
        RECT -64.990 -196.990 -64.820 -196.120 ;
        RECT -62.245 -196.125 -59.815 -196.120 ;
        RECT -62.245 -196.130 -61.890 -196.125 ;
        RECT -60.185 -196.155 -59.815 -196.125 ;
        RECT -67.160 -197.660 -62.470 -197.230 ;
        RECT -81.980 -197.950 -80.640 -197.715 ;
        RECT -118.995 -198.880 -80.640 -197.950 ;
        RECT -62.900 -198.065 -62.470 -197.660 ;
        RECT -62.085 -197.880 -61.915 -196.340 ;
        RECT -61.595 -197.880 -61.425 -196.340 ;
        RECT -61.105 -197.880 -60.935 -196.340 ;
        RECT -60.615 -197.880 -60.445 -196.340 ;
        RECT -60.125 -197.880 -59.955 -196.340 ;
        RECT -61.600 -198.065 -61.425 -197.880 ;
        RECT -58.030 -198.050 -57.725 -196.015 ;
        RECT -59.975 -198.065 -57.725 -198.050 ;
        RECT -62.900 -198.355 -57.725 -198.065 ;
        RECT -62.900 -198.495 -59.575 -198.355 ;
        RECT -129.885 -214.935 -121.675 -214.360 ;
        RECT -129.885 -215.635 -128.195 -214.935 ;
        RECT -118.640 -220.870 -117.710 -198.880 ;
        RECT -81.980 -199.040 -80.640 -198.880 ;
        RECT -64.480 -199.460 -61.340 -199.290 ;
        RECT -71.715 -199.575 -71.545 -199.555 ;
        RECT -71.745 -200.840 -71.515 -199.575 ;
        RECT -70.735 -200.515 -70.565 -199.555 ;
        RECT -69.755 -200.515 -69.585 -199.555 ;
        RECT -67.530 -199.575 -67.360 -199.555 ;
        RECT -68.635 -199.985 -68.350 -199.665 ;
        RECT -69.350 -200.230 -68.350 -199.985 ;
        RECT -70.765 -200.840 -70.535 -200.515 ;
        RECT -69.785 -200.840 -69.555 -200.515 ;
        RECT -71.745 -200.880 -69.555 -200.840 ;
        RECT -69.350 -200.880 -69.120 -200.230 ;
        RECT -68.635 -200.485 -68.350 -200.230 ;
        RECT -72.765 -201.065 -71.925 -200.915 ;
        RECT -72.800 -201.285 -71.925 -201.065 ;
        RECT -71.745 -201.070 -69.120 -200.880 ;
        RECT -67.560 -200.840 -67.330 -199.575 ;
        RECT -66.550 -200.515 -66.380 -199.555 ;
        RECT -65.570 -200.515 -65.400 -199.555 ;
        RECT -64.480 -199.685 -64.300 -199.460 ;
        RECT -66.580 -200.840 -66.350 -200.515 ;
        RECT -65.600 -200.840 -65.370 -200.515 ;
        RECT -67.560 -200.880 -65.370 -200.840 ;
        RECT -65.095 -200.760 -64.725 -199.920 ;
        RECT -64.475 -200.055 -64.305 -199.685 ;
        RECT -65.095 -200.880 -64.730 -200.760 ;
        RECT -68.580 -200.970 -67.740 -200.915 ;
        RECT -68.755 -200.975 -67.740 -200.970 ;
        RECT -72.800 -203.145 -72.560 -201.285 ;
        RECT -72.205 -202.250 -72.035 -201.455 ;
        RECT -71.745 -201.535 -71.515 -201.070 ;
        RECT -71.715 -201.995 -71.545 -201.535 ;
        RECT -71.225 -202.250 -71.055 -201.455 ;
        RECT -70.765 -201.535 -70.535 -201.070 ;
        RECT -69.785 -201.230 -69.120 -201.070 ;
        RECT -70.735 -201.995 -70.565 -201.535 ;
        RECT -70.245 -202.250 -70.075 -201.455 ;
        RECT -69.785 -201.535 -69.555 -201.230 ;
        RECT -68.940 -201.285 -67.740 -200.975 ;
        RECT -67.560 -201.070 -64.730 -200.880 ;
        RECT -69.755 -201.995 -69.585 -201.535 ;
        RECT -68.940 -202.005 -68.640 -201.285 ;
        RECT -68.020 -202.250 -67.850 -201.455 ;
        RECT -67.560 -201.535 -67.330 -201.070 ;
        RECT -67.530 -201.995 -67.360 -201.535 ;
        RECT -67.040 -202.250 -66.870 -201.455 ;
        RECT -66.580 -201.535 -66.350 -201.070 ;
        RECT -65.600 -201.230 -64.730 -201.070 ;
        RECT -64.505 -200.790 -64.270 -200.055 ;
        RECT -63.985 -200.090 -63.815 -199.630 ;
        RECT -63.500 -199.735 -63.290 -199.460 ;
        RECT -63.990 -200.350 -63.810 -200.090 ;
        RECT -63.495 -200.170 -63.325 -199.735 ;
        RECT -63.005 -200.080 -62.835 -199.630 ;
        RECT -62.530 -199.740 -62.320 -199.460 ;
        RECT -63.005 -200.170 -62.820 -200.080 ;
        RECT -62.515 -200.170 -62.345 -199.740 ;
        RECT -62.025 -200.080 -61.855 -199.630 ;
        RECT -61.550 -199.715 -61.340 -199.460 ;
        RECT -50.980 -199.460 -47.840 -199.290 ;
        RECT -58.215 -199.575 -58.045 -199.555 ;
        RECT -63.000 -200.350 -62.820 -200.170 ;
        RECT -62.030 -200.350 -61.850 -200.080 ;
        RECT -61.535 -200.170 -61.365 -199.715 ;
        RECT -61.045 -200.130 -60.875 -199.630 ;
        RECT -61.060 -200.350 -60.850 -200.130 ;
        RECT -63.990 -200.520 -60.850 -200.350 ;
        RECT -64.505 -201.160 -63.645 -200.790 ;
        RECT -61.725 -201.055 -60.850 -200.520 ;
        RECT -58.245 -200.840 -58.015 -199.575 ;
        RECT -57.235 -200.515 -57.065 -199.555 ;
        RECT -56.255 -200.515 -56.085 -199.555 ;
        RECT -54.030 -199.575 -53.860 -199.555 ;
        RECT -55.135 -199.925 -54.850 -199.665 ;
        RECT -55.875 -200.235 -54.850 -199.925 ;
        RECT -57.265 -200.840 -57.035 -200.515 ;
        RECT -56.285 -200.840 -56.055 -200.515 ;
        RECT -58.245 -200.880 -56.055 -200.840 ;
        RECT -55.875 -200.880 -55.565 -200.235 ;
        RECT -55.135 -200.485 -54.850 -200.235 ;
        RECT -59.265 -200.950 -58.425 -200.915 ;
        RECT -66.550 -201.995 -66.380 -201.535 ;
        RECT -66.060 -202.250 -65.890 -201.455 ;
        RECT -65.600 -201.535 -65.370 -201.230 ;
        RECT -65.570 -201.995 -65.400 -201.535 ;
        RECT -64.505 -201.835 -64.270 -201.160 ;
        RECT -61.725 -201.355 -60.395 -201.055 ;
        RECT -59.375 -201.250 -58.425 -200.950 ;
        RECT -59.265 -201.285 -58.425 -201.250 ;
        RECT -58.245 -201.070 -55.565 -200.880 ;
        RECT -54.060 -200.840 -53.830 -199.575 ;
        RECT -53.050 -200.515 -52.880 -199.555 ;
        RECT -52.070 -200.515 -51.900 -199.555 ;
        RECT -50.980 -199.685 -50.800 -199.460 ;
        RECT -53.080 -200.840 -52.850 -200.515 ;
        RECT -52.100 -200.840 -51.870 -200.515 ;
        RECT -54.060 -200.880 -51.870 -200.840 ;
        RECT -51.595 -200.760 -51.225 -199.920 ;
        RECT -50.975 -200.055 -50.805 -199.685 ;
        RECT -51.595 -200.880 -51.230 -200.760 ;
        RECT -55.080 -200.970 -54.240 -200.915 ;
        RECT -64.005 -201.525 -60.850 -201.355 ;
        RECT -64.005 -201.730 -63.800 -201.525 ;
        RECT -64.475 -202.185 -64.305 -201.835 ;
        RECT -72.250 -202.590 -65.395 -202.250 ;
        RECT -64.500 -202.475 -64.280 -202.185 ;
        RECT -63.985 -202.245 -63.815 -201.730 ;
        RECT -63.495 -202.130 -63.325 -201.705 ;
        RECT -63.015 -201.770 -62.810 -201.525 ;
        RECT -63.520 -202.475 -63.300 -202.130 ;
        RECT -63.005 -202.245 -62.835 -201.770 ;
        RECT -62.515 -202.130 -62.345 -201.705 ;
        RECT -62.045 -201.770 -61.840 -201.525 ;
        RECT -61.060 -201.560 -60.850 -201.525 ;
        RECT -62.540 -202.475 -62.320 -202.130 ;
        RECT -62.025 -202.245 -61.855 -201.770 ;
        RECT -61.535 -202.185 -61.365 -201.705 ;
        RECT -61.060 -201.775 -60.855 -201.560 ;
        RECT -61.555 -202.475 -61.335 -202.185 ;
        RECT -61.045 -202.245 -60.875 -201.775 ;
        RECT -58.705 -202.250 -58.535 -201.455 ;
        RECT -58.245 -201.535 -58.015 -201.070 ;
        RECT -58.215 -201.995 -58.045 -201.535 ;
        RECT -57.725 -202.250 -57.555 -201.455 ;
        RECT -57.265 -201.535 -57.035 -201.070 ;
        RECT -56.285 -201.230 -55.565 -201.070 ;
        RECT -57.235 -201.995 -57.065 -201.535 ;
        RECT -56.745 -202.250 -56.575 -201.455 ;
        RECT -56.285 -201.535 -56.055 -201.230 ;
        RECT -55.380 -201.285 -54.240 -200.970 ;
        RECT -54.060 -201.070 -51.230 -200.880 ;
        RECT -56.255 -201.995 -56.085 -201.535 ;
        RECT -55.380 -202.080 -55.080 -201.285 ;
        RECT -54.520 -202.250 -54.350 -201.455 ;
        RECT -54.060 -201.535 -53.830 -201.070 ;
        RECT -54.030 -201.995 -53.860 -201.535 ;
        RECT -53.540 -202.250 -53.370 -201.455 ;
        RECT -53.080 -201.535 -52.850 -201.070 ;
        RECT -52.100 -201.230 -51.230 -201.070 ;
        RECT -51.005 -200.790 -50.770 -200.055 ;
        RECT -50.485 -200.090 -50.315 -199.630 ;
        RECT -50.000 -199.735 -49.790 -199.460 ;
        RECT -50.490 -200.350 -50.310 -200.090 ;
        RECT -49.995 -200.170 -49.825 -199.735 ;
        RECT -49.505 -200.080 -49.335 -199.630 ;
        RECT -49.030 -199.740 -48.820 -199.460 ;
        RECT -49.505 -200.170 -49.320 -200.080 ;
        RECT -49.015 -200.170 -48.845 -199.740 ;
        RECT -48.525 -200.080 -48.355 -199.630 ;
        RECT -48.050 -199.715 -47.840 -199.460 ;
        RECT -39.720 -199.470 -38.520 -199.300 ;
        RECT -49.500 -200.350 -49.320 -200.170 ;
        RECT -48.530 -200.350 -48.350 -200.080 ;
        RECT -48.035 -200.170 -47.865 -199.715 ;
        RECT -47.545 -200.130 -47.375 -199.630 ;
        RECT -47.560 -200.350 -47.350 -200.130 ;
        RECT -50.490 -200.520 -47.350 -200.350 ;
        RECT -51.005 -201.160 -50.145 -200.790 ;
        RECT -48.225 -201.065 -47.350 -200.520 ;
        RECT -53.050 -201.995 -52.880 -201.535 ;
        RECT -52.560 -202.250 -52.390 -201.455 ;
        RECT -52.100 -201.535 -51.870 -201.230 ;
        RECT -52.070 -201.995 -51.900 -201.535 ;
        RECT -51.005 -201.835 -50.770 -201.160 ;
        RECT -48.225 -201.355 -46.975 -201.065 ;
        RECT -50.505 -201.365 -46.975 -201.355 ;
        RECT -50.505 -201.525 -47.350 -201.365 ;
        RECT -50.505 -201.730 -50.300 -201.525 ;
        RECT -50.975 -202.185 -50.805 -201.835 ;
        RECT -71.010 -202.790 -70.455 -202.590 ;
        RECT -71.065 -202.830 -70.380 -202.790 ;
        RECT -66.955 -202.830 -66.400 -202.590 ;
        RECT -64.500 -202.645 -61.335 -202.475 ;
        RECT -58.750 -202.260 -56.080 -202.250 ;
        RECT -54.565 -202.260 -51.895 -202.250 ;
        RECT -58.750 -202.590 -51.895 -202.260 ;
        RECT -51.000 -202.475 -50.780 -202.185 ;
        RECT -50.485 -202.245 -50.315 -201.730 ;
        RECT -49.995 -202.130 -49.825 -201.705 ;
        RECT -49.515 -201.770 -49.310 -201.525 ;
        RECT -50.020 -202.475 -49.800 -202.130 ;
        RECT -49.505 -202.245 -49.335 -201.770 ;
        RECT -49.015 -202.130 -48.845 -201.705 ;
        RECT -48.545 -201.770 -48.340 -201.525 ;
        RECT -47.560 -201.560 -47.350 -201.525 ;
        RECT -49.040 -202.475 -48.820 -202.130 ;
        RECT -48.525 -202.245 -48.355 -201.770 ;
        RECT -48.035 -202.185 -47.865 -201.705 ;
        RECT -47.560 -201.775 -47.355 -201.560 ;
        RECT -48.055 -202.475 -47.835 -202.185 ;
        RECT -47.545 -202.245 -47.375 -201.775 ;
        RECT -57.965 -202.820 -57.410 -202.590 ;
        RECT -57.050 -202.600 -54.450 -202.590 ;
        RECT -58.080 -202.830 -57.395 -202.820 ;
        RECT -53.575 -202.830 -53.020 -202.590 ;
        RECT -51.000 -202.645 -47.835 -202.475 ;
        RECT -40.750 -202.610 -40.580 -199.640 ;
        RECT -39.720 -199.690 -39.510 -199.470 ;
        RECT -44.890 -202.830 -44.230 -202.820 ;
        RECT -71.150 -203.025 -44.225 -202.830 ;
        RECT -71.065 -203.090 -70.380 -203.025 ;
        RECT -58.080 -203.120 -57.395 -203.025 ;
        RECT -44.890 -203.120 -44.230 -203.025 ;
        RECT -72.805 -203.830 -72.505 -203.145 ;
        RECT -60.255 -203.290 -59.570 -203.235 ;
        RECT -55.525 -203.290 -54.865 -203.240 ;
        RECT -71.150 -203.485 -42.500 -203.290 ;
        RECT -60.255 -203.535 -59.570 -203.485 ;
        RECT -55.525 -203.540 -54.865 -203.485 ;
        RECT -69.120 -203.720 -68.460 -203.680 ;
        RECT -46.505 -203.720 -45.845 -203.670 ;
        RECT -102.050 -204.445 -100.830 -204.255 ;
        RECT -107.600 -204.800 -105.285 -204.630 ;
        RECT -109.100 -207.935 -108.930 -204.980 ;
        RECT -109.120 -208.190 -108.915 -207.935 ;
        RECT -108.040 -207.970 -107.870 -204.980 ;
        RECT -107.600 -205.010 -107.335 -204.800 ;
        RECT -108.065 -208.190 -107.855 -207.970 ;
        RECT -107.550 -208.020 -107.380 -205.010 ;
        RECT -107.060 -207.965 -106.890 -204.980 ;
        RECT -106.555 -205.010 -106.275 -204.800 ;
        RECT -107.085 -208.190 -106.875 -207.965 ;
        RECT -106.495 -208.020 -106.325 -205.010 ;
        RECT -106.005 -207.930 -105.835 -204.980 ;
        RECT -105.565 -205.010 -105.285 -204.800 ;
        RECT -109.120 -208.375 -106.875 -208.190 ;
        RECT -106.025 -208.210 -105.815 -207.930 ;
        RECT -105.515 -208.020 -105.345 -205.010 ;
        RECT -103.070 -206.640 -102.900 -204.625 ;
        RECT -102.050 -204.765 -101.820 -204.445 ;
        RECT -103.075 -206.835 -102.895 -206.640 ;
        RECT -102.015 -206.665 -101.845 -204.765 ;
        RECT -101.525 -206.615 -101.355 -204.625 ;
        RECT -101.060 -204.765 -100.830 -204.445 ;
        RECT -97.525 -204.450 -96.305 -204.260 ;
        RECT -101.035 -206.435 -100.865 -204.765 ;
        RECT -101.560 -206.835 -101.335 -206.615 ;
        RECT -103.075 -207.015 -101.335 -206.835 ;
        RECT -101.050 -207.595 -100.800 -206.435 ;
        RECT -98.545 -206.645 -98.375 -204.630 ;
        RECT -97.525 -204.770 -97.295 -204.450 ;
        RECT -99.880 -207.250 -99.590 -206.775 ;
        RECT -98.550 -206.840 -98.370 -206.645 ;
        RECT -97.490 -206.670 -97.320 -204.770 ;
        RECT -97.000 -206.620 -96.830 -204.630 ;
        RECT -96.535 -204.770 -96.305 -204.450 ;
        RECT -87.970 -204.640 -80.585 -204.075 ;
        RECT -96.510 -206.440 -96.340 -204.770 ;
        RECT -92.125 -206.115 -89.880 -206.025 ;
        RECT -87.970 -206.115 -87.665 -204.640 ;
        RECT -84.335 -205.230 -84.100 -204.640 ;
        RECT -94.685 -206.420 -87.665 -206.115 ;
        RECT -97.035 -206.840 -96.810 -206.620 ;
        RECT -98.550 -207.020 -96.810 -206.840 ;
        RECT -97.900 -207.250 -97.185 -207.215 ;
        RECT -99.880 -207.430 -97.185 -207.250 ;
        RECT -99.880 -207.460 -99.590 -207.430 ;
        RECT -97.900 -207.515 -97.185 -207.430 ;
        RECT -104.085 -207.690 -103.795 -207.625 ;
        RECT -103.540 -207.690 -102.810 -207.610 ;
        RECT -101.050 -207.660 -100.320 -207.595 ;
        RECT -96.525 -207.600 -96.275 -206.440 ;
        RECT -104.085 -207.870 -102.810 -207.690 ;
        RECT -101.330 -207.705 -100.320 -207.660 ;
        RECT -106.025 -208.420 -105.185 -208.210 ;
        RECT -104.085 -208.310 -103.795 -207.870 ;
        RECT -103.540 -207.910 -102.810 -207.870 ;
        RECT -102.605 -207.885 -100.320 -207.705 ;
        RECT -99.495 -207.695 -99.205 -207.635 ;
        RECT -99.015 -207.695 -98.285 -207.615 ;
        RECT -96.525 -207.665 -95.665 -207.600 ;
        RECT -99.495 -207.875 -98.285 -207.695 ;
        RECT -96.805 -207.710 -95.665 -207.665 ;
        RECT -105.395 -209.340 -105.185 -208.420 ;
        RECT -103.070 -208.880 -102.900 -208.085 ;
        RECT -102.605 -208.130 -102.380 -207.885 ;
        RECT -105.440 -209.420 -104.755 -209.340 ;
        RECT -108.630 -209.630 -104.755 -209.420 ;
        RECT -109.100 -210.655 -108.930 -209.800 ;
        RECT -108.630 -209.885 -108.420 -209.630 ;
        RECT -109.125 -211.300 -108.885 -210.655 ;
        RECT -108.610 -210.840 -108.440 -209.885 ;
        RECT -108.120 -210.640 -107.950 -209.800 ;
        RECT -107.650 -209.885 -107.440 -209.630 ;
        RECT -103.090 -209.640 -102.870 -208.880 ;
        RECT -102.580 -209.125 -102.410 -208.130 ;
        RECT -102.090 -208.885 -101.920 -208.085 ;
        RECT -99.495 -208.320 -99.205 -207.875 ;
        RECT -99.015 -207.915 -98.285 -207.875 ;
        RECT -98.080 -207.890 -95.665 -207.710 ;
        RECT -98.545 -208.885 -98.375 -208.090 ;
        RECT -98.080 -208.135 -97.855 -207.890 ;
        RECT -102.120 -209.640 -101.900 -208.885 ;
        RECT -103.735 -209.815 -100.750 -209.640 ;
        RECT -98.565 -209.645 -98.345 -208.885 ;
        RECT -98.055 -209.130 -97.885 -208.135 ;
        RECT -97.565 -208.890 -97.395 -208.090 ;
        RECT -94.685 -208.210 -94.380 -206.420 ;
        RECT -91.540 -206.590 -91.365 -206.420 ;
        RECT -92.025 -208.130 -91.855 -206.590 ;
        RECT -91.535 -208.130 -91.365 -206.590 ;
        RECT -91.045 -208.130 -90.875 -206.590 ;
        RECT -90.555 -208.130 -90.385 -206.590 ;
        RECT -90.065 -208.130 -89.895 -206.590 ;
        RECT -96.620 -208.515 -94.380 -208.210 ;
        RECT -92.185 -208.345 -91.830 -208.340 ;
        RECT -90.125 -208.345 -89.755 -208.315 ;
        RECT -92.185 -208.350 -89.755 -208.345 ;
        RECT -97.595 -209.645 -97.375 -208.890 ;
        RECT -96.620 -209.645 -96.315 -208.515 ;
        RECT -93.315 -208.540 -89.755 -208.350 ;
        RECT -87.970 -208.455 -87.665 -206.420 ;
        RECT -84.300 -206.700 -84.130 -205.230 ;
        RECT -83.810 -206.620 -83.640 -205.160 ;
        RECT -83.355 -205.235 -83.120 -204.640 ;
        RECT -84.845 -206.930 -84.070 -206.870 ;
        RECT -85.030 -207.100 -84.070 -206.930 ;
        RECT -84.845 -207.145 -84.070 -207.100 ;
        RECT -83.840 -206.970 -83.615 -206.620 ;
        RECT -83.320 -206.700 -83.150 -205.235 ;
        RECT -82.145 -205.285 -81.910 -204.640 ;
        RECT -82.110 -206.700 -81.940 -205.285 ;
        RECT -81.620 -206.655 -81.450 -205.160 ;
        RECT -72.800 -205.620 -72.560 -203.830 ;
        RECT -71.150 -203.915 -45.845 -203.720 ;
        RECT -69.120 -203.980 -68.460 -203.915 ;
        RECT -46.505 -203.970 -45.845 -203.915 ;
        RECT -42.695 -203.830 -42.500 -203.485 ;
        RECT -40.790 -203.830 -40.575 -202.610 ;
        RECT -39.690 -202.680 -39.520 -199.690 ;
        RECT -39.200 -202.580 -39.030 -199.640 ;
        RECT -38.730 -199.680 -38.520 -199.470 ;
        RECT -39.220 -202.850 -39.010 -202.580 ;
        RECT -38.710 -202.590 -38.540 -199.680 ;
        RECT -37.655 -202.560 -37.485 -199.640 ;
        RECT -6.785 -199.960 -5.295 -195.670 ;
        RECT 1.260 -199.960 2.565 -195.670 ;
        RECT 5.445 -199.960 6.750 -195.670 ;
        RECT 10.645 -199.960 11.950 -195.670 ;
        RECT 17.935 -199.960 19.240 -195.670 ;
        RECT 24.005 -199.960 25.310 -195.670 ;
        RECT 33.735 -199.960 35.040 -195.670 ;
        RECT 41.205 -199.960 42.510 -195.670 ;
        RECT 92.375 -195.665 92.640 -195.455 ;
        RECT 92.915 -195.485 93.085 -192.500 ;
        RECT 93.480 -195.455 93.650 -192.445 ;
        RECT 93.950 -192.535 94.160 -192.255 ;
        RECT 93.420 -195.665 93.700 -195.455 ;
        RECT 93.970 -195.485 94.140 -192.535 ;
        RECT 94.460 -195.455 94.630 -192.445 ;
        RECT 94.410 -195.665 94.690 -195.455 ;
        RECT 92.375 -195.835 94.690 -195.665 ;
        RECT -25.110 -200.795 -21.970 -200.625 ;
        RECT -32.345 -200.910 -32.175 -200.890 ;
        RECT -32.375 -202.175 -32.145 -200.910 ;
        RECT -31.365 -201.850 -31.195 -200.890 ;
        RECT -30.385 -201.850 -30.215 -200.890 ;
        RECT -28.160 -200.910 -27.990 -200.890 ;
        RECT -29.265 -201.320 -28.980 -201.000 ;
        RECT -29.980 -201.565 -28.980 -201.320 ;
        RECT -31.395 -202.175 -31.165 -201.850 ;
        RECT -30.415 -202.175 -30.185 -201.850 ;
        RECT -32.375 -202.215 -30.185 -202.175 ;
        RECT -29.980 -202.215 -29.750 -201.565 ;
        RECT -29.265 -201.820 -28.980 -201.565 ;
        RECT -33.395 -202.400 -32.555 -202.250 ;
        RECT -39.715 -203.045 -39.010 -202.850 ;
        RECT -38.735 -202.855 -38.525 -202.590 ;
        RECT -37.675 -202.855 -37.465 -202.560 ;
        RECT -38.735 -203.035 -37.465 -202.855 ;
        RECT -33.430 -202.620 -32.555 -202.400 ;
        RECT -32.375 -202.405 -29.750 -202.215 ;
        RECT -28.190 -202.175 -27.960 -200.910 ;
        RECT -27.180 -201.850 -27.010 -200.890 ;
        RECT -26.200 -201.850 -26.030 -200.890 ;
        RECT -25.110 -201.020 -24.930 -200.795 ;
        RECT -27.210 -202.175 -26.980 -201.850 ;
        RECT -26.230 -202.175 -26.000 -201.850 ;
        RECT -28.190 -202.215 -26.000 -202.175 ;
        RECT -25.725 -202.095 -25.355 -201.255 ;
        RECT -25.105 -201.390 -24.935 -201.020 ;
        RECT -25.725 -202.215 -25.360 -202.095 ;
        RECT -29.210 -202.305 -28.370 -202.250 ;
        RECT -29.385 -202.310 -28.370 -202.305 ;
        RECT -39.715 -203.105 -39.500 -203.045 ;
        RECT -40.405 -203.380 -39.500 -203.105 ;
        RECT -39.715 -203.730 -39.500 -203.380 ;
        RECT -39.065 -203.265 -38.290 -203.215 ;
        RECT -36.500 -203.265 -35.840 -203.005 ;
        RECT -39.065 -203.445 -35.840 -203.265 ;
        RECT -39.065 -203.490 -38.290 -203.445 ;
        RECT -42.695 -204.030 -39.905 -203.830 ;
        RECT -39.715 -203.930 -37.945 -203.730 ;
        RECT -42.695 -204.045 -40.145 -204.030 ;
        RECT -72.210 -204.490 -69.540 -204.150 ;
        RECT -67.555 -204.265 -64.390 -204.095 ;
        RECT -72.205 -205.205 -72.035 -204.745 ;
        RECT -72.235 -205.510 -72.005 -205.205 ;
        RECT -71.715 -205.285 -71.545 -204.490 ;
        RECT -71.225 -205.205 -71.055 -204.745 ;
        RECT -72.385 -205.620 -72.005 -205.510 ;
        RECT -72.800 -205.670 -72.005 -205.620 ;
        RECT -71.255 -205.670 -71.025 -205.205 ;
        RECT -70.735 -205.285 -70.565 -204.490 ;
        RECT -70.245 -205.205 -70.075 -204.745 ;
        RECT -70.275 -205.670 -70.045 -205.205 ;
        RECT -69.755 -205.285 -69.585 -204.490 ;
        RECT -68.015 -204.965 -67.845 -204.495 ;
        RECT -67.555 -204.555 -67.335 -204.265 ;
        RECT -68.035 -205.180 -67.830 -204.965 ;
        RECT -67.525 -205.035 -67.355 -204.555 ;
        RECT -67.035 -204.970 -66.865 -204.495 ;
        RECT -66.570 -204.610 -66.350 -204.265 ;
        RECT -68.040 -205.215 -67.830 -205.180 ;
        RECT -67.050 -205.215 -66.845 -204.970 ;
        RECT -66.545 -205.035 -66.375 -204.610 ;
        RECT -66.055 -204.970 -65.885 -204.495 ;
        RECT -65.590 -204.610 -65.370 -204.265 ;
        RECT -66.080 -205.215 -65.875 -204.970 ;
        RECT -65.565 -205.035 -65.395 -204.610 ;
        RECT -65.075 -205.010 -64.905 -204.495 ;
        RECT -64.610 -204.555 -64.390 -204.265 ;
        RECT -63.495 -204.490 -56.040 -204.150 ;
        RECT -54.055 -204.265 -50.890 -204.095 ;
        RECT -64.585 -204.905 -64.415 -204.555 ;
        RECT -65.090 -205.215 -64.885 -205.010 ;
        RECT -68.040 -205.385 -64.885 -205.215 ;
        RECT -72.800 -205.805 -70.045 -205.670 ;
        RECT -72.795 -205.815 -70.045 -205.805 ;
        RECT -72.385 -205.860 -70.045 -205.815 ;
        RECT -69.865 -205.530 -69.025 -205.455 ;
        RECT -68.040 -205.530 -67.165 -205.385 ;
        RECT -69.865 -205.795 -67.165 -205.530 ;
        RECT -64.620 -205.580 -64.385 -204.905 ;
        RECT -63.490 -205.205 -63.320 -204.745 ;
        RECT -63.520 -205.510 -63.290 -205.205 ;
        RECT -63.000 -205.285 -62.830 -204.490 ;
        RECT -62.510 -205.205 -62.340 -204.745 ;
        RECT -69.865 -205.825 -69.025 -205.795 ;
        RECT -72.235 -205.900 -70.045 -205.860 ;
        RECT -72.235 -206.225 -72.005 -205.900 ;
        RECT -71.255 -206.225 -71.025 -205.900 ;
        RECT -81.640 -206.855 -81.420 -206.655 ;
        RECT -77.180 -206.855 -76.495 -206.505 ;
        RECT -81.640 -206.870 -76.495 -206.855 ;
        RECT -83.840 -207.170 -82.070 -206.970 ;
        RECT -81.880 -207.070 -76.495 -206.870 ;
        RECT -85.520 -207.455 -85.170 -207.445 ;
        RECT -83.495 -207.455 -82.720 -207.410 ;
        RECT -85.520 -207.635 -82.720 -207.455 ;
        RECT -93.315 -208.550 -92.180 -208.540 ;
        RECT -90.125 -208.670 -89.755 -208.540 ;
        RECT -95.045 -208.840 -94.460 -208.765 ;
        RECT -92.450 -208.830 -91.775 -208.790 ;
        RECT -92.550 -208.840 -91.775 -208.830 ;
        RECT -95.045 -209.020 -91.775 -208.840 ;
        RECT -89.190 -208.885 -86.115 -208.455 ;
        RECT -95.045 -209.380 -94.460 -209.020 ;
        RECT -92.550 -209.030 -91.775 -209.020 ;
        RECT -92.450 -209.060 -91.775 -209.030 ;
        RECT -91.535 -208.945 -89.440 -208.905 ;
        RECT -91.535 -209.095 -89.385 -208.945 ;
        RECT -99.210 -209.815 -96.225 -209.645 ;
        RECT -108.155 -211.300 -107.915 -210.640 ;
        RECT -107.630 -210.840 -107.460 -209.885 ;
        RECT -106.510 -210.090 -96.225 -209.815 ;
        RECT -106.510 -210.395 -97.305 -210.090 ;
        RECT -106.510 -211.300 -105.930 -210.395 ;
        RECT -91.535 -210.815 -91.365 -209.095 ;
        RECT -90.555 -210.815 -90.385 -209.095 ;
        RECT -89.690 -209.840 -89.385 -209.095 ;
        RECT -88.490 -209.665 -88.320 -208.885 ;
        RECT -88.000 -209.665 -87.830 -209.125 ;
        RECT -87.510 -209.665 -87.340 -208.885 ;
        RECT -87.020 -209.665 -86.850 -209.125 ;
        RECT -85.520 -209.610 -85.170 -207.635 ;
        RECT -83.495 -207.685 -82.720 -207.635 ;
        RECT -82.285 -207.520 -82.070 -207.170 ;
        RECT -82.285 -207.795 -81.380 -207.520 ;
        RECT -82.285 -207.855 -82.070 -207.795 ;
        RECT -84.320 -208.045 -83.050 -207.865 ;
        RECT -84.320 -208.340 -84.110 -208.045 ;
        RECT -83.260 -208.310 -83.050 -208.045 ;
        RECT -82.775 -208.050 -82.070 -207.855 ;
        RECT -89.080 -209.840 -88.715 -209.810 ;
        RECT -89.690 -209.905 -88.715 -209.840 ;
        RECT -89.580 -210.045 -88.715 -209.905 ;
        RECT -89.080 -210.110 -88.715 -210.045 ;
        RECT -86.530 -209.960 -85.140 -209.610 ;
        RECT -88.490 -210.820 -88.320 -210.280 ;
        RECT -87.510 -210.820 -87.340 -210.280 ;
        RECT -86.530 -210.820 -86.360 -209.960 ;
        RECT -84.300 -211.260 -84.130 -208.340 ;
        RECT -83.245 -211.220 -83.075 -208.310 ;
        RECT -82.775 -208.320 -82.565 -208.050 ;
        RECT -109.800 -211.385 -105.780 -211.300 ;
        RECT -109.800 -211.915 -105.360 -211.385 ;
        RECT -83.265 -211.430 -83.055 -211.220 ;
        RECT -82.755 -211.260 -82.585 -208.320 ;
        RECT -82.265 -211.210 -82.095 -208.220 ;
        RECT -81.210 -208.290 -80.995 -207.070 ;
        RECT -77.180 -207.335 -76.495 -207.070 ;
        RECT -72.205 -207.185 -72.035 -206.225 ;
        RECT -71.225 -207.185 -71.055 -206.225 ;
        RECT -70.275 -207.165 -70.045 -205.900 ;
        RECT -68.040 -206.220 -67.165 -205.795 ;
        RECT -65.245 -205.950 -64.385 -205.580 ;
        RECT -68.040 -206.390 -64.900 -206.220 ;
        RECT -68.040 -206.610 -67.830 -206.390 ;
        RECT -68.015 -207.110 -67.845 -206.610 ;
        RECT -67.525 -207.025 -67.355 -206.570 ;
        RECT -67.040 -206.660 -66.860 -206.390 ;
        RECT -66.070 -206.570 -65.890 -206.390 ;
        RECT -70.245 -207.185 -70.075 -207.165 ;
        RECT -67.550 -207.280 -67.340 -207.025 ;
        RECT -67.035 -207.110 -66.865 -206.660 ;
        RECT -66.545 -207.000 -66.375 -206.570 ;
        RECT -66.070 -206.660 -65.885 -206.570 ;
        RECT -66.570 -207.280 -66.360 -207.000 ;
        RECT -66.055 -207.110 -65.885 -206.660 ;
        RECT -65.565 -207.005 -65.395 -206.570 ;
        RECT -65.080 -206.650 -64.900 -206.390 ;
        RECT -65.600 -207.280 -65.390 -207.005 ;
        RECT -65.075 -207.110 -64.905 -206.650 ;
        RECT -64.620 -206.685 -64.385 -205.950 ;
        RECT -64.160 -205.670 -63.290 -205.510 ;
        RECT -62.540 -205.670 -62.310 -205.205 ;
        RECT -62.020 -205.285 -61.850 -204.490 ;
        RECT -61.530 -205.205 -61.360 -204.745 ;
        RECT -61.560 -205.670 -61.330 -205.205 ;
        RECT -61.040 -205.285 -60.870 -204.490 ;
        RECT -64.160 -205.860 -61.330 -205.670 ;
        RECT -61.150 -205.480 -60.310 -205.455 ;
        RECT -60.010 -205.480 -59.710 -205.115 ;
        RECT -61.150 -205.770 -59.710 -205.480 ;
        RECT -59.435 -205.565 -59.135 -204.990 ;
        RECT -58.705 -205.205 -58.535 -204.745 ;
        RECT -58.735 -205.510 -58.505 -205.205 ;
        RECT -58.215 -205.285 -58.045 -204.490 ;
        RECT -57.725 -205.205 -57.555 -204.745 ;
        RECT -58.885 -205.565 -58.505 -205.510 ;
        RECT -61.150 -205.825 -60.310 -205.770 ;
        RECT -60.010 -205.775 -59.710 -205.770 ;
        RECT -59.460 -205.670 -58.505 -205.565 ;
        RECT -57.755 -205.670 -57.525 -205.205 ;
        RECT -57.235 -205.285 -57.065 -204.490 ;
        RECT -56.745 -205.205 -56.575 -204.745 ;
        RECT -56.775 -205.670 -56.545 -205.205 ;
        RECT -56.255 -205.285 -56.085 -204.490 ;
        RECT -54.530 -204.965 -54.300 -204.355 ;
        RECT -54.055 -204.555 -53.835 -204.265 ;
        RECT -54.535 -205.015 -54.300 -204.965 ;
        RECT -54.535 -205.180 -54.330 -205.015 ;
        RECT -54.025 -205.035 -53.855 -204.555 ;
        RECT -53.535 -204.970 -53.365 -204.495 ;
        RECT -53.070 -204.610 -52.850 -204.265 ;
        RECT -54.540 -205.215 -54.330 -205.180 ;
        RECT -53.550 -205.215 -53.345 -204.970 ;
        RECT -53.045 -205.035 -52.875 -204.610 ;
        RECT -52.555 -204.970 -52.385 -204.495 ;
        RECT -52.090 -204.610 -51.870 -204.265 ;
        RECT -52.580 -205.215 -52.375 -204.970 ;
        RECT -52.065 -205.035 -51.895 -204.610 ;
        RECT -51.575 -205.010 -51.405 -204.495 ;
        RECT -51.110 -204.555 -50.890 -204.265 ;
        RECT -49.995 -204.490 -42.915 -204.150 ;
        RECT -51.085 -204.905 -50.915 -204.555 ;
        RECT -51.590 -205.215 -51.385 -205.010 ;
        RECT -54.540 -205.385 -51.385 -205.215 ;
        RECT -59.460 -205.790 -56.545 -205.670 ;
        RECT -64.160 -205.980 -63.795 -205.860 ;
        RECT -64.585 -207.055 -64.415 -206.685 ;
        RECT -64.165 -206.820 -63.795 -205.980 ;
        RECT -63.520 -205.900 -61.330 -205.860 ;
        RECT -63.520 -206.225 -63.290 -205.900 ;
        RECT -62.540 -206.225 -62.310 -205.900 ;
        RECT -64.590 -207.280 -64.410 -207.055 ;
        RECT -63.490 -207.185 -63.320 -206.225 ;
        RECT -62.510 -207.185 -62.340 -206.225 ;
        RECT -61.560 -207.165 -61.330 -205.900 ;
        RECT -60.540 -206.460 -60.255 -206.255 ;
        RECT -59.460 -206.460 -59.235 -205.790 ;
        RECT -58.885 -205.860 -56.545 -205.790 ;
        RECT -56.365 -205.495 -55.525 -205.455 ;
        RECT -54.540 -205.495 -53.665 -205.385 ;
        RECT -56.365 -205.780 -53.665 -205.495 ;
        RECT -51.120 -205.580 -50.885 -204.905 ;
        RECT -49.990 -205.205 -49.820 -204.745 ;
        RECT -50.020 -205.510 -49.790 -205.205 ;
        RECT -49.500 -205.285 -49.330 -204.490 ;
        RECT -49.010 -205.205 -48.840 -204.745 ;
        RECT -56.365 -205.825 -55.525 -205.780 ;
        RECT -58.735 -205.900 -56.545 -205.860 ;
        RECT -58.735 -206.225 -58.505 -205.900 ;
        RECT -57.755 -206.225 -57.525 -205.900 ;
        RECT -60.540 -206.685 -59.235 -206.460 ;
        RECT -60.540 -207.075 -60.255 -206.685 ;
        RECT -61.530 -207.185 -61.360 -207.165 ;
        RECT -58.705 -207.185 -58.535 -206.225 ;
        RECT -57.725 -207.185 -57.555 -206.225 ;
        RECT -56.775 -207.165 -56.545 -205.900 ;
        RECT -54.540 -206.220 -53.665 -205.780 ;
        RECT -51.745 -205.950 -50.885 -205.580 ;
        RECT -54.540 -206.390 -51.400 -206.220 ;
        RECT -54.540 -206.610 -54.330 -206.390 ;
        RECT -54.515 -207.110 -54.345 -206.610 ;
        RECT -54.025 -207.025 -53.855 -206.570 ;
        RECT -53.540 -206.660 -53.360 -206.390 ;
        RECT -52.570 -206.570 -52.390 -206.390 ;
        RECT -56.745 -207.185 -56.575 -207.165 ;
        RECT -67.550 -207.450 -64.410 -207.280 ;
        RECT -54.050 -207.280 -53.840 -207.025 ;
        RECT -53.535 -207.110 -53.365 -206.660 ;
        RECT -53.045 -207.000 -52.875 -206.570 ;
        RECT -52.570 -206.660 -52.385 -206.570 ;
        RECT -53.070 -207.280 -52.860 -207.000 ;
        RECT -52.555 -207.110 -52.385 -206.660 ;
        RECT -52.065 -207.005 -51.895 -206.570 ;
        RECT -51.580 -206.650 -51.400 -206.390 ;
        RECT -52.100 -207.280 -51.890 -207.005 ;
        RECT -51.575 -207.110 -51.405 -206.650 ;
        RECT -51.120 -206.685 -50.885 -205.950 ;
        RECT -50.660 -205.670 -49.790 -205.510 ;
        RECT -49.040 -205.670 -48.810 -205.205 ;
        RECT -48.520 -205.285 -48.350 -204.490 ;
        RECT -48.030 -205.205 -47.860 -204.745 ;
        RECT -48.060 -205.670 -47.830 -205.205 ;
        RECT -47.540 -205.285 -47.370 -204.490 ;
        RECT -50.660 -205.860 -47.830 -205.670 ;
        RECT -47.650 -205.480 -46.810 -205.455 ;
        RECT -47.650 -205.540 -46.635 -205.480 ;
        RECT -46.350 -205.540 -46.050 -205.110 ;
        RECT -45.580 -205.205 -45.410 -204.745 ;
        RECT -45.610 -205.510 -45.380 -205.205 ;
        RECT -45.090 -205.285 -44.920 -204.490 ;
        RECT -44.600 -205.205 -44.430 -204.745 ;
        RECT -45.760 -205.540 -45.380 -205.510 ;
        RECT -47.650 -205.670 -45.380 -205.540 ;
        RECT -44.630 -205.670 -44.400 -205.205 ;
        RECT -44.110 -205.285 -43.940 -204.490 ;
        RECT -43.620 -205.205 -43.450 -204.745 ;
        RECT -43.650 -205.670 -43.420 -205.205 ;
        RECT -43.130 -205.285 -42.960 -204.490 ;
        RECT -42.695 -205.455 -42.500 -204.045 ;
        RECT -40.365 -204.245 -40.145 -204.045 ;
        RECT -47.650 -205.750 -43.420 -205.670 ;
        RECT -47.650 -205.770 -46.635 -205.750 ;
        RECT -46.350 -205.770 -46.050 -205.750 ;
        RECT -47.650 -205.825 -46.810 -205.770 ;
        RECT -45.760 -205.860 -43.420 -205.750 ;
        RECT -43.240 -205.825 -42.400 -205.455 ;
        RECT -40.335 -205.740 -40.165 -204.245 ;
        RECT -39.845 -205.615 -39.675 -204.200 ;
        RECT -50.660 -205.980 -50.295 -205.860 ;
        RECT -51.085 -207.055 -50.915 -206.685 ;
        RECT -50.665 -206.820 -50.295 -205.980 ;
        RECT -50.020 -205.900 -47.830 -205.860 ;
        RECT -50.020 -206.225 -49.790 -205.900 ;
        RECT -49.040 -206.225 -48.810 -205.900 ;
        RECT -51.090 -207.280 -50.910 -207.055 ;
        RECT -49.990 -207.185 -49.820 -206.225 ;
        RECT -49.010 -207.185 -48.840 -206.225 ;
        RECT -48.060 -207.165 -47.830 -205.900 ;
        RECT -45.610 -205.900 -43.420 -205.860 ;
        RECT -45.610 -206.225 -45.380 -205.900 ;
        RECT -44.630 -206.225 -44.400 -205.900 ;
        RECT -47.040 -207.075 -46.755 -206.255 ;
        RECT -48.030 -207.185 -47.860 -207.165 ;
        RECT -45.580 -207.185 -45.410 -206.225 ;
        RECT -44.600 -207.185 -44.430 -206.225 ;
        RECT -43.650 -207.165 -43.420 -205.900 ;
        RECT -39.875 -206.265 -39.640 -205.615 ;
        RECT -38.635 -205.665 -38.465 -204.200 ;
        RECT -38.170 -204.280 -37.945 -203.930 ;
        RECT -37.715 -203.800 -36.940 -203.755 ;
        RECT -35.125 -203.800 -34.415 -203.715 ;
        RECT -37.715 -203.970 -34.415 -203.800 ;
        RECT -37.715 -204.030 -36.940 -203.970 ;
        RECT -35.125 -204.035 -34.415 -203.970 ;
        RECT -38.665 -206.265 -38.430 -205.665 ;
        RECT -38.145 -205.740 -37.975 -204.280 ;
        RECT -37.655 -205.670 -37.485 -204.200 ;
        RECT -33.430 -204.480 -33.190 -202.620 ;
        RECT -32.835 -203.585 -32.665 -202.790 ;
        RECT -32.375 -202.870 -32.145 -202.405 ;
        RECT -32.345 -203.330 -32.175 -202.870 ;
        RECT -31.855 -203.585 -31.685 -202.790 ;
        RECT -31.395 -202.870 -31.165 -202.405 ;
        RECT -30.415 -202.565 -29.750 -202.405 ;
        RECT -31.365 -203.330 -31.195 -202.870 ;
        RECT -30.875 -203.585 -30.705 -202.790 ;
        RECT -30.415 -202.870 -30.185 -202.565 ;
        RECT -29.570 -202.620 -28.370 -202.310 ;
        RECT -28.190 -202.405 -25.360 -202.215 ;
        RECT -30.385 -203.330 -30.215 -202.870 ;
        RECT -29.570 -203.340 -29.270 -202.620 ;
        RECT -28.650 -203.585 -28.480 -202.790 ;
        RECT -28.190 -202.870 -27.960 -202.405 ;
        RECT -28.160 -203.330 -27.990 -202.870 ;
        RECT -27.670 -203.585 -27.500 -202.790 ;
        RECT -27.210 -202.870 -26.980 -202.405 ;
        RECT -26.230 -202.565 -25.360 -202.405 ;
        RECT -25.135 -202.125 -24.900 -201.390 ;
        RECT -24.615 -201.425 -24.445 -200.965 ;
        RECT -24.130 -201.070 -23.920 -200.795 ;
        RECT -24.620 -201.685 -24.440 -201.425 ;
        RECT -24.125 -201.505 -23.955 -201.070 ;
        RECT -23.635 -201.415 -23.465 -200.965 ;
        RECT -23.160 -201.075 -22.950 -200.795 ;
        RECT -23.635 -201.505 -23.450 -201.415 ;
        RECT -23.145 -201.505 -22.975 -201.075 ;
        RECT -22.655 -201.415 -22.485 -200.965 ;
        RECT -22.180 -201.050 -21.970 -200.795 ;
        RECT -11.610 -200.795 -8.470 -200.625 ;
        RECT -18.845 -200.910 -18.675 -200.890 ;
        RECT -23.630 -201.685 -23.450 -201.505 ;
        RECT -22.660 -201.685 -22.480 -201.415 ;
        RECT -22.165 -201.505 -21.995 -201.050 ;
        RECT -21.675 -201.465 -21.505 -200.965 ;
        RECT -21.690 -201.685 -21.480 -201.465 ;
        RECT -24.620 -201.855 -21.480 -201.685 ;
        RECT -25.135 -202.495 -24.275 -202.125 ;
        RECT -22.355 -202.390 -21.480 -201.855 ;
        RECT -18.875 -202.175 -18.645 -200.910 ;
        RECT -17.865 -201.850 -17.695 -200.890 ;
        RECT -16.885 -201.850 -16.715 -200.890 ;
        RECT -14.660 -200.910 -14.490 -200.890 ;
        RECT -15.765 -201.260 -15.480 -201.000 ;
        RECT -16.505 -201.570 -15.480 -201.260 ;
        RECT -17.895 -202.175 -17.665 -201.850 ;
        RECT -16.915 -202.175 -16.685 -201.850 ;
        RECT -18.875 -202.215 -16.685 -202.175 ;
        RECT -16.505 -202.215 -16.195 -201.570 ;
        RECT -15.765 -201.820 -15.480 -201.570 ;
        RECT -19.895 -202.285 -19.055 -202.250 ;
        RECT -27.180 -203.330 -27.010 -202.870 ;
        RECT -26.690 -203.585 -26.520 -202.790 ;
        RECT -26.230 -202.870 -26.000 -202.565 ;
        RECT -26.200 -203.330 -26.030 -202.870 ;
        RECT -25.135 -203.170 -24.900 -202.495 ;
        RECT -22.355 -202.690 -21.025 -202.390 ;
        RECT -20.005 -202.585 -19.055 -202.285 ;
        RECT -19.895 -202.620 -19.055 -202.585 ;
        RECT -18.875 -202.405 -16.195 -202.215 ;
        RECT -24.635 -202.860 -21.480 -202.690 ;
        RECT -24.635 -203.065 -24.430 -202.860 ;
        RECT -25.105 -203.520 -24.935 -203.170 ;
        RECT -32.880 -203.925 -26.025 -203.585 ;
        RECT -25.130 -203.810 -24.910 -203.520 ;
        RECT -24.615 -203.580 -24.445 -203.065 ;
        RECT -24.125 -203.465 -23.955 -203.040 ;
        RECT -23.645 -203.105 -23.440 -202.860 ;
        RECT -24.150 -203.810 -23.930 -203.465 ;
        RECT -23.635 -203.580 -23.465 -203.105 ;
        RECT -23.145 -203.465 -22.975 -203.040 ;
        RECT -22.675 -203.105 -22.470 -202.860 ;
        RECT -21.690 -202.895 -21.480 -202.860 ;
        RECT -23.170 -203.810 -22.950 -203.465 ;
        RECT -22.655 -203.580 -22.485 -203.105 ;
        RECT -22.165 -203.520 -21.995 -203.040 ;
        RECT -21.690 -203.110 -21.485 -202.895 ;
        RECT -22.185 -203.810 -21.965 -203.520 ;
        RECT -21.675 -203.580 -21.505 -203.110 ;
        RECT -19.335 -203.585 -19.165 -202.790 ;
        RECT -18.875 -202.870 -18.645 -202.405 ;
        RECT -18.845 -203.330 -18.675 -202.870 ;
        RECT -18.355 -203.585 -18.185 -202.790 ;
        RECT -17.895 -202.870 -17.665 -202.405 ;
        RECT -16.915 -202.565 -16.195 -202.405 ;
        RECT -14.690 -202.175 -14.460 -200.910 ;
        RECT -13.680 -201.850 -13.510 -200.890 ;
        RECT -12.700 -201.850 -12.530 -200.890 ;
        RECT -11.610 -201.020 -11.430 -200.795 ;
        RECT -13.710 -202.175 -13.480 -201.850 ;
        RECT -12.730 -202.175 -12.500 -201.850 ;
        RECT -14.690 -202.215 -12.500 -202.175 ;
        RECT -12.225 -202.095 -11.855 -201.255 ;
        RECT -11.605 -201.390 -11.435 -201.020 ;
        RECT -12.225 -202.215 -11.860 -202.095 ;
        RECT -14.690 -202.405 -11.860 -202.215 ;
        RECT -17.865 -203.330 -17.695 -202.870 ;
        RECT -17.375 -203.585 -17.205 -202.790 ;
        RECT -16.915 -202.870 -16.685 -202.565 ;
        RECT -16.885 -203.330 -16.715 -202.870 ;
        RECT -15.150 -203.585 -14.980 -202.790 ;
        RECT -14.690 -202.870 -14.460 -202.405 ;
        RECT -14.660 -203.330 -14.490 -202.870 ;
        RECT -14.170 -203.585 -14.000 -202.790 ;
        RECT -13.710 -202.870 -13.480 -202.405 ;
        RECT -12.730 -202.565 -11.860 -202.405 ;
        RECT -11.635 -202.125 -11.400 -201.390 ;
        RECT -11.115 -201.425 -10.945 -200.965 ;
        RECT -10.630 -201.070 -10.420 -200.795 ;
        RECT -11.120 -201.685 -10.940 -201.425 ;
        RECT -10.625 -201.505 -10.455 -201.070 ;
        RECT -10.135 -201.415 -9.965 -200.965 ;
        RECT -9.660 -201.075 -9.450 -200.795 ;
        RECT -10.135 -201.505 -9.950 -201.415 ;
        RECT -9.645 -201.505 -9.475 -201.075 ;
        RECT -9.155 -201.415 -8.985 -200.965 ;
        RECT -8.680 -201.050 -8.470 -200.795 ;
        RECT -10.130 -201.685 -9.950 -201.505 ;
        RECT -9.160 -201.685 -8.980 -201.415 ;
        RECT -8.665 -201.505 -8.495 -201.050 ;
        RECT -8.175 -201.465 -8.005 -200.965 ;
        RECT -6.785 -201.265 42.510 -199.960 ;
        RECT 71.240 -199.325 73.810 -198.510 ;
        RECT 80.040 -199.325 81.145 -199.185 ;
        RECT 71.240 -199.975 81.145 -199.325 ;
        RECT 71.240 -200.635 73.810 -199.975 ;
        RECT -8.190 -201.685 -7.980 -201.465 ;
        RECT -11.120 -201.855 -7.980 -201.685 ;
        RECT -11.635 -202.495 -10.775 -202.125 ;
        RECT -8.855 -202.400 -7.980 -201.855 ;
        RECT -13.680 -203.330 -13.510 -202.870 ;
        RECT -13.190 -203.585 -13.020 -202.790 ;
        RECT -12.730 -202.870 -12.500 -202.565 ;
        RECT -12.700 -203.330 -12.530 -202.870 ;
        RECT -11.635 -203.170 -11.400 -202.495 ;
        RECT -8.855 -202.690 -7.605 -202.400 ;
        RECT -11.135 -202.700 -7.605 -202.690 ;
        RECT -11.135 -202.860 -7.980 -202.700 ;
        RECT -11.135 -203.065 -10.930 -202.860 ;
        RECT -11.605 -203.520 -11.435 -203.170 ;
        RECT -31.640 -204.125 -31.085 -203.925 ;
        RECT -31.695 -204.165 -31.010 -204.125 ;
        RECT -27.585 -204.165 -27.030 -203.925 ;
        RECT -25.130 -203.980 -21.965 -203.810 ;
        RECT -19.380 -203.595 -16.710 -203.585 ;
        RECT -15.195 -203.595 -12.525 -203.585 ;
        RECT -19.380 -203.925 -12.525 -203.595 ;
        RECT -11.630 -203.810 -11.410 -203.520 ;
        RECT -11.115 -203.580 -10.945 -203.065 ;
        RECT -10.625 -203.465 -10.455 -203.040 ;
        RECT -10.145 -203.105 -9.940 -202.860 ;
        RECT -10.650 -203.810 -10.430 -203.465 ;
        RECT -10.135 -203.580 -9.965 -203.105 ;
        RECT -9.645 -203.465 -9.475 -203.040 ;
        RECT -9.175 -203.105 -8.970 -202.860 ;
        RECT -8.190 -202.895 -7.980 -202.860 ;
        RECT -9.670 -203.810 -9.450 -203.465 ;
        RECT -9.155 -203.580 -8.985 -203.105 ;
        RECT -8.665 -203.520 -8.495 -203.040 ;
        RECT -8.190 -203.110 -7.985 -202.895 ;
        RECT -8.685 -203.810 -8.465 -203.520 ;
        RECT -8.175 -203.580 -8.005 -203.110 ;
        RECT -18.595 -204.155 -18.040 -203.925 ;
        RECT -17.680 -203.935 -15.080 -203.925 ;
        RECT -18.710 -204.165 -18.025 -204.155 ;
        RECT -14.205 -204.165 -13.650 -203.925 ;
        RECT -11.630 -203.980 -8.465 -203.810 ;
        RECT -6.785 -204.155 -5.295 -201.265 ;
        RECT -1.555 -202.590 -0.905 -201.265 ;
        RECT -0.025 -202.590 0.625 -201.265 ;
        RECT 1.560 -202.590 2.210 -201.265 ;
        RECT 3.790 -202.590 4.440 -201.265 ;
        RECT -1.620 -202.915 4.750 -202.590 ;
        RECT -6.785 -204.165 -4.860 -204.155 ;
        RECT -31.780 -204.360 -4.855 -204.165 ;
        RECT -31.695 -204.425 -31.010 -204.360 ;
        RECT -18.710 -204.455 -18.025 -204.360 ;
        RECT -5.520 -204.455 -4.860 -204.360 ;
        RECT -33.435 -205.165 -33.135 -204.480 ;
        RECT -29.750 -205.055 -29.090 -205.015 ;
        RECT -7.135 -205.055 -6.475 -205.005 ;
        RECT -37.685 -206.265 -37.450 -205.670 ;
        RECT -35.130 -206.265 -34.605 -206.235 ;
        RECT -40.775 -206.675 -34.605 -206.265 ;
        RECT -35.130 -206.710 -34.605 -206.675 ;
        RECT -33.430 -206.955 -33.190 -205.165 ;
        RECT -31.780 -205.250 -6.475 -205.055 ;
        RECT -29.750 -205.315 -29.090 -205.250 ;
        RECT -7.135 -205.305 -6.475 -205.250 ;
        RECT -32.840 -205.825 -30.170 -205.485 ;
        RECT -28.185 -205.600 -25.020 -205.430 ;
        RECT -32.835 -206.540 -32.665 -206.080 ;
        RECT -32.865 -206.845 -32.635 -206.540 ;
        RECT -32.345 -206.620 -32.175 -205.825 ;
        RECT -31.855 -206.540 -31.685 -206.080 ;
        RECT -33.015 -206.955 -32.635 -206.845 ;
        RECT -33.430 -207.005 -32.635 -206.955 ;
        RECT -31.885 -207.005 -31.655 -206.540 ;
        RECT -31.365 -206.620 -31.195 -205.825 ;
        RECT -30.875 -206.540 -30.705 -206.080 ;
        RECT -30.905 -207.005 -30.675 -206.540 ;
        RECT -30.385 -206.620 -30.215 -205.825 ;
        RECT -28.645 -206.300 -28.475 -205.830 ;
        RECT -28.185 -205.890 -27.965 -205.600 ;
        RECT -28.665 -206.515 -28.460 -206.300 ;
        RECT -28.155 -206.370 -27.985 -205.890 ;
        RECT -27.665 -206.305 -27.495 -205.830 ;
        RECT -27.200 -205.945 -26.980 -205.600 ;
        RECT -28.670 -206.550 -28.460 -206.515 ;
        RECT -27.680 -206.550 -27.475 -206.305 ;
        RECT -27.175 -206.370 -27.005 -205.945 ;
        RECT -26.685 -206.305 -26.515 -205.830 ;
        RECT -26.220 -205.945 -26.000 -205.600 ;
        RECT -26.710 -206.550 -26.505 -206.305 ;
        RECT -26.195 -206.370 -26.025 -205.945 ;
        RECT -25.705 -206.345 -25.535 -205.830 ;
        RECT -25.240 -205.890 -25.020 -205.600 ;
        RECT -24.125 -205.825 -16.670 -205.485 ;
        RECT -14.685 -205.600 -11.520 -205.430 ;
        RECT -25.215 -206.240 -25.045 -205.890 ;
        RECT -25.720 -206.550 -25.515 -206.345 ;
        RECT -28.670 -206.720 -25.515 -206.550 ;
        RECT -33.430 -207.140 -30.675 -207.005 ;
        RECT -33.425 -207.150 -30.675 -207.140 ;
        RECT -43.620 -207.185 -43.450 -207.165 ;
        RECT -33.015 -207.195 -30.675 -207.150 ;
        RECT -30.495 -206.865 -29.655 -206.790 ;
        RECT -28.670 -206.865 -27.795 -206.720 ;
        RECT -30.495 -207.130 -27.795 -206.865 ;
        RECT -25.250 -206.915 -25.015 -206.240 ;
        RECT -24.120 -206.540 -23.950 -206.080 ;
        RECT -24.150 -206.845 -23.920 -206.540 ;
        RECT -23.630 -206.620 -23.460 -205.825 ;
        RECT -23.140 -206.540 -22.970 -206.080 ;
        RECT -30.495 -207.160 -29.655 -207.130 ;
        RECT -54.050 -207.450 -50.910 -207.280 ;
        RECT -32.865 -207.235 -30.675 -207.195 ;
        RECT -32.865 -207.560 -32.635 -207.235 ;
        RECT -31.885 -207.560 -31.655 -207.235 ;
        RECT -80.080 -207.945 -79.555 -207.585 ;
        RECT -82.275 -211.430 -82.065 -211.210 ;
        RECT -81.205 -211.260 -81.035 -208.290 ;
        RECT -83.265 -211.600 -82.065 -211.430 ;
        RECT -109.800 -212.050 -105.780 -211.915 ;
        RECT -113.370 -212.875 -113.080 -212.860 ;
        RECT -104.095 -212.875 -103.805 -212.395 ;
        RECT -113.370 -213.080 -103.805 -212.875 ;
        RECT -113.370 -213.545 -113.080 -213.080 ;
        RECT -112.800 -213.270 -112.510 -213.265 ;
        RECT -99.990 -213.270 -99.700 -212.790 ;
        RECT -112.800 -213.475 -99.700 -213.270 ;
        RECT -112.800 -213.950 -112.510 -213.475 ;
        RECT -99.525 -213.655 -99.235 -213.175 ;
        RECT -112.075 -213.860 -99.235 -213.655 ;
        RECT -112.075 -214.340 -111.785 -213.860 ;
        RECT -110.865 -214.265 -105.950 -214.110 ;
        RECT -110.865 -214.590 -104.475 -214.265 ;
        RECT -110.865 -214.685 -105.950 -214.590 ;
        RECT -110.785 -220.110 -110.615 -215.530 ;
        RECT -110.295 -216.570 -110.125 -214.685 ;
        RECT -108.230 -215.040 -106.025 -214.870 ;
        RECT -108.720 -217.390 -108.550 -215.530 ;
        RECT -108.230 -217.070 -108.060 -215.040 ;
        RECT -107.180 -215.055 -106.025 -215.040 ;
        RECT -107.740 -217.390 -107.570 -215.530 ;
        RECT -107.180 -215.585 -107.005 -215.055 ;
        RECT -107.175 -217.070 -107.005 -215.585 ;
        RECT -106.685 -217.070 -106.515 -215.530 ;
        RECT -106.200 -215.575 -106.025 -215.055 ;
        RECT -106.195 -217.070 -106.025 -215.575 ;
        RECT -106.690 -217.385 -106.515 -217.070 ;
        RECT -105.625 -217.385 -105.455 -215.535 ;
        RECT -105.135 -217.075 -104.965 -214.590 ;
        RECT -91.405 -215.460 -91.235 -214.420 ;
        RECT -90.425 -215.460 -90.255 -214.420 ;
        RECT -89.445 -215.460 -89.275 -214.420 ;
        RECT -86.540 -215.495 -86.370 -213.775 ;
        RECT -85.560 -215.495 -85.390 -213.775 ;
        RECT -83.495 -214.310 -83.325 -213.770 ;
        RECT -82.515 -214.310 -82.345 -213.770 ;
        RECT -84.085 -214.545 -83.720 -214.480 ;
        RECT -84.585 -214.685 -83.720 -214.545 ;
        RECT -84.695 -214.750 -83.720 -214.685 ;
        RECT -84.695 -215.495 -84.390 -214.750 ;
        RECT -84.085 -214.780 -83.720 -214.750 ;
        RECT -81.535 -214.630 -81.365 -213.770 ;
        RECT -80.025 -214.630 -79.675 -207.945 ;
        RECT -32.835 -208.520 -32.665 -207.560 ;
        RECT -31.855 -208.520 -31.685 -207.560 ;
        RECT -30.905 -208.500 -30.675 -207.235 ;
        RECT -28.670 -207.555 -27.795 -207.130 ;
        RECT -25.875 -207.285 -25.015 -206.915 ;
        RECT -28.670 -207.725 -25.530 -207.555 ;
        RECT -28.670 -207.945 -28.460 -207.725 ;
        RECT -28.645 -208.445 -28.475 -207.945 ;
        RECT -28.155 -208.360 -27.985 -207.905 ;
        RECT -27.670 -207.995 -27.490 -207.725 ;
        RECT -26.700 -207.905 -26.520 -207.725 ;
        RECT -30.875 -208.520 -30.705 -208.500 ;
        RECT -28.180 -208.615 -27.970 -208.360 ;
        RECT -27.665 -208.445 -27.495 -207.995 ;
        RECT -27.175 -208.335 -27.005 -207.905 ;
        RECT -26.700 -207.995 -26.515 -207.905 ;
        RECT -27.200 -208.615 -26.990 -208.335 ;
        RECT -26.685 -208.445 -26.515 -207.995 ;
        RECT -26.195 -208.340 -26.025 -207.905 ;
        RECT -25.710 -207.985 -25.530 -207.725 ;
        RECT -26.230 -208.615 -26.020 -208.340 ;
        RECT -25.705 -208.445 -25.535 -207.985 ;
        RECT -25.250 -208.020 -25.015 -207.285 ;
        RECT -24.790 -207.005 -23.920 -206.845 ;
        RECT -23.170 -207.005 -22.940 -206.540 ;
        RECT -22.650 -206.620 -22.480 -205.825 ;
        RECT -22.160 -206.540 -21.990 -206.080 ;
        RECT -22.190 -207.005 -21.960 -206.540 ;
        RECT -21.670 -206.620 -21.500 -205.825 ;
        RECT -20.065 -206.900 -19.765 -206.325 ;
        RECT -19.335 -206.540 -19.165 -206.080 ;
        RECT -19.365 -206.845 -19.135 -206.540 ;
        RECT -18.845 -206.620 -18.675 -205.825 ;
        RECT -18.355 -206.540 -18.185 -206.080 ;
        RECT -19.515 -206.900 -19.135 -206.845 ;
        RECT -24.790 -207.195 -21.960 -207.005 ;
        RECT -24.790 -207.315 -24.425 -207.195 ;
        RECT -25.215 -208.390 -25.045 -208.020 ;
        RECT -24.795 -208.155 -24.425 -207.315 ;
        RECT -24.150 -207.235 -21.960 -207.195 ;
        RECT -24.150 -207.560 -23.920 -207.235 ;
        RECT -23.170 -207.560 -22.940 -207.235 ;
        RECT -25.220 -208.615 -25.040 -208.390 ;
        RECT -24.120 -208.520 -23.950 -207.560 ;
        RECT -23.140 -208.520 -22.970 -207.560 ;
        RECT -22.190 -208.500 -21.960 -207.235 ;
        RECT -20.090 -207.005 -19.135 -206.900 ;
        RECT -18.385 -207.005 -18.155 -206.540 ;
        RECT -17.865 -206.620 -17.695 -205.825 ;
        RECT -17.375 -206.540 -17.205 -206.080 ;
        RECT -17.405 -207.005 -17.175 -206.540 ;
        RECT -16.885 -206.620 -16.715 -205.825 ;
        RECT -15.160 -206.300 -14.930 -205.690 ;
        RECT -14.685 -205.890 -14.465 -205.600 ;
        RECT -15.165 -206.350 -14.930 -206.300 ;
        RECT -15.165 -206.515 -14.960 -206.350 ;
        RECT -14.655 -206.370 -14.485 -205.890 ;
        RECT -14.165 -206.305 -13.995 -205.830 ;
        RECT -13.700 -205.945 -13.480 -205.600 ;
        RECT -15.170 -206.550 -14.960 -206.515 ;
        RECT -14.180 -206.550 -13.975 -206.305 ;
        RECT -13.675 -206.370 -13.505 -205.945 ;
        RECT -13.185 -206.305 -13.015 -205.830 ;
        RECT -12.720 -205.945 -12.500 -205.600 ;
        RECT -13.210 -206.550 -13.005 -206.305 ;
        RECT -12.695 -206.370 -12.525 -205.945 ;
        RECT -12.205 -206.345 -12.035 -205.830 ;
        RECT -11.740 -205.890 -11.520 -205.600 ;
        RECT -10.625 -205.825 -3.545 -205.485 ;
        RECT -11.715 -206.240 -11.545 -205.890 ;
        RECT -12.220 -206.550 -12.015 -206.345 ;
        RECT -15.170 -206.720 -12.015 -206.550 ;
        RECT -20.090 -207.125 -17.175 -207.005 ;
        RECT -21.170 -207.795 -20.885 -207.590 ;
        RECT -20.090 -207.795 -19.865 -207.125 ;
        RECT -19.515 -207.195 -17.175 -207.125 ;
        RECT -16.995 -206.830 -16.155 -206.790 ;
        RECT -15.170 -206.830 -14.295 -206.720 ;
        RECT -16.995 -207.115 -14.295 -206.830 ;
        RECT -11.750 -206.915 -11.515 -206.240 ;
        RECT -10.620 -206.540 -10.450 -206.080 ;
        RECT -10.650 -206.845 -10.420 -206.540 ;
        RECT -10.130 -206.620 -9.960 -205.825 ;
        RECT -9.640 -206.540 -9.470 -206.080 ;
        RECT -16.995 -207.160 -16.155 -207.115 ;
        RECT -19.365 -207.235 -17.175 -207.195 ;
        RECT -19.365 -207.560 -19.135 -207.235 ;
        RECT -18.385 -207.560 -18.155 -207.235 ;
        RECT -21.170 -208.020 -19.865 -207.795 ;
        RECT -21.170 -208.410 -20.885 -208.020 ;
        RECT -22.160 -208.520 -21.990 -208.500 ;
        RECT -19.335 -208.520 -19.165 -207.560 ;
        RECT -18.355 -208.520 -18.185 -207.560 ;
        RECT -17.405 -208.500 -17.175 -207.235 ;
        RECT -15.170 -207.555 -14.295 -207.115 ;
        RECT -12.375 -207.285 -11.515 -206.915 ;
        RECT -15.170 -207.725 -12.030 -207.555 ;
        RECT -15.170 -207.945 -14.960 -207.725 ;
        RECT -15.145 -208.445 -14.975 -207.945 ;
        RECT -14.655 -208.360 -14.485 -207.905 ;
        RECT -14.170 -207.995 -13.990 -207.725 ;
        RECT -13.200 -207.905 -13.020 -207.725 ;
        RECT -17.375 -208.520 -17.205 -208.500 ;
        RECT -28.180 -208.785 -25.040 -208.615 ;
        RECT -14.680 -208.615 -14.470 -208.360 ;
        RECT -14.165 -208.445 -13.995 -207.995 ;
        RECT -13.675 -208.335 -13.505 -207.905 ;
        RECT -13.200 -207.995 -13.015 -207.905 ;
        RECT -13.700 -208.615 -13.490 -208.335 ;
        RECT -13.185 -208.445 -13.015 -207.995 ;
        RECT -12.695 -208.340 -12.525 -207.905 ;
        RECT -12.210 -207.985 -12.030 -207.725 ;
        RECT -12.730 -208.615 -12.520 -208.340 ;
        RECT -12.205 -208.445 -12.035 -207.985 ;
        RECT -11.750 -208.020 -11.515 -207.285 ;
        RECT -11.290 -207.005 -10.420 -206.845 ;
        RECT -9.670 -207.005 -9.440 -206.540 ;
        RECT -9.150 -206.620 -8.980 -205.825 ;
        RECT -8.660 -206.540 -8.490 -206.080 ;
        RECT -8.690 -207.005 -8.460 -206.540 ;
        RECT -8.170 -206.620 -8.000 -205.825 ;
        RECT -11.290 -207.195 -8.460 -207.005 ;
        RECT -8.280 -206.815 -7.440 -206.790 ;
        RECT -8.280 -206.875 -7.265 -206.815 ;
        RECT -6.980 -206.875 -6.680 -206.445 ;
        RECT -6.210 -206.540 -6.040 -206.080 ;
        RECT -6.240 -206.845 -6.010 -206.540 ;
        RECT -5.720 -206.620 -5.550 -205.825 ;
        RECT -5.230 -206.540 -5.060 -206.080 ;
        RECT -6.390 -206.875 -6.010 -206.845 ;
        RECT -8.280 -207.005 -6.010 -206.875 ;
        RECT -5.260 -207.005 -5.030 -206.540 ;
        RECT -4.740 -206.620 -4.570 -205.825 ;
        RECT -4.250 -206.540 -4.080 -206.080 ;
        RECT -4.280 -207.005 -4.050 -206.540 ;
        RECT -3.760 -206.620 -3.590 -205.825 ;
        RECT -1.560 -206.120 -1.390 -203.855 ;
        RECT -1.070 -204.895 -0.900 -202.915 ;
        RECT 0.995 -203.365 3.200 -203.195 ;
        RECT 0.505 -205.715 0.675 -203.855 ;
        RECT 0.995 -205.395 1.165 -203.365 ;
        RECT 2.045 -203.380 3.200 -203.365 ;
        RECT 1.485 -205.715 1.655 -203.855 ;
        RECT 2.045 -203.910 2.220 -203.380 ;
        RECT 2.050 -205.395 2.220 -203.910 ;
        RECT 2.540 -205.395 2.710 -203.855 ;
        RECT 3.025 -203.900 3.200 -203.380 ;
        RECT 3.030 -205.395 3.200 -203.900 ;
        RECT 2.535 -205.710 2.710 -205.395 ;
        RECT 3.600 -205.710 3.770 -203.860 ;
        RECT 4.090 -205.400 4.260 -202.915 ;
        RECT 8.410 -203.665 9.165 -201.265 ;
        RECT 10.295 -203.575 10.915 -201.265 ;
        RECT 11.945 -203.575 12.565 -201.265 ;
        RECT 13.980 -203.475 14.660 -203.245 ;
        RECT 10.295 -203.665 12.870 -203.575 ;
        RECT 2.535 -205.715 3.770 -205.710 ;
        RECT 4.580 -205.715 4.750 -203.860 ;
        RECT 0.505 -205.885 1.670 -205.715 ;
        RECT 2.535 -205.885 4.750 -205.715 ;
        RECT 8.410 -203.880 12.870 -203.665 ;
        RECT 8.410 -203.970 10.660 -203.880 ;
        RECT -2.315 -206.385 -1.390 -206.120 ;
        RECT -8.280 -207.085 -4.050 -207.005 ;
        RECT -8.280 -207.105 -7.265 -207.085 ;
        RECT -6.980 -207.105 -6.680 -207.085 ;
        RECT -8.280 -207.160 -7.440 -207.105 ;
        RECT -6.390 -207.195 -4.050 -207.085 ;
        RECT -11.290 -207.315 -10.925 -207.195 ;
        RECT -11.715 -208.390 -11.545 -208.020 ;
        RECT -11.295 -208.155 -10.925 -207.315 ;
        RECT -10.650 -207.235 -8.460 -207.195 ;
        RECT -10.650 -207.560 -10.420 -207.235 ;
        RECT -9.670 -207.560 -9.440 -207.235 ;
        RECT -11.720 -208.615 -11.540 -208.390 ;
        RECT -10.620 -208.520 -10.450 -207.560 ;
        RECT -9.640 -208.520 -9.470 -207.560 ;
        RECT -8.690 -208.500 -8.460 -207.235 ;
        RECT -6.240 -207.235 -4.050 -207.195 ;
        RECT -6.240 -207.560 -6.010 -207.235 ;
        RECT -5.260 -207.560 -5.030 -207.235 ;
        RECT -7.670 -208.410 -7.385 -207.590 ;
        RECT -8.660 -208.520 -8.490 -208.500 ;
        RECT -6.210 -208.520 -6.040 -207.560 ;
        RECT -5.230 -208.520 -5.060 -207.560 ;
        RECT -4.280 -208.500 -4.050 -207.235 ;
        RECT -1.560 -208.435 -1.390 -206.385 ;
        RECT -1.215 -206.155 -0.540 -206.120 ;
        RECT 1.485 -206.155 1.670 -205.885 ;
        RECT 8.410 -206.005 8.715 -203.970 ;
        RECT 12.110 -204.140 12.285 -203.880 ;
        RECT 10.640 -205.680 10.810 -204.140 ;
        RECT 11.130 -205.680 11.300 -204.140 ;
        RECT 11.620 -205.680 11.790 -204.140 ;
        RECT 12.110 -205.680 12.280 -204.140 ;
        RECT 12.600 -205.680 12.770 -204.140 ;
        RECT 10.500 -205.895 10.870 -205.865 ;
        RECT 12.575 -205.895 12.930 -205.890 ;
        RECT 10.500 -205.900 12.930 -205.895 ;
        RECT -1.215 -206.340 1.670 -206.155 ;
        RECT -1.215 -206.390 -0.540 -206.340 ;
        RECT 1.485 -207.030 1.670 -206.340 ;
        RECT 1.840 -206.165 2.515 -206.130 ;
        RECT 1.840 -206.335 6.620 -206.165 ;
        RECT 1.840 -206.400 2.515 -206.335 ;
        RECT 2.780 -206.555 3.455 -206.520 ;
        RECT 5.595 -206.555 6.275 -206.520 ;
        RECT 2.780 -206.745 6.275 -206.555 ;
        RECT 2.780 -206.790 3.455 -206.745 ;
        RECT 5.595 -206.750 6.275 -206.745 ;
        RECT 1.485 -207.215 4.260 -207.030 ;
        RECT 4.460 -207.200 5.420 -206.930 ;
        RECT 6.450 -207.160 6.620 -206.335 ;
        RECT 6.860 -206.435 9.935 -206.005 ;
        RECT 10.500 -206.090 13.835 -205.900 ;
        RECT 10.500 -206.220 10.870 -206.090 ;
        RECT 12.925 -206.100 13.835 -206.090 ;
        RECT 12.520 -206.370 13.195 -206.340 ;
        RECT 12.520 -206.390 13.345 -206.370 ;
        RECT 2.130 -208.435 2.300 -207.215 ;
        RECT 3.110 -208.435 3.280 -207.215 ;
        RECT 4.090 -208.435 4.260 -207.215 ;
        RECT 5.190 -207.620 5.420 -207.200 ;
        RECT 6.420 -207.510 7.275 -207.160 ;
        RECT 7.595 -207.215 7.765 -206.675 ;
        RECT 8.085 -207.215 8.255 -206.435 ;
        RECT 8.575 -207.215 8.745 -206.675 ;
        RECT 9.065 -207.215 9.235 -206.435 ;
        RECT 10.185 -206.495 12.280 -206.455 ;
        RECT 10.130 -206.645 12.280 -206.495 ;
        RECT 12.520 -206.570 13.455 -206.390 ;
        RECT 12.520 -206.610 13.410 -206.570 ;
        RECT 7.105 -208.370 7.275 -207.510 ;
        RECT 9.460 -207.390 9.825 -207.360 ;
        RECT 10.130 -207.390 10.435 -206.645 ;
        RECT 9.460 -207.455 10.435 -207.390 ;
        RECT 9.460 -207.595 10.325 -207.455 ;
        RECT 9.460 -207.660 9.825 -207.595 ;
        RECT 8.085 -208.370 8.255 -207.830 ;
        RECT 9.065 -208.370 9.235 -207.830 ;
        RECT 11.130 -208.365 11.300 -206.645 ;
        RECT 12.110 -208.365 12.280 -206.645 ;
        RECT -4.250 -208.520 -4.080 -208.500 ;
        RECT -14.680 -208.785 -11.540 -208.615 ;
        RECT 13.230 -210.360 13.410 -206.610 ;
        RECT -34.490 -210.635 -33.810 -210.405 ;
        RECT 12.635 -210.590 13.410 -210.360 ;
        RECT -106.690 -217.390 -105.455 -217.385 ;
        RECT -104.645 -217.390 -104.475 -215.535 ;
        RECT -87.455 -215.560 -86.780 -215.530 ;
        RECT -87.555 -215.570 -86.780 -215.560 ;
        RECT -92.865 -215.695 -92.215 -215.610 ;
        RECT -91.995 -215.695 -91.630 -215.630 ;
        RECT -95.540 -215.725 -95.250 -215.720 ;
        RECT -92.865 -215.725 -91.630 -215.695 ;
        RECT -95.540 -215.900 -91.630 -215.725 ;
        RECT -88.590 -215.750 -86.780 -215.570 ;
        RECT -86.540 -215.645 -84.390 -215.495 ;
        RECT -86.540 -215.685 -84.445 -215.645 ;
        RECT -83.495 -215.705 -83.325 -214.925 ;
        RECT -83.005 -215.465 -82.835 -214.925 ;
        RECT -82.515 -215.705 -82.345 -214.925 ;
        RECT -82.025 -215.465 -81.855 -214.925 ;
        RECT -81.535 -214.980 -79.675 -214.630 ;
        RECT -87.555 -215.760 -86.780 -215.750 ;
        RECT -87.455 -215.800 -86.780 -215.760 ;
        RECT -95.540 -216.065 -92.215 -215.900 ;
        RECT -91.995 -215.930 -91.630 -215.900 ;
        RECT -95.540 -216.405 -95.250 -216.065 ;
        RECT -92.865 -216.360 -92.215 -216.065 ;
        RECT -89.930 -216.050 -87.185 -216.040 ;
        RECT -85.130 -216.050 -84.760 -215.920 ;
        RECT -89.930 -216.070 -84.760 -216.050 ;
        RECT -108.720 -217.560 -107.555 -217.390 ;
        RECT -106.690 -217.560 -104.475 -217.390 ;
        RECT -110.440 -217.830 -109.765 -217.795 ;
        RECT -107.740 -217.830 -107.555 -217.560 ;
        RECT -110.440 -218.015 -107.555 -217.830 ;
        RECT -110.440 -218.065 -109.765 -218.015 ;
        RECT -107.740 -218.705 -107.555 -218.015 ;
        RECT -107.385 -217.840 -106.710 -217.805 ;
        RECT -104.240 -217.840 -103.950 -217.325 ;
        RECT -91.405 -217.350 -91.235 -216.070 ;
        RECT -90.915 -217.110 -90.745 -216.070 ;
        RECT -90.425 -217.350 -90.255 -216.070 ;
        RECT -89.935 -216.240 -84.760 -216.070 ;
        RECT -84.195 -216.135 -80.270 -215.705 ;
        RECT -89.935 -217.110 -89.765 -216.240 ;
        RECT -87.190 -216.245 -84.760 -216.240 ;
        RECT -87.190 -216.250 -86.835 -216.245 ;
        RECT -85.130 -216.275 -84.760 -216.245 ;
        RECT -107.385 -218.010 -103.950 -217.840 ;
        RECT -107.385 -218.075 -106.710 -218.010 ;
        RECT -106.445 -218.230 -105.770 -218.195 ;
        RECT -100.590 -218.230 -100.300 -217.735 ;
        RECT -92.105 -217.780 -87.415 -217.350 ;
        RECT -106.445 -218.420 -100.300 -218.230 ;
        RECT -106.445 -218.465 -105.770 -218.420 ;
        RECT -104.765 -218.650 -104.090 -218.605 ;
        RECT -95.965 -218.650 -95.675 -218.165 ;
        RECT -87.845 -218.185 -87.415 -217.780 ;
        RECT -87.030 -218.000 -86.860 -216.460 ;
        RECT -86.540 -218.000 -86.370 -216.460 ;
        RECT -86.050 -218.000 -85.880 -216.460 ;
        RECT -85.560 -218.000 -85.390 -216.460 ;
        RECT -85.070 -218.000 -84.900 -216.460 ;
        RECT -86.545 -218.185 -86.370 -218.000 ;
        RECT -82.975 -218.170 -82.670 -216.135 ;
        RECT -84.920 -218.185 -82.670 -218.170 ;
        RECT -87.845 -218.475 -82.670 -218.185 ;
        RECT -34.290 -218.290 -34.120 -210.635 ;
        RECT -22.090 -211.000 -21.410 -210.770 ;
        RECT 13.635 -210.780 13.835 -206.100 ;
        RECT 14.310 -207.150 14.660 -203.475 ;
        RECT 16.435 -203.655 17.190 -201.265 ;
        RECT 18.645 -203.565 19.400 -201.265 ;
        RECT 20.110 -203.565 20.865 -201.265 ;
        RECT 23.310 -202.635 24.040 -201.265 ;
        RECT 25.535 -202.635 26.265 -201.265 ;
        RECT 26.865 -202.635 27.595 -201.265 ;
        RECT 28.665 -202.635 29.395 -201.265 ;
        RECT 21.820 -202.915 22.500 -202.685 ;
        RECT 18.645 -203.655 20.895 -203.565 ;
        RECT 16.435 -203.870 20.895 -203.655 ;
        RECT 16.435 -203.960 18.685 -203.870 ;
        RECT 16.435 -205.995 16.740 -203.960 ;
        RECT 20.135 -204.130 20.310 -203.870 ;
        RECT 18.665 -205.670 18.835 -204.130 ;
        RECT 19.155 -205.670 19.325 -204.130 ;
        RECT 19.645 -205.670 19.815 -204.130 ;
        RECT 20.135 -205.670 20.305 -204.130 ;
        RECT 20.625 -205.670 20.795 -204.130 ;
        RECT 22.170 -205.190 22.495 -202.915 ;
        RECT 23.190 -202.960 29.560 -202.635 ;
        RECT 23.250 -205.190 23.420 -203.900 ;
        RECT 23.740 -204.940 23.910 -202.960 ;
        RECT 25.805 -203.410 28.010 -203.240 ;
        RECT 22.170 -205.480 23.420 -205.190 ;
        RECT 18.525 -205.885 18.895 -205.855 ;
        RECT 20.600 -205.885 20.955 -205.880 ;
        RECT 18.525 -205.890 20.955 -205.885 ;
        RECT 14.885 -206.425 17.960 -205.995 ;
        RECT 18.525 -206.080 21.975 -205.890 ;
        RECT 18.525 -206.210 18.895 -206.080 ;
        RECT 20.950 -206.090 21.975 -206.080 ;
        RECT 20.545 -206.370 21.220 -206.330 ;
        RECT 20.545 -206.380 21.480 -206.370 ;
        RECT 14.310 -207.500 15.300 -207.150 ;
        RECT 15.620 -207.205 15.790 -206.665 ;
        RECT 16.110 -207.205 16.280 -206.425 ;
        RECT 16.600 -207.205 16.770 -206.665 ;
        RECT 17.090 -207.205 17.260 -206.425 ;
        RECT 18.210 -206.485 20.305 -206.445 ;
        RECT 18.155 -206.635 20.305 -206.485 ;
        RECT 20.545 -206.570 21.580 -206.380 ;
        RECT 20.545 -206.600 21.220 -206.570 ;
        RECT 15.130 -208.360 15.300 -207.500 ;
        RECT 17.485 -207.380 17.850 -207.350 ;
        RECT 18.155 -207.380 18.460 -206.635 ;
        RECT 17.485 -207.445 18.460 -207.380 ;
        RECT 17.485 -207.585 18.350 -207.445 ;
        RECT 17.485 -207.650 17.850 -207.585 ;
        RECT 16.110 -208.360 16.280 -207.820 ;
        RECT 17.090 -208.360 17.260 -207.820 ;
        RECT 19.155 -208.355 19.325 -206.635 ;
        RECT 20.135 -208.355 20.305 -206.635 ;
        RECT -22.090 -212.265 -21.890 -211.000 ;
        RECT 13.155 -211.010 13.835 -210.780 ;
        RECT -22.105 -212.945 -21.875 -212.265 ;
        RECT 21.400 -213.205 21.580 -206.570 ;
        RECT 13.975 -213.385 21.580 -213.205 ;
        RECT 13.975 -213.945 14.155 -213.385 ;
        RECT 21.775 -213.555 21.975 -206.090 ;
        RECT 23.250 -208.480 23.420 -205.480 ;
        RECT 25.315 -205.760 25.485 -203.900 ;
        RECT 25.805 -205.440 25.975 -203.410 ;
        RECT 26.855 -203.425 28.010 -203.410 ;
        RECT 26.295 -205.760 26.465 -203.900 ;
        RECT 26.855 -203.955 27.030 -203.425 ;
        RECT 26.860 -205.440 27.030 -203.955 ;
        RECT 27.350 -205.440 27.520 -203.900 ;
        RECT 27.835 -203.945 28.010 -203.425 ;
        RECT 27.840 -205.440 28.010 -203.945 ;
        RECT 27.345 -205.755 27.520 -205.440 ;
        RECT 28.410 -205.755 28.580 -203.905 ;
        RECT 28.900 -205.445 29.070 -202.960 ;
        RECT 31.485 -203.535 32.470 -201.265 ;
        RECT 34.150 -203.535 35.135 -201.265 ;
        RECT 36.715 -203.490 37.700 -201.265 ;
        RECT 39.230 -203.490 40.215 -201.265 ;
        RECT 41.205 -203.400 42.510 -201.265 ;
        RECT 48.930 -200.950 49.250 -200.835 ;
        RECT 75.755 -200.950 76.170 -199.975 ;
        RECT 80.040 -200.085 81.145 -199.975 ;
        RECT 48.930 -201.365 76.170 -200.950 ;
        RECT 48.930 -201.425 49.250 -201.365 ;
        RECT 95.455 -201.755 96.200 -189.080 ;
        RECT 98.260 -191.730 99.180 -189.080 ;
        RECT 101.380 -189.250 101.590 -189.030 ;
        RECT 101.895 -189.070 102.065 -188.615 ;
        RECT 102.385 -188.980 102.555 -188.530 ;
        RECT 102.850 -188.640 103.060 -188.360 ;
        RECT 102.380 -189.250 102.560 -188.980 ;
        RECT 102.875 -189.070 103.045 -188.640 ;
        RECT 103.365 -188.980 103.535 -188.530 ;
        RECT 103.820 -188.635 104.030 -188.360 ;
        RECT 103.350 -189.070 103.535 -188.980 ;
        RECT 103.855 -189.070 104.025 -188.635 ;
        RECT 104.345 -188.990 104.515 -188.530 ;
        RECT 104.830 -188.585 105.010 -188.360 ;
        RECT 115.370 -188.360 118.510 -188.190 ;
        RECT 104.835 -188.955 105.005 -188.585 ;
        RECT 103.350 -189.250 103.530 -189.070 ;
        RECT 104.340 -189.250 104.520 -188.990 ;
        RECT 101.380 -189.420 104.520 -189.250 ;
        RECT 101.380 -189.965 102.255 -189.420 ;
        RECT 104.800 -189.690 105.035 -188.955 ;
        RECT 105.255 -189.660 105.625 -188.820 ;
        RECT 105.930 -189.415 106.100 -188.455 ;
        RECT 106.910 -189.415 107.080 -188.455 ;
        RECT 107.890 -188.475 108.060 -188.455 ;
        RECT 101.005 -190.255 102.255 -189.965 ;
        RECT 104.175 -190.060 105.035 -189.690 ;
        RECT 101.005 -190.265 104.535 -190.255 ;
        RECT 101.380 -190.425 104.535 -190.265 ;
        RECT 101.380 -190.460 101.590 -190.425 ;
        RECT 101.385 -190.675 101.590 -190.460 ;
        RECT 101.405 -191.145 101.575 -190.675 ;
        RECT 101.895 -191.085 102.065 -190.605 ;
        RECT 102.370 -190.670 102.575 -190.425 ;
        RECT 101.865 -191.375 102.085 -191.085 ;
        RECT 102.385 -191.145 102.555 -190.670 ;
        RECT 102.875 -191.030 103.045 -190.605 ;
        RECT 103.340 -190.670 103.545 -190.425 ;
        RECT 102.850 -191.375 103.070 -191.030 ;
        RECT 103.365 -191.145 103.535 -190.670 ;
        RECT 103.855 -191.030 104.025 -190.605 ;
        RECT 104.330 -190.630 104.535 -190.425 ;
        RECT 103.830 -191.375 104.050 -191.030 ;
        RECT 104.345 -191.145 104.515 -190.630 ;
        RECT 104.800 -190.735 105.035 -190.060 ;
        RECT 105.260 -189.780 105.625 -189.660 ;
        RECT 105.900 -189.740 106.130 -189.415 ;
        RECT 106.880 -189.740 107.110 -189.415 ;
        RECT 107.860 -189.740 108.090 -188.475 ;
        RECT 108.880 -188.825 109.165 -188.565 ;
        RECT 108.880 -189.135 109.905 -188.825 ;
        RECT 108.880 -189.385 109.165 -189.135 ;
        RECT 105.900 -189.780 108.090 -189.740 ;
        RECT 105.260 -189.970 108.090 -189.780 ;
        RECT 105.260 -190.130 106.130 -189.970 ;
        RECT 105.900 -190.435 106.130 -190.130 ;
        RECT 104.835 -191.085 105.005 -190.735 ;
        RECT 105.930 -190.895 106.100 -190.435 ;
        RECT 104.810 -191.375 105.030 -191.085 ;
        RECT 106.420 -191.150 106.590 -190.355 ;
        RECT 106.880 -190.435 107.110 -189.970 ;
        RECT 106.910 -190.895 107.080 -190.435 ;
        RECT 107.400 -191.150 107.570 -190.355 ;
        RECT 107.860 -190.435 108.090 -189.970 ;
        RECT 109.595 -189.780 109.905 -189.135 ;
        RECT 110.115 -189.415 110.285 -188.455 ;
        RECT 111.095 -189.415 111.265 -188.455 ;
        RECT 112.075 -188.475 112.245 -188.455 ;
        RECT 110.085 -189.740 110.315 -189.415 ;
        RECT 111.065 -189.740 111.295 -189.415 ;
        RECT 112.045 -189.740 112.275 -188.475 ;
        RECT 114.905 -189.030 115.075 -188.530 ;
        RECT 115.370 -188.615 115.580 -188.360 ;
        RECT 110.085 -189.780 112.275 -189.740 ;
        RECT 109.595 -189.970 112.275 -189.780 ;
        RECT 114.880 -189.250 115.090 -189.030 ;
        RECT 115.395 -189.070 115.565 -188.615 ;
        RECT 115.885 -188.980 116.055 -188.530 ;
        RECT 116.350 -188.640 116.560 -188.360 ;
        RECT 115.880 -189.250 116.060 -188.980 ;
        RECT 116.375 -189.070 116.545 -188.640 ;
        RECT 116.865 -188.980 117.035 -188.530 ;
        RECT 117.320 -188.635 117.530 -188.360 ;
        RECT 116.850 -189.070 117.035 -188.980 ;
        RECT 117.355 -189.070 117.525 -188.635 ;
        RECT 117.845 -188.990 118.015 -188.530 ;
        RECT 118.330 -188.585 118.510 -188.360 ;
        RECT 143.635 -188.375 143.805 -186.655 ;
        RECT 144.615 -188.375 144.785 -186.655 ;
        RECT 145.480 -187.400 145.785 -186.655 ;
        RECT 146.680 -187.225 146.850 -186.445 ;
        RECT 147.170 -187.225 147.340 -186.685 ;
        RECT 147.660 -187.225 147.830 -186.445 ;
        RECT 179.510 -186.510 180.745 -186.305 ;
        RECT 184.920 -186.445 185.595 -186.405 ;
        RECT 184.820 -186.455 185.595 -186.445 ;
        RECT 179.510 -186.595 180.160 -186.510 ;
        RECT 180.380 -186.575 180.745 -186.510 ;
        RECT 183.785 -186.635 185.595 -186.455 ;
        RECT 188.180 -186.500 192.105 -186.070 ;
        RECT 223.825 -186.500 224.475 -186.040 ;
        RECT 225.285 -186.330 225.455 -185.050 ;
        RECT 225.775 -186.330 225.945 -185.290 ;
        RECT 226.265 -186.330 226.435 -185.050 ;
        RECT 226.755 -186.160 226.925 -185.290 ;
        RECT 229.660 -185.940 229.830 -184.400 ;
        RECT 230.150 -185.940 230.320 -184.400 ;
        RECT 230.640 -185.940 230.810 -184.400 ;
        RECT 231.130 -185.940 231.300 -184.400 ;
        RECT 231.620 -185.940 231.790 -184.400 ;
        RECT 229.500 -186.155 229.855 -186.150 ;
        RECT 231.560 -186.155 231.930 -186.125 ;
        RECT 229.500 -186.160 231.930 -186.155 ;
        RECT 226.755 -186.330 231.930 -186.160 ;
        RECT 233.715 -186.265 234.020 -184.230 ;
        RECT 257.490 -184.070 258.620 -184.025 ;
        RECT 265.755 -184.070 266.985 -183.670 ;
        RECT 257.490 -184.735 266.985 -184.070 ;
        RECT 274.835 -183.755 278.160 -183.615 ;
        RECT 274.835 -184.045 280.010 -183.755 ;
        RECT 274.835 -184.450 275.265 -184.045 ;
        RECT 276.135 -184.230 276.310 -184.045 ;
        RECT 277.760 -184.060 280.010 -184.045 ;
        RECT 257.490 -185.195 258.620 -184.735 ;
        RECT 265.755 -184.770 266.985 -184.735 ;
        RECT 270.575 -184.880 275.265 -184.450 ;
        RECT 226.760 -186.350 231.930 -186.330 ;
        RECT 226.760 -186.360 229.505 -186.350 ;
        RECT 224.695 -186.500 225.060 -186.470 ;
        RECT 231.560 -186.480 231.930 -186.350 ;
        RECT 184.820 -186.645 185.595 -186.635 ;
        RECT 184.920 -186.675 185.595 -186.645 ;
        RECT 185.835 -186.560 187.930 -186.520 ;
        RECT 148.150 -187.225 148.320 -186.685 ;
        RECT 185.835 -186.710 187.985 -186.560 ;
        RECT 146.090 -187.400 146.455 -187.370 ;
        RECT 145.480 -187.465 146.455 -187.400 ;
        RECT 145.590 -187.605 146.455 -187.465 ;
        RECT 146.090 -187.670 146.455 -187.605 ;
        RECT 148.640 -187.520 150.500 -187.170 ;
        RECT 146.680 -188.380 146.850 -187.840 ;
        RECT 147.660 -188.380 147.830 -187.840 ;
        RECT 148.640 -188.380 148.810 -187.520 ;
        RECT 118.335 -188.955 118.505 -188.585 ;
        RECT 116.850 -189.250 117.030 -189.070 ;
        RECT 117.840 -189.250 118.020 -188.990 ;
        RECT 114.880 -189.420 118.020 -189.250 ;
        RECT 109.595 -190.130 110.315 -189.970 ;
        RECT 107.890 -190.895 108.060 -190.435 ;
        RECT 108.380 -191.150 108.550 -190.355 ;
        RECT 110.085 -190.435 110.315 -190.130 ;
        RECT 110.115 -190.895 110.285 -190.435 ;
        RECT 110.605 -191.150 110.775 -190.355 ;
        RECT 111.065 -190.435 111.295 -189.970 ;
        RECT 111.095 -190.895 111.265 -190.435 ;
        RECT 111.585 -191.150 111.755 -190.355 ;
        RECT 112.045 -190.435 112.275 -189.970 ;
        RECT 112.455 -189.850 113.295 -189.815 ;
        RECT 112.455 -190.150 113.405 -189.850 ;
        RECT 114.880 -189.955 115.755 -189.420 ;
        RECT 118.300 -189.690 118.535 -188.955 ;
        RECT 118.755 -189.660 119.125 -188.820 ;
        RECT 119.430 -189.415 119.600 -188.455 ;
        RECT 120.410 -189.415 120.580 -188.455 ;
        RECT 121.390 -188.475 121.560 -188.455 ;
        RECT 112.455 -190.185 113.295 -190.150 ;
        RECT 114.425 -190.255 115.755 -189.955 ;
        RECT 117.675 -190.060 118.535 -189.690 ;
        RECT 112.075 -190.895 112.245 -190.435 ;
        RECT 112.565 -191.150 112.735 -190.355 ;
        RECT 114.880 -190.425 118.035 -190.255 ;
        RECT 114.880 -190.460 115.090 -190.425 ;
        RECT 114.885 -190.675 115.090 -190.460 ;
        RECT 114.905 -191.145 115.075 -190.675 ;
        RECT 115.395 -191.085 115.565 -190.605 ;
        RECT 115.870 -190.670 116.075 -190.425 ;
        RECT 101.865 -191.545 105.030 -191.375 ;
        RECT 105.925 -191.160 108.595 -191.150 ;
        RECT 110.110 -191.160 112.780 -191.150 ;
        RECT 105.925 -191.490 112.780 -191.160 ;
        RECT 115.365 -191.375 115.585 -191.085 ;
        RECT 115.885 -191.145 116.055 -190.670 ;
        RECT 116.375 -191.030 116.545 -190.605 ;
        RECT 116.840 -190.670 117.045 -190.425 ;
        RECT 116.350 -191.375 116.570 -191.030 ;
        RECT 116.865 -191.145 117.035 -190.670 ;
        RECT 117.355 -191.030 117.525 -190.605 ;
        RECT 117.830 -190.630 118.035 -190.425 ;
        RECT 117.330 -191.375 117.550 -191.030 ;
        RECT 117.845 -191.145 118.015 -190.630 ;
        RECT 118.300 -190.735 118.535 -190.060 ;
        RECT 118.760 -189.780 119.125 -189.660 ;
        RECT 119.400 -189.740 119.630 -189.415 ;
        RECT 120.380 -189.740 120.610 -189.415 ;
        RECT 121.360 -189.740 121.590 -188.475 ;
        RECT 122.380 -188.885 122.665 -188.565 ;
        RECT 122.380 -189.130 123.380 -188.885 ;
        RECT 122.380 -189.385 122.665 -189.130 ;
        RECT 119.400 -189.780 121.590 -189.740 ;
        RECT 118.760 -189.970 121.590 -189.780 ;
        RECT 123.150 -189.780 123.380 -189.130 ;
        RECT 123.615 -189.415 123.785 -188.455 ;
        RECT 124.595 -189.415 124.765 -188.455 ;
        RECT 125.575 -188.475 125.745 -188.455 ;
        RECT 123.585 -189.740 123.815 -189.415 ;
        RECT 124.565 -189.740 124.795 -189.415 ;
        RECT 125.545 -189.740 125.775 -188.475 ;
        RECT 123.585 -189.780 125.775 -189.740 ;
        RECT 118.760 -190.130 119.630 -189.970 ;
        RECT 119.400 -190.435 119.630 -190.130 ;
        RECT 118.335 -191.085 118.505 -190.735 ;
        RECT 119.430 -190.895 119.600 -190.435 ;
        RECT 118.310 -191.375 118.530 -191.085 ;
        RECT 119.920 -191.150 120.090 -190.355 ;
        RECT 120.380 -190.435 120.610 -189.970 ;
        RECT 120.410 -190.895 120.580 -190.435 ;
        RECT 120.900 -191.150 121.070 -190.355 ;
        RECT 121.360 -190.435 121.590 -189.970 ;
        RECT 121.770 -189.870 122.610 -189.815 ;
        RECT 121.770 -189.875 122.785 -189.870 ;
        RECT 121.770 -190.185 122.970 -189.875 ;
        RECT 123.150 -189.970 125.775 -189.780 ;
        RECT 123.150 -190.130 123.815 -189.970 ;
        RECT 121.390 -190.895 121.560 -190.435 ;
        RECT 121.880 -191.150 122.050 -190.355 ;
        RECT 122.670 -190.905 122.970 -190.185 ;
        RECT 123.585 -190.435 123.815 -190.130 ;
        RECT 123.615 -190.895 123.785 -190.435 ;
        RECT 124.105 -191.150 124.275 -190.355 ;
        RECT 124.565 -190.435 124.795 -189.970 ;
        RECT 124.595 -190.895 124.765 -190.435 ;
        RECT 125.085 -191.150 125.255 -190.355 ;
        RECT 125.545 -190.435 125.775 -189.970 ;
        RECT 125.955 -189.965 126.795 -189.815 ;
        RECT 125.955 -190.185 126.830 -189.965 ;
        RECT 125.575 -190.895 125.745 -190.435 ;
        RECT 126.065 -191.150 126.235 -190.355 ;
        RECT 107.050 -191.730 107.605 -191.490 ;
        RECT 108.480 -191.500 111.080 -191.490 ;
        RECT 111.440 -191.720 111.995 -191.490 ;
        RECT 115.365 -191.545 118.530 -191.375 ;
        RECT 119.425 -191.490 126.280 -191.150 ;
        RECT 111.425 -191.730 112.110 -191.720 ;
        RECT 120.430 -191.730 120.985 -191.490 ;
        RECT 124.485 -191.690 125.040 -191.490 ;
        RECT 124.410 -191.730 125.095 -191.690 ;
        RECT 98.255 -191.925 125.180 -191.730 ;
        RECT 98.260 -192.020 98.920 -191.925 ;
        RECT 111.425 -192.020 112.110 -191.925 ;
        RECT 124.410 -191.990 125.095 -191.925 ;
        RECT 126.590 -192.045 126.830 -190.185 ;
        RECT 146.910 -190.720 148.110 -190.550 ;
        RECT 99.875 -192.620 100.535 -192.570 ;
        RECT 122.490 -192.620 123.150 -192.580 ;
        RECT 99.875 -192.815 125.180 -192.620 ;
        RECT 126.535 -192.730 126.835 -192.045 ;
        RECT 99.875 -192.870 100.535 -192.815 ;
        RECT 122.490 -192.880 123.150 -192.815 ;
        RECT 96.945 -193.390 104.025 -193.050 ;
        RECT 104.920 -193.165 108.085 -192.995 ;
        RECT 96.990 -194.185 97.160 -193.390 ;
        RECT 97.480 -194.105 97.650 -193.645 ;
        RECT 97.450 -194.570 97.680 -194.105 ;
        RECT 97.970 -194.185 98.140 -193.390 ;
        RECT 98.460 -194.105 98.630 -193.645 ;
        RECT 98.430 -194.570 98.660 -194.105 ;
        RECT 98.950 -194.185 99.120 -193.390 ;
        RECT 99.440 -194.105 99.610 -193.645 ;
        RECT 99.410 -194.410 99.640 -194.105 ;
        RECT 99.410 -194.440 99.790 -194.410 ;
        RECT 100.080 -194.440 100.380 -194.010 ;
        RECT 101.400 -194.185 101.570 -193.390 ;
        RECT 101.890 -194.105 102.060 -193.645 ;
        RECT 100.840 -194.380 101.680 -194.355 ;
        RECT 100.665 -194.440 101.680 -194.380 ;
        RECT 99.410 -194.570 101.680 -194.440 ;
        RECT 97.450 -194.650 101.680 -194.570 ;
        RECT 97.450 -194.760 99.790 -194.650 ;
        RECT 100.080 -194.670 100.380 -194.650 ;
        RECT 100.665 -194.670 101.680 -194.650 ;
        RECT 100.840 -194.725 101.680 -194.670 ;
        RECT 101.860 -194.570 102.090 -194.105 ;
        RECT 102.380 -194.185 102.550 -193.390 ;
        RECT 102.870 -194.105 103.040 -193.645 ;
        RECT 102.840 -194.570 103.070 -194.105 ;
        RECT 103.360 -194.185 103.530 -193.390 ;
        RECT 104.920 -193.455 105.140 -193.165 ;
        RECT 103.850 -194.105 104.020 -193.645 ;
        RECT 104.945 -193.805 105.115 -193.455 ;
        RECT 103.820 -194.410 104.050 -194.105 ;
        RECT 103.820 -194.570 104.690 -194.410 ;
        RECT 101.860 -194.760 104.690 -194.570 ;
        RECT 97.450 -194.800 99.640 -194.760 ;
        RECT 97.450 -196.065 97.680 -194.800 ;
        RECT 98.430 -195.125 98.660 -194.800 ;
        RECT 99.410 -195.125 99.640 -194.800 ;
        RECT 101.860 -194.800 104.050 -194.760 ;
        RECT 97.480 -196.085 97.650 -196.065 ;
        RECT 98.460 -196.085 98.630 -195.125 ;
        RECT 99.440 -196.085 99.610 -195.125 ;
        RECT 100.785 -195.975 101.070 -195.155 ;
        RECT 101.860 -196.065 102.090 -194.800 ;
        RECT 102.840 -195.125 103.070 -194.800 ;
        RECT 103.820 -195.125 104.050 -194.800 ;
        RECT 104.325 -194.880 104.690 -194.760 ;
        RECT 104.915 -194.480 105.150 -193.805 ;
        RECT 105.435 -193.910 105.605 -193.395 ;
        RECT 105.900 -193.510 106.120 -193.165 ;
        RECT 105.415 -194.115 105.620 -193.910 ;
        RECT 105.925 -193.935 106.095 -193.510 ;
        RECT 106.415 -193.870 106.585 -193.395 ;
        RECT 106.880 -193.510 107.100 -193.165 ;
        RECT 106.405 -194.115 106.610 -193.870 ;
        RECT 106.905 -193.935 107.075 -193.510 ;
        RECT 107.395 -193.870 107.565 -193.395 ;
        RECT 107.865 -193.455 108.085 -193.165 ;
        RECT 107.375 -194.115 107.580 -193.870 ;
        RECT 107.885 -193.935 108.055 -193.455 ;
        RECT 108.330 -193.865 108.560 -193.255 ;
        RECT 110.070 -193.390 117.525 -193.050 ;
        RECT 118.420 -193.165 121.585 -192.995 ;
        RECT 108.330 -193.915 108.565 -193.865 ;
        RECT 108.360 -194.080 108.565 -193.915 ;
        RECT 108.360 -194.115 108.570 -194.080 ;
        RECT 105.415 -194.285 108.570 -194.115 ;
        RECT 110.115 -194.185 110.285 -193.390 ;
        RECT 110.605 -194.105 110.775 -193.645 ;
        RECT 107.695 -194.395 108.570 -194.285 ;
        RECT 109.555 -194.395 110.395 -194.355 ;
        RECT 104.915 -194.850 105.775 -194.480 ;
        RECT 107.695 -194.680 110.395 -194.395 ;
        RECT 101.890 -196.085 102.060 -196.065 ;
        RECT 102.870 -196.085 103.040 -195.125 ;
        RECT 103.850 -196.085 104.020 -195.125 ;
        RECT 104.325 -195.720 104.695 -194.880 ;
        RECT 104.915 -195.585 105.150 -194.850 ;
        RECT 107.695 -195.120 108.570 -194.680 ;
        RECT 109.555 -194.725 110.395 -194.680 ;
        RECT 110.575 -194.570 110.805 -194.105 ;
        RECT 111.095 -194.185 111.265 -193.390 ;
        RECT 111.585 -194.105 111.755 -193.645 ;
        RECT 111.555 -194.570 111.785 -194.105 ;
        RECT 112.075 -194.185 112.245 -193.390 ;
        RECT 112.565 -194.105 112.735 -193.645 ;
        RECT 112.535 -194.410 112.765 -194.105 ;
        RECT 112.535 -194.465 112.915 -194.410 ;
        RECT 113.165 -194.465 113.465 -193.890 ;
        RECT 114.900 -194.185 115.070 -193.390 ;
        RECT 115.390 -194.105 115.560 -193.645 ;
        RECT 112.535 -194.570 113.490 -194.465 ;
        RECT 110.575 -194.690 113.490 -194.570 ;
        RECT 105.430 -195.290 108.570 -195.120 ;
        RECT 105.430 -195.550 105.610 -195.290 ;
        RECT 106.420 -195.470 106.600 -195.290 ;
        RECT 104.945 -195.955 105.115 -195.585 ;
        RECT 104.940 -196.180 105.120 -195.955 ;
        RECT 105.435 -196.010 105.605 -195.550 ;
        RECT 105.925 -195.905 106.095 -195.470 ;
        RECT 106.415 -195.560 106.600 -195.470 ;
        RECT 105.920 -196.180 106.130 -195.905 ;
        RECT 106.415 -196.010 106.585 -195.560 ;
        RECT 106.905 -195.900 107.075 -195.470 ;
        RECT 107.390 -195.560 107.570 -195.290 ;
        RECT 106.890 -196.180 107.100 -195.900 ;
        RECT 107.395 -196.010 107.565 -195.560 ;
        RECT 107.885 -195.925 108.055 -195.470 ;
        RECT 108.360 -195.510 108.570 -195.290 ;
        RECT 110.575 -194.760 112.915 -194.690 ;
        RECT 110.575 -194.800 112.765 -194.760 ;
        RECT 107.870 -196.180 108.080 -195.925 ;
        RECT 108.375 -196.010 108.545 -195.510 ;
        RECT 110.575 -196.065 110.805 -194.800 ;
        RECT 111.555 -195.125 111.785 -194.800 ;
        RECT 112.535 -195.125 112.765 -194.800 ;
        RECT 110.605 -196.085 110.775 -196.065 ;
        RECT 111.585 -196.085 111.755 -195.125 ;
        RECT 112.565 -196.085 112.735 -195.125 ;
        RECT 113.265 -195.360 113.490 -194.690 ;
        RECT 115.360 -194.570 115.590 -194.105 ;
        RECT 115.880 -194.185 116.050 -193.390 ;
        RECT 116.370 -194.105 116.540 -193.645 ;
        RECT 116.340 -194.570 116.570 -194.105 ;
        RECT 116.860 -194.185 117.030 -193.390 ;
        RECT 118.420 -193.455 118.640 -193.165 ;
        RECT 117.350 -194.105 117.520 -193.645 ;
        RECT 118.445 -193.805 118.615 -193.455 ;
        RECT 117.320 -194.410 117.550 -194.105 ;
        RECT 117.320 -194.570 118.190 -194.410 ;
        RECT 115.360 -194.760 118.190 -194.570 ;
        RECT 115.360 -194.800 117.550 -194.760 ;
        RECT 114.285 -195.360 114.570 -195.155 ;
        RECT 113.265 -195.585 114.570 -195.360 ;
        RECT 114.285 -195.975 114.570 -195.585 ;
        RECT 115.360 -196.065 115.590 -194.800 ;
        RECT 116.340 -195.125 116.570 -194.800 ;
        RECT 117.320 -195.125 117.550 -194.800 ;
        RECT 117.825 -194.880 118.190 -194.760 ;
        RECT 118.415 -194.480 118.650 -193.805 ;
        RECT 118.935 -193.910 119.105 -193.395 ;
        RECT 119.400 -193.510 119.620 -193.165 ;
        RECT 118.915 -194.115 119.120 -193.910 ;
        RECT 119.425 -193.935 119.595 -193.510 ;
        RECT 119.915 -193.870 120.085 -193.395 ;
        RECT 120.380 -193.510 120.600 -193.165 ;
        RECT 119.905 -194.115 120.110 -193.870 ;
        RECT 120.405 -193.935 120.575 -193.510 ;
        RECT 120.895 -193.870 121.065 -193.395 ;
        RECT 121.365 -193.455 121.585 -193.165 ;
        RECT 123.570 -193.390 126.240 -193.050 ;
        RECT 120.875 -194.115 121.080 -193.870 ;
        RECT 121.385 -193.935 121.555 -193.455 ;
        RECT 121.875 -193.865 122.045 -193.395 ;
        RECT 121.860 -194.080 122.065 -193.865 ;
        RECT 121.860 -194.115 122.070 -194.080 ;
        RECT 118.915 -194.285 122.070 -194.115 ;
        RECT 123.615 -194.185 123.785 -193.390 ;
        RECT 124.105 -194.105 124.275 -193.645 ;
        RECT 121.195 -194.430 122.070 -194.285 ;
        RECT 123.055 -194.430 123.895 -194.355 ;
        RECT 118.415 -194.850 119.275 -194.480 ;
        RECT 121.195 -194.695 123.895 -194.430 ;
        RECT 115.390 -196.085 115.560 -196.065 ;
        RECT 116.370 -196.085 116.540 -195.125 ;
        RECT 117.350 -196.085 117.520 -195.125 ;
        RECT 117.825 -195.720 118.195 -194.880 ;
        RECT 118.415 -195.585 118.650 -194.850 ;
        RECT 121.195 -195.120 122.070 -194.695 ;
        RECT 123.055 -194.725 123.895 -194.695 ;
        RECT 124.075 -194.570 124.305 -194.105 ;
        RECT 124.595 -194.185 124.765 -193.390 ;
        RECT 125.085 -194.105 125.255 -193.645 ;
        RECT 125.055 -194.570 125.285 -194.105 ;
        RECT 125.575 -194.185 125.745 -193.390 ;
        RECT 126.065 -194.105 126.235 -193.645 ;
        RECT 126.035 -194.410 126.265 -194.105 ;
        RECT 126.035 -194.520 126.415 -194.410 ;
        RECT 126.590 -194.520 126.830 -192.730 ;
        RECT 138.640 -193.055 138.810 -191.335 ;
        RECT 139.620 -193.055 139.790 -191.335 ;
        RECT 141.685 -191.870 141.855 -191.330 ;
        RECT 142.665 -191.870 142.835 -191.330 ;
        RECT 141.095 -192.105 141.460 -192.040 ;
        RECT 140.595 -192.245 141.460 -192.105 ;
        RECT 140.485 -192.310 141.460 -192.245 ;
        RECT 140.485 -193.055 140.790 -192.310 ;
        RECT 141.095 -192.340 141.460 -192.310 ;
        RECT 143.645 -192.190 143.815 -191.330 ;
        RECT 138.640 -193.205 140.790 -193.055 ;
        RECT 138.640 -193.245 140.735 -193.205 ;
        RECT 141.685 -193.265 141.855 -192.485 ;
        RECT 142.175 -193.025 142.345 -192.485 ;
        RECT 142.665 -193.265 142.835 -192.485 ;
        RECT 143.155 -193.025 143.325 -192.485 ;
        RECT 143.645 -192.540 145.035 -192.190 ;
        RECT 136.860 -193.610 137.995 -193.600 ;
        RECT 140.050 -193.610 140.420 -193.480 ;
        RECT 136.860 -193.800 140.420 -193.610 ;
        RECT 140.985 -193.695 144.060 -193.265 ;
        RECT 126.035 -194.570 126.830 -194.520 ;
        RECT 124.075 -194.705 126.830 -194.570 ;
        RECT 124.075 -194.715 126.825 -194.705 ;
        RECT 118.930 -195.290 122.070 -195.120 ;
        RECT 118.930 -195.550 119.110 -195.290 ;
        RECT 119.920 -195.470 120.100 -195.290 ;
        RECT 118.445 -195.955 118.615 -195.585 ;
        RECT 104.940 -196.350 108.080 -196.180 ;
        RECT 118.440 -196.180 118.620 -195.955 ;
        RECT 118.935 -196.010 119.105 -195.550 ;
        RECT 119.425 -195.905 119.595 -195.470 ;
        RECT 119.915 -195.560 120.100 -195.470 ;
        RECT 119.420 -196.180 119.630 -195.905 ;
        RECT 119.915 -196.010 120.085 -195.560 ;
        RECT 120.405 -195.900 120.575 -195.470 ;
        RECT 120.890 -195.560 121.070 -195.290 ;
        RECT 120.390 -196.180 120.600 -195.900 ;
        RECT 120.895 -196.010 121.065 -195.560 ;
        RECT 121.385 -195.925 121.555 -195.470 ;
        RECT 121.860 -195.510 122.070 -195.290 ;
        RECT 124.075 -194.760 126.415 -194.715 ;
        RECT 124.075 -194.800 126.265 -194.760 ;
        RECT 121.370 -196.180 121.580 -195.925 ;
        RECT 121.875 -196.010 122.045 -195.510 ;
        RECT 124.075 -196.065 124.305 -194.800 ;
        RECT 125.055 -195.125 125.285 -194.800 ;
        RECT 126.035 -195.125 126.265 -194.800 ;
        RECT 124.105 -196.085 124.275 -196.065 ;
        RECT 125.085 -196.085 125.255 -195.125 ;
        RECT 126.065 -196.085 126.235 -195.125 ;
        RECT 118.440 -196.350 121.580 -196.180 ;
        RECT 107.105 -197.855 107.905 -197.195 ;
        RECT 107.140 -198.770 107.815 -197.855 ;
        RECT 111.895 -198.465 126.515 -197.980 ;
        RECT 107.090 -199.430 107.890 -198.770 ;
        RECT 109.705 -201.025 109.875 -198.805 ;
        RECT 110.685 -201.025 110.855 -198.805 ;
        RECT 109.705 -201.030 110.855 -201.025 ;
        RECT 106.575 -201.095 107.235 -201.045 ;
        RECT 108.790 -201.090 109.465 -201.060 ;
        RECT 108.690 -201.095 109.465 -201.090 ;
        RECT 106.575 -201.275 109.465 -201.095 ;
        RECT 109.705 -201.215 110.925 -201.030 ;
        RECT 106.575 -201.345 107.235 -201.275 ;
        RECT 108.690 -201.290 109.465 -201.275 ;
        RECT 108.790 -201.330 109.465 -201.290 ;
        RECT 110.755 -201.390 110.925 -201.215 ;
        RECT 111.405 -201.390 111.705 -201.090 ;
        RECT 99.430 -201.755 107.410 -201.540 ;
        RECT 90.185 -201.865 107.410 -201.755 ;
        RECT 108.340 -201.555 109.135 -201.550 ;
        RECT 108.340 -201.580 109.140 -201.555 ;
        RECT 109.880 -201.580 110.555 -201.550 ;
        RECT 108.340 -201.775 110.555 -201.580 ;
        RECT 108.340 -201.780 109.410 -201.775 ;
        RECT 108.340 -201.845 109.140 -201.780 ;
        RECT 109.880 -201.820 110.555 -201.775 ;
        RECT 110.755 -201.695 111.705 -201.390 ;
        RECT 108.340 -201.850 109.135 -201.845 ;
        RECT 90.185 -202.200 100.330 -201.865 ;
        RECT 47.325 -202.470 47.620 -202.435 ;
        RECT 47.325 -202.885 67.205 -202.470 ;
        RECT 47.325 -202.910 47.620 -202.885 ;
        RECT 36.715 -203.535 40.460 -203.490 ;
        RECT 31.295 -203.800 40.460 -203.535 ;
        RECT 27.345 -205.760 28.580 -205.755 ;
        RECT 29.390 -205.760 29.560 -203.905 ;
        RECT 31.295 -204.415 31.490 -203.800 ;
        RECT 37.300 -203.970 40.460 -203.800 ;
        RECT 31.805 -204.170 36.845 -203.990 ;
        RECT 31.315 -205.360 31.485 -204.415 ;
        RECT 25.315 -205.930 26.480 -205.760 ;
        RECT 27.345 -205.930 29.560 -205.760 ;
        RECT 31.305 -205.775 31.490 -205.360 ;
        RECT 31.805 -205.395 31.975 -204.170 ;
        RECT 33.385 -205.365 33.555 -204.355 ;
        RECT 33.875 -205.350 34.045 -204.355 ;
        RECT 35.195 -205.350 35.365 -204.355 ;
        RECT 33.370 -205.470 33.555 -205.365 ;
        RECT 32.775 -205.655 33.555 -205.470 ;
        RECT 33.865 -205.545 35.365 -205.350 ;
        RECT 32.775 -205.775 32.960 -205.655 ;
        RECT 23.595 -206.200 24.270 -206.165 ;
        RECT 26.295 -206.200 26.480 -205.930 ;
        RECT 31.305 -205.960 32.960 -205.775 ;
        RECT 35.685 -205.810 35.855 -204.355 ;
        RECT 36.665 -204.440 36.845 -204.170 ;
        RECT 36.665 -205.395 36.835 -204.440 ;
        RECT 37.155 -205.810 37.325 -204.355 ;
        RECT 38.215 -205.310 38.385 -204.355 ;
        RECT 38.680 -204.390 38.895 -203.970 ;
        RECT 38.190 -205.535 38.405 -205.310 ;
        RECT 38.705 -205.395 38.875 -204.390 ;
        RECT 39.760 -205.300 39.930 -204.355 ;
        RECT 40.225 -204.400 40.440 -203.970 ;
        RECT 37.710 -205.765 38.405 -205.535 ;
        RECT 34.520 -205.980 37.325 -205.810 ;
        RECT 23.595 -206.385 26.480 -206.200 ;
        RECT 23.595 -206.435 24.270 -206.385 ;
        RECT 26.295 -207.075 26.480 -206.385 ;
        RECT 26.650 -206.210 27.325 -206.175 ;
        RECT 26.650 -206.380 30.745 -206.210 ;
        RECT 34.520 -206.290 34.690 -205.980 ;
        RECT 26.650 -206.445 27.325 -206.380 ;
        RECT 27.590 -206.600 28.265 -206.565 ;
        RECT 27.590 -206.790 30.395 -206.600 ;
        RECT 27.590 -206.835 28.265 -206.790 ;
        RECT 29.265 -207.020 29.945 -206.975 ;
        RECT 26.295 -207.260 29.070 -207.075 ;
        RECT 29.265 -207.205 30.040 -207.020 ;
        RECT 29.270 -207.245 29.945 -207.205 ;
        RECT 26.940 -208.480 27.110 -207.260 ;
        RECT 27.920 -208.480 28.090 -207.260 ;
        RECT 28.900 -208.480 29.070 -207.260 ;
        RECT -8.105 -214.125 14.155 -213.945 ;
        RECT 14.465 -213.725 21.975 -213.555 ;
        RECT 30.225 -213.635 30.395 -206.790 ;
        RECT -8.105 -214.365 -7.860 -214.125 ;
        RECT 3.945 -214.345 4.625 -214.300 ;
        RECT 14.465 -214.345 14.635 -213.725 ;
        RECT 28.695 -213.805 30.395 -213.635 ;
        RECT 14.860 -214.000 15.540 -213.985 ;
        RECT 28.695 -214.000 28.865 -213.805 ;
        RECT 14.860 -214.170 28.865 -214.000 ;
        RECT 29.385 -214.095 30.065 -214.065 ;
        RECT 30.575 -214.095 30.745 -206.380 ;
        RECT 31.310 -206.635 32.005 -206.365 ;
        RECT 33.960 -206.460 34.690 -206.290 ;
        RECT 33.960 -207.035 34.130 -206.460 ;
        RECT 35.055 -206.485 35.750 -206.215 ;
        RECT 31.060 -207.205 34.130 -207.035 ;
        RECT 34.435 -206.840 36.835 -206.670 ;
        RECT 31.315 -208.945 31.485 -207.385 ;
        RECT 31.805 -208.425 31.975 -207.205 ;
        RECT 32.295 -208.945 32.465 -207.385 ;
        RECT 32.895 -208.600 33.065 -207.385 ;
        RECT 33.385 -208.425 33.555 -207.205 ;
        RECT 33.875 -208.600 34.045 -207.385 ;
        RECT 34.435 -208.600 34.605 -206.840 ;
        RECT 32.895 -208.770 34.605 -208.600 ;
        RECT 34.785 -207.210 35.855 -207.040 ;
        RECT 34.785 -208.945 34.955 -207.210 ;
        RECT 35.685 -208.425 35.855 -207.210 ;
        RECT 36.665 -208.425 36.835 -206.840 ;
        RECT 37.100 -206.855 37.795 -206.585 ;
        RECT 38.190 -207.460 38.405 -205.765 ;
        RECT 39.740 -206.255 39.955 -205.300 ;
        RECT 40.250 -205.395 40.420 -204.400 ;
        RECT 41.205 -204.705 46.980 -203.400 ;
        RECT 63.890 -203.830 65.315 -203.540 ;
        RECT 66.790 -203.830 67.205 -202.885 ;
        RECT 90.830 -202.960 91.050 -202.200 ;
        RECT 90.850 -203.755 91.020 -202.960 ;
        RECT 91.340 -203.710 91.510 -202.715 ;
        RECT 91.800 -202.955 92.020 -202.200 ;
        RECT 63.890 -203.970 88.690 -203.830 ;
        RECT 90.380 -203.970 91.110 -203.930 ;
        RECT 63.890 -204.150 91.110 -203.970 ;
        RECT 91.315 -203.955 91.540 -203.710 ;
        RECT 91.830 -203.755 92.000 -202.955 ;
        RECT 95.560 -202.960 95.780 -202.200 ;
        RECT 95.580 -203.755 95.750 -202.960 ;
        RECT 96.070 -203.710 96.240 -202.715 ;
        RECT 96.530 -202.955 96.750 -202.200 ;
        RECT 91.315 -203.960 93.285 -203.955 ;
        RECT 91.315 -204.135 93.530 -203.960 ;
        RECT 95.110 -203.970 95.840 -203.930 ;
        RECT 63.890 -204.300 88.690 -204.150 ;
        RECT 90.380 -204.230 91.110 -204.150 ;
        RECT 92.590 -204.180 93.530 -204.135 ;
        RECT 94.815 -204.150 95.840 -203.970 ;
        RECT 96.045 -203.955 96.270 -203.710 ;
        RECT 96.560 -203.755 96.730 -202.955 ;
        RECT 96.045 -204.135 99.395 -203.955 ;
        RECT 92.870 -204.260 93.530 -204.180 ;
        RECT 95.110 -204.230 95.840 -204.150 ;
        RECT 97.320 -204.180 99.395 -204.135 ;
        RECT 63.890 -204.635 65.315 -204.300 ;
        RECT 91.495 -204.415 92.210 -204.330 ;
        RECT 89.205 -204.595 92.210 -204.415 ;
        RECT 39.240 -206.485 39.955 -206.255 ;
        RECT 38.215 -208.425 38.385 -207.460 ;
        RECT 39.740 -207.470 39.955 -206.485 ;
        RECT 40.175 -206.825 40.870 -206.555 ;
        RECT 39.760 -208.425 39.930 -207.470 ;
        RECT 31.315 -209.115 34.955 -208.945 ;
        RECT 14.860 -214.215 15.540 -214.170 ;
        RECT 29.385 -214.265 30.745 -214.095 ;
        RECT 29.385 -214.295 30.065 -214.265 ;
        RECT -8.540 -214.595 -7.860 -214.365 ;
        RECT 3.780 -214.515 14.635 -214.345 ;
        RECT 3.945 -214.530 4.625 -214.515 ;
        RECT 41.205 -214.680 42.510 -204.705 ;
        RECT 45.675 -208.675 46.980 -204.705 ;
        RECT 89.205 -204.860 89.385 -204.595 ;
        RECT 91.495 -204.630 92.210 -204.595 ;
        RECT 68.800 -205.670 89.385 -204.860 ;
        RECT 90.845 -205.005 92.585 -204.825 ;
        RECT 90.845 -205.200 91.025 -205.005 ;
        RECT 48.090 -206.485 48.435 -206.395 ;
        RECT 74.155 -206.485 74.710 -205.670 ;
        RECT 48.090 -207.040 74.710 -206.485 ;
        RECT 48.090 -207.090 48.435 -207.040 ;
        RECT 90.850 -207.215 91.020 -205.200 ;
        RECT 91.905 -207.075 92.075 -205.175 ;
        RECT 92.360 -205.225 92.585 -205.005 ;
        RECT 91.870 -207.395 92.100 -207.075 ;
        RECT 92.395 -207.215 92.565 -205.225 ;
        RECT 92.870 -205.405 93.120 -204.260 ;
        RECT 96.225 -204.415 96.940 -204.330 ;
        RECT 94.810 -204.595 96.940 -204.415 ;
        RECT 96.225 -204.630 96.940 -204.595 ;
        RECT 95.575 -205.005 97.315 -204.825 ;
        RECT 95.575 -205.200 95.755 -205.005 ;
        RECT 92.885 -207.075 93.055 -205.405 ;
        RECT 92.860 -207.395 93.090 -207.075 ;
        RECT 95.580 -207.215 95.750 -205.200 ;
        RECT 96.635 -207.075 96.805 -205.175 ;
        RECT 97.090 -205.225 97.315 -205.005 ;
        RECT 91.870 -207.585 93.090 -207.395 ;
        RECT 96.600 -207.395 96.830 -207.075 ;
        RECT 97.125 -207.215 97.295 -205.225 ;
        RECT 97.600 -205.405 97.850 -204.180 ;
        RECT 97.615 -207.075 97.785 -205.405 ;
        RECT 98.050 -205.505 98.350 -204.675 ;
        RECT 99.225 -205.115 99.395 -204.180 ;
        RECT 99.670 -204.665 99.840 -202.810 ;
        RECT 100.160 -204.350 100.330 -202.200 ;
        RECT 101.220 -202.315 103.425 -202.145 ;
        RECT 101.220 -202.330 102.375 -202.315 ;
        RECT 100.650 -204.660 100.820 -202.810 ;
        RECT 101.220 -202.850 101.395 -202.330 ;
        RECT 101.220 -204.345 101.390 -202.850 ;
        RECT 101.710 -204.345 101.880 -202.805 ;
        RECT 102.200 -202.860 102.375 -202.330 ;
        RECT 102.200 -204.345 102.370 -202.860 ;
        RECT 101.710 -204.660 101.885 -204.345 ;
        RECT 100.650 -204.665 101.885 -204.660 ;
        RECT 102.765 -204.665 102.935 -202.805 ;
        RECT 103.255 -204.345 103.425 -202.315 ;
        RECT 103.745 -204.665 103.915 -202.805 ;
        RECT 105.320 -203.845 105.490 -201.865 ;
        RECT 105.830 -201.945 107.410 -201.865 ;
        RECT 105.830 -202.120 107.405 -201.945 ;
        RECT 99.670 -204.835 101.885 -204.665 ;
        RECT 102.750 -204.835 103.915 -204.665 ;
        RECT 105.810 -204.770 105.980 -202.805 ;
        RECT 107.000 -203.650 107.405 -202.120 ;
        RECT 109.215 -203.635 109.385 -202.075 ;
        RECT 109.705 -203.215 109.875 -202.075 ;
        RECT 110.265 -203.215 110.435 -202.075 ;
        RECT 110.755 -203.115 110.925 -201.695 ;
        RECT 111.405 -201.760 111.705 -201.695 ;
        RECT 109.705 -203.390 110.435 -203.215 ;
        RECT 109.050 -203.650 111.445 -203.635 ;
        RECT 111.895 -203.650 112.245 -198.465 ;
        RECT 107.000 -204.440 112.245 -203.650 ;
        RECT 108.920 -204.655 112.245 -204.440 ;
        RECT 112.530 -202.860 112.880 -199.190 ;
        RECT 113.365 -202.570 113.535 -198.465 ;
        RECT 113.855 -202.850 114.025 -199.030 ;
        RECT 115.365 -202.570 115.535 -198.465 ;
        RECT 115.015 -202.850 115.685 -202.785 ;
        RECT 112.530 -203.130 113.675 -202.860 ;
        RECT 113.855 -203.020 115.685 -202.850 ;
        RECT 101.905 -205.115 102.580 -205.080 ;
        RECT 99.200 -205.285 102.580 -205.115 ;
        RECT 101.905 -205.350 102.580 -205.285 ;
        RECT 102.750 -205.105 102.935 -204.835 ;
        RECT 105.810 -204.950 107.195 -204.770 ;
        RECT 104.960 -205.105 105.635 -205.070 ;
        RECT 102.750 -205.290 105.635 -205.105 ;
        RECT 100.965 -205.505 101.640 -205.470 ;
        RECT 98.050 -205.695 101.640 -205.505 ;
        RECT 100.965 -205.740 101.640 -205.695 ;
        RECT 99.285 -205.925 99.960 -205.880 ;
        RECT 98.625 -206.100 99.960 -205.925 ;
        RECT 102.750 -205.980 102.935 -205.290 ;
        RECT 104.960 -205.340 105.635 -205.290 ;
        RECT 98.625 -206.585 98.925 -206.100 ;
        RECT 99.190 -206.110 99.960 -206.100 ;
        RECT 99.285 -206.150 99.960 -206.110 ;
        RECT 100.160 -206.165 102.935 -205.980 ;
        RECT 97.590 -207.395 97.820 -207.075 ;
        RECT 100.160 -207.385 100.330 -206.165 ;
        RECT 101.140 -207.385 101.310 -206.165 ;
        RECT 102.120 -207.385 102.290 -206.165 ;
        RECT 105.810 -207.385 105.980 -204.950 ;
        RECT 106.540 -205.070 107.195 -204.950 ;
        RECT 108.965 -205.450 109.135 -204.655 ;
        RECT 109.455 -205.370 109.625 -204.910 ;
        RECT 108.405 -205.990 109.245 -205.620 ;
        RECT 109.425 -205.835 109.655 -205.370 ;
        RECT 109.945 -205.450 110.115 -204.655 ;
        RECT 110.435 -205.370 110.605 -204.910 ;
        RECT 110.405 -205.835 110.635 -205.370 ;
        RECT 110.925 -205.450 111.095 -204.655 ;
        RECT 111.415 -205.370 111.585 -204.910 ;
        RECT 111.385 -205.675 111.615 -205.370 ;
        RECT 112.530 -205.675 112.880 -203.130 ;
        RECT 111.385 -205.835 112.880 -205.675 ;
        RECT 109.425 -206.025 112.880 -205.835 ;
        RECT 109.425 -206.065 111.615 -206.025 ;
        RECT 109.425 -207.330 109.655 -206.065 ;
        RECT 110.405 -206.390 110.635 -206.065 ;
        RECT 111.385 -206.390 111.615 -206.065 ;
        RECT 109.455 -207.350 109.625 -207.330 ;
        RECT 110.435 -207.350 110.605 -206.390 ;
        RECT 111.415 -207.350 111.585 -206.390 ;
        RECT 113.855 -206.995 114.025 -203.020 ;
        RECT 115.015 -203.055 115.685 -203.020 ;
        RECT 115.855 -202.800 116.025 -199.030 ;
        RECT 116.395 -202.800 116.985 -202.740 ;
        RECT 115.855 -202.970 116.985 -202.800 ;
        RECT 115.855 -206.995 116.025 -202.970 ;
        RECT 116.395 -203.030 116.985 -202.970 ;
        RECT 117.750 -202.850 118.100 -201.945 ;
        RECT 118.365 -202.570 118.535 -198.465 ;
        RECT 117.750 -203.120 118.620 -202.850 ;
        RECT 118.855 -202.900 119.025 -199.030 ;
        RECT 120.365 -202.570 120.535 -198.465 ;
        RECT 120.015 -202.900 120.685 -202.860 ;
        RECT 118.855 -203.095 120.685 -202.900 ;
        RECT 118.855 -206.995 119.025 -203.095 ;
        RECT 120.015 -203.130 120.685 -203.095 ;
        RECT 120.855 -202.935 121.025 -199.030 ;
        RECT 121.780 -202.935 122.370 -202.875 ;
        RECT 120.855 -203.105 122.370 -202.935 ;
        RECT 120.855 -206.995 121.025 -203.105 ;
        RECT 121.780 -203.165 122.370 -203.105 ;
        RECT 122.705 -202.885 123.055 -201.950 ;
        RECT 123.365 -202.570 123.535 -198.465 ;
        RECT 122.705 -203.155 123.620 -202.885 ;
        RECT 123.855 -202.905 124.025 -199.030 ;
        RECT 125.365 -202.570 125.535 -198.465 ;
        RECT 125.855 -202.855 126.025 -199.030 ;
        RECT 136.915 -199.160 137.295 -193.800 ;
        RECT 137.990 -193.805 140.420 -193.800 ;
        RECT 137.990 -193.810 138.345 -193.805 ;
        RECT 140.050 -193.835 140.420 -193.805 ;
        RECT 138.150 -195.560 138.320 -194.020 ;
        RECT 138.640 -195.560 138.810 -194.020 ;
        RECT 139.130 -195.560 139.300 -194.020 ;
        RECT 139.620 -195.560 139.790 -194.020 ;
        RECT 140.110 -195.560 140.280 -194.020 ;
        RECT 138.635 -195.820 138.810 -195.560 ;
        RECT 142.205 -195.730 142.510 -193.695 ;
        RECT 144.655 -194.515 145.005 -192.540 ;
        RECT 145.875 -193.810 146.045 -190.890 ;
        RECT 146.910 -190.930 147.120 -190.720 ;
        RECT 145.855 -194.105 146.065 -193.810 ;
        RECT 146.930 -193.840 147.100 -190.930 ;
        RECT 147.420 -193.830 147.590 -190.890 ;
        RECT 147.900 -190.940 148.110 -190.720 ;
        RECT 146.915 -194.105 147.125 -193.840 ;
        RECT 145.855 -194.285 147.125 -194.105 ;
        RECT 147.400 -194.100 147.610 -193.830 ;
        RECT 147.910 -193.930 148.080 -190.940 ;
        RECT 148.970 -193.860 149.140 -190.890 ;
        RECT 147.400 -194.295 148.105 -194.100 ;
        RECT 147.890 -194.355 148.105 -194.295 ;
        RECT 146.680 -194.515 147.455 -194.465 ;
        RECT 144.655 -194.695 147.455 -194.515 ;
        RECT 144.655 -194.705 145.005 -194.695 ;
        RECT 146.680 -194.740 147.455 -194.695 ;
        RECT 147.890 -194.630 148.795 -194.355 ;
        RECT 147.890 -194.980 148.105 -194.630 ;
        RECT 145.330 -195.050 146.105 -195.005 ;
        RECT 145.145 -195.220 146.105 -195.050 ;
        RECT 145.330 -195.280 146.105 -195.220 ;
        RECT 146.335 -195.180 148.105 -194.980 ;
        RECT 148.965 -195.080 149.180 -193.860 ;
        RECT 150.150 -194.205 150.500 -187.520 ;
        RECT 180.970 -187.785 181.140 -186.745 ;
        RECT 181.950 -187.785 182.120 -186.745 ;
        RECT 182.930 -187.785 183.100 -186.745 ;
        RECT 185.835 -188.430 186.005 -186.710 ;
        RECT 186.815 -188.430 186.985 -186.710 ;
        RECT 187.680 -187.455 187.985 -186.710 ;
        RECT 188.880 -187.280 189.050 -186.500 ;
        RECT 189.370 -187.280 189.540 -186.740 ;
        RECT 189.860 -187.280 190.030 -186.500 ;
        RECT 223.825 -186.705 225.060 -186.500 ;
        RECT 229.235 -186.640 229.910 -186.600 ;
        RECT 229.135 -186.650 229.910 -186.640 ;
        RECT 190.350 -187.280 190.520 -186.740 ;
        RECT 223.825 -186.790 224.475 -186.705 ;
        RECT 224.695 -186.770 225.060 -186.705 ;
        RECT 228.100 -186.830 229.910 -186.650 ;
        RECT 232.495 -186.695 236.420 -186.265 ;
        RECT 269.815 -186.330 270.465 -185.870 ;
        RECT 271.275 -186.160 271.445 -184.880 ;
        RECT 271.765 -186.160 271.935 -185.120 ;
        RECT 272.255 -186.160 272.425 -184.880 ;
        RECT 272.745 -185.990 272.915 -185.120 ;
        RECT 275.650 -185.770 275.820 -184.230 ;
        RECT 276.140 -185.770 276.310 -184.230 ;
        RECT 276.630 -185.770 276.800 -184.230 ;
        RECT 277.120 -185.770 277.290 -184.230 ;
        RECT 277.610 -185.770 277.780 -184.230 ;
        RECT 275.490 -185.985 275.845 -185.980 ;
        RECT 277.550 -185.985 277.920 -185.955 ;
        RECT 275.490 -185.990 277.920 -185.985 ;
        RECT 272.745 -186.160 277.920 -185.990 ;
        RECT 279.705 -186.095 280.010 -184.060 ;
        RECT 302.945 -184.210 312.200 -183.455 ;
        RECT 318.605 -183.425 321.930 -183.285 ;
        RECT 318.605 -183.715 323.780 -183.425 ;
        RECT 318.605 -184.120 319.035 -183.715 ;
        RECT 319.905 -183.900 320.080 -183.715 ;
        RECT 321.530 -183.730 323.780 -183.715 ;
        RECT 302.945 -184.550 304.825 -184.210 ;
        RECT 310.950 -184.465 312.200 -184.210 ;
        RECT 314.345 -184.550 319.035 -184.120 ;
        RECT 313.585 -186.000 314.235 -185.540 ;
        RECT 315.045 -185.830 315.215 -184.550 ;
        RECT 315.535 -185.830 315.705 -184.790 ;
        RECT 316.025 -185.830 316.195 -184.550 ;
        RECT 316.515 -185.660 316.685 -184.790 ;
        RECT 319.420 -185.440 319.590 -183.900 ;
        RECT 319.910 -185.440 320.080 -183.900 ;
        RECT 320.400 -185.440 320.570 -183.900 ;
        RECT 320.890 -185.440 321.060 -183.900 ;
        RECT 321.380 -185.440 321.550 -183.900 ;
        RECT 319.260 -185.655 319.615 -185.650 ;
        RECT 321.320 -185.655 321.690 -185.625 ;
        RECT 319.260 -185.660 321.690 -185.655 ;
        RECT 316.515 -185.830 321.690 -185.660 ;
        RECT 323.475 -185.765 323.780 -183.730 ;
        RECT 346.825 -183.485 348.515 -183.005 ;
        RECT 365.705 -183.200 367.405 -181.230 ;
        RECT 392.975 -183.180 394.325 -182.575 ;
        RECT 403.040 -183.180 404.515 -182.970 ;
        RECT 412.385 -183.010 413.440 -181.230 ;
        RECT 356.765 -183.485 358.105 -183.280 ;
        RECT 346.825 -184.140 358.105 -183.485 ;
        RECT 364.370 -183.340 367.695 -183.200 ;
        RECT 364.370 -183.630 369.545 -183.340 ;
        RECT 364.370 -184.035 364.800 -183.630 ;
        RECT 365.670 -183.815 365.845 -183.630 ;
        RECT 367.295 -183.645 369.545 -183.630 ;
        RECT 346.825 -184.460 348.515 -184.140 ;
        RECT 356.765 -184.480 358.105 -184.140 ;
        RECT 360.110 -184.465 364.800 -184.035 ;
        RECT 316.520 -185.850 321.690 -185.830 ;
        RECT 316.520 -185.860 319.265 -185.850 ;
        RECT 314.455 -186.000 314.820 -185.970 ;
        RECT 321.320 -185.980 321.690 -185.850 ;
        RECT 272.750 -186.180 277.920 -186.160 ;
        RECT 272.750 -186.190 275.495 -186.180 ;
        RECT 270.685 -186.330 271.050 -186.300 ;
        RECT 277.550 -186.310 277.920 -186.180 ;
        RECT 269.815 -186.535 271.050 -186.330 ;
        RECT 275.225 -186.470 275.900 -186.430 ;
        RECT 275.125 -186.480 275.900 -186.470 ;
        RECT 269.815 -186.620 270.465 -186.535 ;
        RECT 270.685 -186.600 271.050 -186.535 ;
        RECT 274.090 -186.660 275.900 -186.480 ;
        RECT 278.485 -186.525 282.410 -186.095 ;
        RECT 313.585 -186.205 314.820 -186.000 ;
        RECT 318.995 -186.140 319.670 -186.100 ;
        RECT 318.895 -186.150 319.670 -186.140 ;
        RECT 313.585 -186.290 314.235 -186.205 ;
        RECT 314.455 -186.270 314.820 -186.205 ;
        RECT 317.860 -186.330 319.670 -186.150 ;
        RECT 322.255 -186.195 326.180 -185.765 ;
        RECT 359.350 -185.915 360.000 -185.455 ;
        RECT 360.810 -185.745 360.980 -184.465 ;
        RECT 361.300 -185.745 361.470 -184.705 ;
        RECT 361.790 -185.745 361.960 -184.465 ;
        RECT 362.280 -185.575 362.450 -184.705 ;
        RECT 365.185 -185.355 365.355 -183.815 ;
        RECT 365.675 -185.355 365.845 -183.815 ;
        RECT 366.165 -185.355 366.335 -183.815 ;
        RECT 366.655 -185.355 366.825 -183.815 ;
        RECT 367.145 -185.355 367.315 -183.815 ;
        RECT 365.025 -185.570 365.380 -185.565 ;
        RECT 367.085 -185.570 367.455 -185.540 ;
        RECT 365.025 -185.575 367.455 -185.570 ;
        RECT 362.280 -185.745 367.455 -185.575 ;
        RECT 369.240 -185.680 369.545 -183.645 ;
        RECT 392.975 -183.875 404.515 -183.180 ;
        RECT 411.190 -183.150 414.515 -183.010 ;
        RECT 411.190 -183.440 416.365 -183.150 ;
        RECT 411.190 -183.845 411.620 -183.440 ;
        RECT 412.490 -183.625 412.665 -183.440 ;
        RECT 414.115 -183.455 416.365 -183.440 ;
        RECT 392.975 -184.000 394.325 -183.875 ;
        RECT 403.040 -184.335 404.515 -183.875 ;
        RECT 406.930 -184.275 411.620 -183.845 ;
        RECT 362.285 -185.765 367.455 -185.745 ;
        RECT 362.285 -185.775 365.030 -185.765 ;
        RECT 360.220 -185.915 360.585 -185.885 ;
        RECT 367.085 -185.895 367.455 -185.765 ;
        RECT 359.350 -186.120 360.585 -185.915 ;
        RECT 364.760 -186.055 365.435 -186.015 ;
        RECT 364.660 -186.065 365.435 -186.055 ;
        RECT 318.895 -186.340 319.670 -186.330 ;
        RECT 318.995 -186.370 319.670 -186.340 ;
        RECT 319.910 -186.255 322.005 -186.215 ;
        RECT 319.910 -186.405 322.060 -186.255 ;
        RECT 275.125 -186.670 275.900 -186.660 ;
        RECT 229.135 -186.840 229.910 -186.830 ;
        RECT 229.235 -186.870 229.910 -186.840 ;
        RECT 230.150 -186.755 232.245 -186.715 ;
        RECT 230.150 -186.905 232.300 -186.755 ;
        RECT 188.290 -187.455 188.655 -187.425 ;
        RECT 187.680 -187.520 188.655 -187.455 ;
        RECT 187.790 -187.660 188.655 -187.520 ;
        RECT 188.290 -187.725 188.655 -187.660 ;
        RECT 190.840 -187.575 192.700 -187.225 ;
        RECT 188.880 -188.435 189.050 -187.895 ;
        RECT 189.860 -188.435 190.030 -187.895 ;
        RECT 190.840 -188.435 191.010 -187.575 ;
        RECT 156.730 -190.000 158.335 -189.830 ;
        RECT 155.835 -192.680 156.005 -190.180 ;
        RECT 155.830 -192.910 156.005 -192.680 ;
        RECT 156.730 -192.910 156.930 -190.000 ;
        RECT 157.175 -190.200 157.350 -190.000 ;
        RECT 157.180 -192.720 157.350 -190.200 ;
        RECT 157.670 -192.685 157.840 -190.180 ;
        RECT 158.160 -190.195 158.335 -190.000 ;
        RECT 155.830 -193.110 156.930 -192.910 ;
        RECT 157.655 -193.285 157.845 -192.685 ;
        RECT 158.160 -192.720 158.330 -190.195 ;
        RECT 158.810 -193.100 158.980 -190.180 ;
        RECT 160.440 -192.750 160.610 -190.180 ;
        RECT 161.580 -191.630 161.750 -190.180 ;
        RECT 189.110 -190.775 190.310 -190.605 ;
        RECT 161.575 -192.095 161.760 -191.630 ;
        RECT 161.575 -192.280 162.260 -192.095 ;
        RECT 160.440 -192.920 161.235 -192.750 ;
        RECT 159.555 -193.100 160.245 -193.045 ;
        RECT 155.835 -193.475 157.845 -193.285 ;
        RECT 158.180 -193.270 160.245 -193.100 ;
        RECT 154.650 -193.530 155.340 -193.480 ;
        RECT 152.700 -193.700 155.340 -193.530 ;
        RECT 150.095 -194.565 150.620 -194.205 ;
        RECT 152.700 -195.080 152.915 -193.700 ;
        RECT 154.650 -193.750 155.340 -193.700 ;
        RECT 154.930 -194.205 155.620 -194.160 ;
        RECT 153.880 -194.375 155.620 -194.205 ;
        RECT 153.880 -195.010 154.240 -194.375 ;
        RECT 154.930 -194.430 155.620 -194.375 ;
        RECT 153.880 -195.055 154.300 -195.010 ;
        RECT 140.260 -195.820 142.510 -195.730 ;
        RECT 138.050 -196.035 142.510 -195.820 ;
        RECT 138.050 -196.125 140.295 -196.035 ;
        RECT 142.205 -197.510 142.510 -196.035 ;
        RECT 145.875 -196.920 146.045 -195.450 ;
        RECT 146.335 -195.530 146.560 -195.180 ;
        RECT 148.295 -195.280 152.915 -195.080 ;
        RECT 148.535 -195.295 152.915 -195.280 ;
        RECT 145.840 -197.510 146.075 -196.920 ;
        RECT 146.365 -196.990 146.535 -195.530 ;
        RECT 146.855 -196.915 147.025 -195.450 ;
        RECT 148.065 -196.865 148.235 -195.450 ;
        RECT 148.535 -195.495 148.755 -195.295 ;
        RECT 153.905 -195.405 154.300 -195.055 ;
        RECT 146.820 -197.510 147.055 -196.915 ;
        RECT 148.030 -197.510 148.265 -196.865 ;
        RECT 148.555 -196.990 148.725 -195.495 ;
        RECT 155.345 -196.615 155.515 -195.160 ;
        RECT 155.335 -197.170 155.520 -196.615 ;
        RECT 155.835 -196.700 156.005 -193.475 ;
        RECT 156.980 -193.825 157.170 -193.475 ;
        RECT 158.180 -193.665 158.350 -193.270 ;
        RECT 159.555 -193.315 160.245 -193.270 ;
        RECT 156.930 -194.515 157.200 -193.825 ;
        RECT 157.695 -193.835 158.350 -193.665 ;
        RECT 158.680 -193.750 159.370 -193.480 ;
        RECT 160.605 -193.825 160.875 -193.135 ;
        RECT 161.065 -193.140 161.235 -192.920 ;
        RECT 161.065 -193.410 161.895 -193.140 ;
        RECT 157.695 -196.700 157.865 -193.835 ;
        RECT 161.065 -193.985 161.235 -193.410 ;
        RECT 161.495 -193.985 161.765 -193.900 ;
        RECT 158.185 -194.180 158.980 -194.005 ;
        RECT 161.065 -194.010 161.765 -193.985 ;
        RECT 160.925 -194.155 161.765 -194.010 ;
        RECT 158.185 -196.700 158.355 -194.180 ;
        RECT 158.810 -196.700 158.980 -194.180 ;
        RECT 159.300 -196.615 159.470 -194.160 ;
        RECT 159.950 -196.610 160.120 -194.160 ;
        RECT 152.650 -197.190 155.705 -197.170 ;
        RECT 159.295 -197.190 159.480 -196.615 ;
        RECT 159.935 -197.190 160.120 -196.610 ;
        RECT 160.440 -196.700 160.610 -194.160 ;
        RECT 160.925 -194.180 161.235 -194.155 ;
        RECT 160.930 -196.700 161.100 -194.180 ;
        RECT 161.495 -194.195 161.765 -194.155 ;
        RECT 162.070 -194.745 162.260 -192.280 ;
        RECT 180.840 -193.110 181.010 -191.390 ;
        RECT 181.820 -193.110 181.990 -191.390 ;
        RECT 183.885 -191.925 184.055 -191.385 ;
        RECT 184.865 -191.925 185.035 -191.385 ;
        RECT 183.295 -192.160 183.660 -192.095 ;
        RECT 182.795 -192.300 183.660 -192.160 ;
        RECT 182.685 -192.365 183.660 -192.300 ;
        RECT 182.685 -193.110 182.990 -192.365 ;
        RECT 183.295 -192.395 183.660 -192.365 ;
        RECT 185.845 -192.245 186.015 -191.385 ;
        RECT 180.840 -193.260 182.990 -193.110 ;
        RECT 180.840 -193.300 182.935 -193.260 ;
        RECT 183.885 -193.320 184.055 -192.540 ;
        RECT 184.375 -193.080 184.545 -192.540 ;
        RECT 184.865 -193.320 185.035 -192.540 ;
        RECT 185.355 -193.080 185.525 -192.540 ;
        RECT 185.845 -192.595 187.235 -192.245 ;
        RECT 179.060 -193.665 180.195 -193.655 ;
        RECT 182.250 -193.665 182.620 -193.535 ;
        RECT 179.060 -193.855 182.620 -193.665 ;
        RECT 183.185 -193.750 186.260 -193.320 ;
        RECT 162.070 -194.935 163.530 -194.745 ;
        RECT 161.580 -196.605 161.750 -195.160 ;
        RECT 162.070 -195.185 162.260 -194.935 ;
        RECT 161.570 -197.190 161.755 -196.605 ;
        RECT 162.070 -196.700 162.240 -195.185 ;
        RECT 152.650 -197.510 162.320 -197.190 ;
        RECT 142.205 -197.735 162.320 -197.510 ;
        RECT 142.205 -198.075 153.215 -197.735 ;
        RECT 154.955 -197.995 162.320 -197.735 ;
        RECT 132.935 -199.440 137.295 -199.160 ;
        RECT 163.340 -199.410 163.530 -194.935 ;
        RECT 179.115 -198.105 179.495 -193.855 ;
        RECT 180.190 -193.860 182.620 -193.855 ;
        RECT 180.190 -193.865 180.545 -193.860 ;
        RECT 182.250 -193.890 182.620 -193.860 ;
        RECT 180.350 -195.615 180.520 -194.075 ;
        RECT 180.840 -195.615 181.010 -194.075 ;
        RECT 181.330 -195.615 181.500 -194.075 ;
        RECT 181.820 -195.615 181.990 -194.075 ;
        RECT 182.310 -195.615 182.480 -194.075 ;
        RECT 180.835 -195.875 181.010 -195.615 ;
        RECT 184.405 -195.785 184.710 -193.750 ;
        RECT 186.855 -194.570 187.205 -192.595 ;
        RECT 188.075 -193.865 188.245 -190.945 ;
        RECT 189.110 -190.985 189.320 -190.775 ;
        RECT 188.055 -194.160 188.265 -193.865 ;
        RECT 189.130 -193.895 189.300 -190.985 ;
        RECT 189.620 -193.885 189.790 -190.945 ;
        RECT 190.100 -190.995 190.310 -190.775 ;
        RECT 189.115 -194.160 189.325 -193.895 ;
        RECT 188.055 -194.340 189.325 -194.160 ;
        RECT 189.600 -194.155 189.810 -193.885 ;
        RECT 190.110 -193.985 190.280 -190.995 ;
        RECT 191.170 -193.915 191.340 -190.945 ;
        RECT 189.600 -194.350 190.305 -194.155 ;
        RECT 190.090 -194.410 190.305 -194.350 ;
        RECT 188.880 -194.570 189.655 -194.520 ;
        RECT 186.855 -194.750 189.655 -194.570 ;
        RECT 186.855 -194.760 187.205 -194.750 ;
        RECT 188.880 -194.795 189.655 -194.750 ;
        RECT 190.090 -194.685 190.995 -194.410 ;
        RECT 190.090 -195.035 190.305 -194.685 ;
        RECT 187.530 -195.105 188.305 -195.060 ;
        RECT 187.345 -195.275 188.305 -195.105 ;
        RECT 187.530 -195.335 188.305 -195.275 ;
        RECT 188.535 -195.235 190.305 -195.035 ;
        RECT 191.165 -195.135 191.380 -193.915 ;
        RECT 192.350 -194.260 192.700 -187.575 ;
        RECT 225.285 -187.980 225.455 -186.940 ;
        RECT 226.265 -187.980 226.435 -186.940 ;
        RECT 227.245 -187.980 227.415 -186.940 ;
        RECT 230.150 -188.625 230.320 -186.905 ;
        RECT 231.130 -188.625 231.300 -186.905 ;
        RECT 231.995 -187.650 232.300 -186.905 ;
        RECT 233.195 -187.475 233.365 -186.695 ;
        RECT 233.685 -187.475 233.855 -186.935 ;
        RECT 234.175 -187.475 234.345 -186.695 ;
        RECT 275.225 -186.700 275.900 -186.670 ;
        RECT 276.140 -186.585 278.235 -186.545 ;
        RECT 276.140 -186.735 278.290 -186.585 ;
        RECT 234.665 -187.475 234.835 -186.935 ;
        RECT 232.605 -187.650 232.970 -187.620 ;
        RECT 231.995 -187.715 232.970 -187.650 ;
        RECT 232.105 -187.855 232.970 -187.715 ;
        RECT 232.605 -187.920 232.970 -187.855 ;
        RECT 235.155 -187.770 237.015 -187.420 ;
        RECT 233.195 -188.630 233.365 -188.090 ;
        RECT 234.175 -188.630 234.345 -188.090 ;
        RECT 235.155 -188.630 235.325 -187.770 ;
        RECT 198.930 -190.055 200.535 -189.885 ;
        RECT 198.035 -192.735 198.205 -190.235 ;
        RECT 198.030 -192.965 198.205 -192.735 ;
        RECT 198.930 -192.965 199.130 -190.055 ;
        RECT 199.375 -190.255 199.550 -190.055 ;
        RECT 199.380 -192.775 199.550 -190.255 ;
        RECT 199.870 -192.740 200.040 -190.235 ;
        RECT 200.360 -190.250 200.535 -190.055 ;
        RECT 198.030 -193.165 199.130 -192.965 ;
        RECT 199.855 -193.340 200.045 -192.740 ;
        RECT 200.360 -192.775 200.530 -190.250 ;
        RECT 201.010 -193.155 201.180 -190.235 ;
        RECT 202.640 -192.805 202.810 -190.235 ;
        RECT 203.780 -191.685 203.950 -190.235 ;
        RECT 233.425 -190.970 234.625 -190.800 ;
        RECT 203.775 -192.150 203.960 -191.685 ;
        RECT 203.775 -192.335 204.460 -192.150 ;
        RECT 202.640 -192.975 203.435 -192.805 ;
        RECT 201.755 -193.155 202.445 -193.100 ;
        RECT 198.035 -193.530 200.045 -193.340 ;
        RECT 200.380 -193.325 202.445 -193.155 ;
        RECT 196.850 -193.585 197.540 -193.535 ;
        RECT 194.900 -193.755 197.540 -193.585 ;
        RECT 192.295 -194.620 192.820 -194.260 ;
        RECT 194.900 -195.135 195.115 -193.755 ;
        RECT 196.850 -193.805 197.540 -193.755 ;
        RECT 197.130 -194.260 197.820 -194.215 ;
        RECT 196.080 -194.430 197.820 -194.260 ;
        RECT 196.080 -195.065 196.440 -194.430 ;
        RECT 197.130 -194.485 197.820 -194.430 ;
        RECT 196.080 -195.110 196.500 -195.065 ;
        RECT 182.460 -195.875 184.710 -195.785 ;
        RECT 180.250 -196.090 184.710 -195.875 ;
        RECT 180.250 -196.180 182.495 -196.090 ;
        RECT 132.935 -199.820 153.465 -199.440 ;
        RECT 132.935 -199.890 137.295 -199.820 ;
        RECT 126.260 -202.855 126.850 -202.815 ;
        RECT 124.980 -202.905 125.650 -202.870 ;
        RECT 123.855 -203.100 125.650 -202.905 ;
        RECT 123.855 -206.995 124.025 -203.100 ;
        RECT 124.980 -203.140 125.650 -203.100 ;
        RECT 125.855 -203.025 126.865 -202.855 ;
        RECT 125.855 -206.995 126.025 -203.025 ;
        RECT 126.260 -203.105 126.850 -203.025 ;
        RECT 96.600 -207.585 97.820 -207.395 ;
        RECT 45.675 -209.980 50.525 -208.675 ;
        RECT 46.415 -212.195 47.155 -211.955 ;
        RECT 45.635 -212.870 46.250 -212.650 ;
        RECT -27.750 -214.790 -24.590 -214.745 ;
        RECT -15.250 -214.790 -12.090 -214.745 ;
        RECT -2.750 -214.790 0.410 -214.745 ;
        RECT 9.750 -214.790 12.910 -214.745 ;
        RECT 22.250 -214.790 25.410 -214.745 ;
        RECT 37.170 -214.790 42.510 -214.680 ;
        RECT -33.755 -214.795 -24.590 -214.790 ;
        RECT -21.255 -214.795 42.510 -214.790 ;
        RECT -33.755 -215.055 42.510 -214.795 ;
        RECT -33.755 -215.670 -33.560 -215.055 ;
        RECT -27.750 -215.225 -21.060 -215.055 ;
        RECT -15.250 -215.225 -12.090 -215.055 ;
        RECT -33.245 -215.425 -28.205 -215.245 ;
        RECT -33.735 -216.615 -33.565 -215.670 ;
        RECT -33.745 -217.030 -33.560 -216.615 ;
        RECT -33.245 -216.650 -33.075 -215.425 ;
        RECT -31.665 -216.620 -31.495 -215.610 ;
        RECT -31.175 -216.605 -31.005 -215.610 ;
        RECT -29.855 -216.605 -29.685 -215.610 ;
        RECT -31.680 -216.725 -31.495 -216.620 ;
        RECT -32.275 -216.910 -31.495 -216.725 ;
        RECT -31.185 -216.800 -29.685 -216.605 ;
        RECT -32.275 -217.030 -32.090 -216.910 ;
        RECT -33.745 -217.215 -32.090 -217.030 ;
        RECT -29.365 -217.065 -29.195 -215.610 ;
        RECT -28.385 -215.695 -28.205 -215.425 ;
        RECT -28.385 -216.650 -28.215 -215.695 ;
        RECT -27.895 -217.065 -27.725 -215.610 ;
        RECT -26.835 -216.565 -26.665 -215.610 ;
        RECT -26.370 -215.645 -26.155 -215.225 ;
        RECT -25.195 -215.230 -21.060 -215.225 ;
        RECT -26.860 -216.790 -26.645 -216.565 ;
        RECT -26.345 -216.650 -26.175 -215.645 ;
        RECT -25.290 -216.555 -25.120 -215.610 ;
        RECT -24.825 -215.655 -24.610 -215.230 ;
        RECT -27.340 -217.020 -26.645 -216.790 ;
        RECT -30.530 -217.235 -27.725 -217.065 ;
        RECT -30.530 -217.545 -30.360 -217.235 ;
        RECT -33.740 -217.890 -33.045 -217.620 ;
        RECT -31.090 -217.715 -30.360 -217.545 ;
        RECT -31.090 -218.290 -30.920 -217.715 ;
        RECT -29.995 -217.740 -29.300 -217.470 ;
        RECT -34.290 -218.460 -30.920 -218.290 ;
        RECT -30.615 -218.095 -28.215 -217.925 ;
        RECT -87.845 -218.615 -84.520 -218.475 ;
        RECT -107.740 -218.890 -104.965 -218.705 ;
        RECT -104.765 -218.825 -95.675 -218.650 ;
        RECT -104.765 -218.835 -103.995 -218.825 ;
        RECT -104.765 -218.875 -104.090 -218.835 ;
        RECT -95.965 -218.850 -95.675 -218.825 ;
        RECT -107.095 -220.110 -106.925 -218.890 ;
        RECT -106.115 -220.110 -105.945 -218.890 ;
        RECT -105.135 -220.110 -104.965 -218.890 ;
        RECT -42.240 -219.430 -41.240 -219.310 ;
        RECT -94.145 -220.110 -41.240 -219.430 ;
        RECT -42.240 -220.165 -41.240 -220.110 ;
        RECT -33.735 -220.200 -33.565 -218.640 ;
        RECT -33.245 -219.680 -33.075 -218.460 ;
        RECT -32.755 -220.200 -32.585 -218.640 ;
        RECT -32.155 -219.855 -31.985 -218.640 ;
        RECT -31.665 -219.680 -31.495 -218.460 ;
        RECT -31.175 -219.855 -31.005 -218.640 ;
        RECT -30.615 -219.855 -30.445 -218.095 ;
        RECT -32.155 -220.025 -30.445 -219.855 ;
        RECT -30.265 -218.465 -29.195 -218.295 ;
        RECT -30.265 -220.200 -30.095 -218.465 ;
        RECT -29.365 -219.680 -29.195 -218.465 ;
        RECT -28.385 -219.680 -28.215 -218.095 ;
        RECT -27.950 -218.110 -27.255 -217.840 ;
        RECT -26.860 -218.715 -26.645 -217.020 ;
        RECT -25.310 -217.510 -25.095 -216.555 ;
        RECT -24.800 -216.650 -24.630 -215.655 ;
        RECT -21.255 -215.670 -21.060 -215.230 ;
        RECT -20.745 -215.425 -15.705 -215.245 ;
        RECT -22.105 -216.475 -21.875 -215.795 ;
        RECT -25.810 -217.740 -25.095 -217.510 ;
        RECT -26.835 -219.680 -26.665 -218.715 ;
        RECT -25.310 -218.725 -25.095 -217.740 ;
        RECT -24.875 -218.080 -24.180 -217.810 ;
        RECT -22.075 -218.290 -21.905 -216.475 ;
        RECT -21.235 -216.615 -21.065 -215.670 ;
        RECT -21.245 -217.030 -21.060 -216.615 ;
        RECT -20.745 -216.650 -20.575 -215.425 ;
        RECT -19.165 -216.620 -18.995 -215.610 ;
        RECT -18.675 -216.605 -18.505 -215.610 ;
        RECT -17.355 -216.605 -17.185 -215.610 ;
        RECT -19.180 -216.725 -18.995 -216.620 ;
        RECT -19.775 -216.910 -18.995 -216.725 ;
        RECT -18.685 -216.800 -17.185 -216.605 ;
        RECT -19.775 -217.030 -19.590 -216.910 ;
        RECT -21.245 -217.215 -19.590 -217.030 ;
        RECT -16.865 -217.065 -16.695 -215.610 ;
        RECT -15.885 -215.695 -15.705 -215.425 ;
        RECT -15.885 -216.650 -15.715 -215.695 ;
        RECT -15.395 -217.065 -15.225 -215.610 ;
        RECT -14.335 -216.565 -14.165 -215.610 ;
        RECT -13.870 -215.645 -13.655 -215.225 ;
        RECT -14.360 -216.790 -14.145 -216.565 ;
        RECT -13.845 -216.650 -13.675 -215.645 ;
        RECT -12.790 -216.555 -12.620 -215.610 ;
        RECT -12.325 -215.655 -12.110 -215.225 ;
        RECT -14.840 -217.020 -14.145 -216.790 ;
        RECT -19.330 -217.370 -18.635 -217.100 ;
        RECT -18.030 -217.235 -15.225 -217.065 ;
        RECT -18.030 -217.545 -17.860 -217.235 ;
        RECT -21.240 -217.890 -20.545 -217.620 ;
        RECT -18.590 -217.715 -17.860 -217.545 ;
        RECT -18.590 -218.290 -18.420 -217.715 ;
        RECT -17.495 -217.740 -16.800 -217.470 ;
        RECT -22.075 -218.460 -18.420 -218.290 ;
        RECT -18.115 -218.095 -15.715 -217.925 ;
        RECT -25.290 -219.680 -25.120 -218.725 ;
        RECT -33.735 -220.370 -30.095 -220.200 ;
        RECT -21.235 -220.200 -21.065 -218.640 ;
        RECT -20.745 -219.680 -20.575 -218.460 ;
        RECT -20.255 -220.200 -20.085 -218.640 ;
        RECT -19.655 -219.855 -19.485 -218.640 ;
        RECT -19.165 -219.680 -18.995 -218.460 ;
        RECT -18.675 -219.855 -18.505 -218.640 ;
        RECT -18.115 -219.855 -17.945 -218.095 ;
        RECT -19.655 -220.025 -17.945 -219.855 ;
        RECT -17.765 -218.465 -16.695 -218.295 ;
        RECT -17.765 -220.200 -17.595 -218.465 ;
        RECT -16.865 -219.680 -16.695 -218.465 ;
        RECT -15.885 -219.680 -15.715 -218.095 ;
        RECT -15.450 -218.110 -14.755 -217.840 ;
        RECT -14.360 -218.715 -14.145 -217.020 ;
        RECT -13.940 -217.340 -13.245 -217.070 ;
        RECT -12.810 -217.510 -12.595 -216.555 ;
        RECT -12.300 -216.650 -12.130 -215.655 ;
        RECT -8.755 -215.670 -8.560 -215.055 ;
        RECT -2.750 -215.225 0.410 -215.055 ;
        RECT -8.245 -215.425 -3.205 -215.245 ;
        RECT -9.365 -216.455 -9.135 -215.775 ;
        RECT -13.310 -217.740 -12.595 -217.510 ;
        RECT -14.335 -219.680 -14.165 -218.715 ;
        RECT -12.810 -218.725 -12.595 -217.740 ;
        RECT -12.375 -218.080 -11.680 -217.810 ;
        RECT -9.335 -218.290 -9.165 -216.455 ;
        RECT -8.735 -216.615 -8.565 -215.670 ;
        RECT -8.745 -217.030 -8.560 -216.615 ;
        RECT -8.245 -216.650 -8.075 -215.425 ;
        RECT -6.665 -216.620 -6.495 -215.610 ;
        RECT -6.175 -216.605 -6.005 -215.610 ;
        RECT -4.855 -216.605 -4.685 -215.610 ;
        RECT -6.680 -216.725 -6.495 -216.620 ;
        RECT -7.275 -216.910 -6.495 -216.725 ;
        RECT -6.185 -216.800 -4.685 -216.605 ;
        RECT -7.275 -217.030 -7.090 -216.910 ;
        RECT -8.745 -217.215 -7.090 -217.030 ;
        RECT -4.365 -217.065 -4.195 -215.610 ;
        RECT -3.385 -215.695 -3.205 -215.425 ;
        RECT -3.385 -216.650 -3.215 -215.695 ;
        RECT -2.895 -217.065 -2.725 -215.610 ;
        RECT -1.835 -216.565 -1.665 -215.610 ;
        RECT -1.370 -215.645 -1.155 -215.225 ;
        RECT -1.860 -216.790 -1.645 -216.565 ;
        RECT -1.345 -216.650 -1.175 -215.645 ;
        RECT -0.290 -216.555 -0.120 -215.610 ;
        RECT 0.175 -215.655 0.390 -215.225 ;
        RECT -2.340 -217.020 -1.645 -216.790 ;
        RECT -6.830 -217.370 -6.135 -217.100 ;
        RECT -5.530 -217.235 -2.725 -217.065 ;
        RECT -5.530 -217.545 -5.360 -217.235 ;
        RECT -8.740 -217.890 -8.045 -217.620 ;
        RECT -6.090 -217.715 -5.360 -217.545 ;
        RECT -6.090 -218.290 -5.920 -217.715 ;
        RECT -4.995 -217.740 -4.300 -217.470 ;
        RECT -9.335 -218.460 -5.920 -218.290 ;
        RECT -5.615 -218.095 -3.215 -217.925 ;
        RECT -12.790 -219.680 -12.620 -218.725 ;
        RECT -21.235 -220.370 -17.595 -220.200 ;
        RECT -8.735 -220.200 -8.565 -218.640 ;
        RECT -8.245 -219.680 -8.075 -218.460 ;
        RECT -7.755 -220.200 -7.585 -218.640 ;
        RECT -7.155 -219.855 -6.985 -218.640 ;
        RECT -6.665 -219.680 -6.495 -218.460 ;
        RECT -6.175 -219.855 -6.005 -218.640 ;
        RECT -5.615 -219.855 -5.445 -218.095 ;
        RECT -7.155 -220.025 -5.445 -219.855 ;
        RECT -5.265 -218.465 -4.195 -218.295 ;
        RECT -5.265 -220.200 -5.095 -218.465 ;
        RECT -4.365 -219.680 -4.195 -218.465 ;
        RECT -3.385 -219.680 -3.215 -218.095 ;
        RECT -2.950 -218.110 -2.255 -217.840 ;
        RECT -1.860 -218.715 -1.645 -217.020 ;
        RECT -1.440 -217.340 -0.745 -217.070 ;
        RECT -0.310 -217.510 -0.095 -216.555 ;
        RECT 0.200 -216.650 0.370 -215.655 ;
        RECT 3.745 -215.670 3.940 -215.055 ;
        RECT 9.750 -215.225 12.910 -215.055 ;
        RECT 4.255 -215.425 9.295 -215.245 ;
        RECT 3.035 -216.455 3.265 -215.775 ;
        RECT -0.810 -217.740 -0.095 -217.510 ;
        RECT -1.835 -219.680 -1.665 -218.715 ;
        RECT -0.310 -218.725 -0.095 -217.740 ;
        RECT 0.125 -218.080 0.820 -217.810 ;
        RECT 3.065 -218.290 3.235 -216.455 ;
        RECT 3.765 -216.615 3.935 -215.670 ;
        RECT 3.755 -217.030 3.940 -216.615 ;
        RECT 4.255 -216.650 4.425 -215.425 ;
        RECT 5.835 -216.620 6.005 -215.610 ;
        RECT 6.325 -216.605 6.495 -215.610 ;
        RECT 7.645 -216.605 7.815 -215.610 ;
        RECT 5.820 -216.725 6.005 -216.620 ;
        RECT 5.225 -216.910 6.005 -216.725 ;
        RECT 6.315 -216.800 7.815 -216.605 ;
        RECT 5.225 -217.030 5.410 -216.910 ;
        RECT 3.755 -217.215 5.410 -217.030 ;
        RECT 8.135 -217.065 8.305 -215.610 ;
        RECT 9.115 -215.695 9.295 -215.425 ;
        RECT 9.115 -216.650 9.285 -215.695 ;
        RECT 9.605 -217.065 9.775 -215.610 ;
        RECT 10.665 -216.565 10.835 -215.610 ;
        RECT 11.130 -215.645 11.345 -215.225 ;
        RECT 10.640 -216.790 10.855 -216.565 ;
        RECT 11.155 -216.650 11.325 -215.645 ;
        RECT 12.210 -216.555 12.380 -215.610 ;
        RECT 12.675 -215.655 12.890 -215.225 ;
        RECT 10.160 -217.020 10.855 -216.790 ;
        RECT 5.670 -217.370 6.365 -217.100 ;
        RECT 6.970 -217.235 9.775 -217.065 ;
        RECT 6.970 -217.545 7.140 -217.235 ;
        RECT 3.760 -217.890 4.455 -217.620 ;
        RECT 6.410 -217.715 7.140 -217.545 ;
        RECT 6.410 -218.290 6.580 -217.715 ;
        RECT 7.505 -217.740 8.200 -217.470 ;
        RECT 3.065 -218.460 6.580 -218.290 ;
        RECT 6.885 -218.095 9.285 -217.925 ;
        RECT 3.065 -218.465 3.235 -218.460 ;
        RECT -0.290 -219.680 -0.120 -218.725 ;
        RECT -8.735 -220.370 -5.095 -220.200 ;
        RECT 3.765 -220.200 3.935 -218.640 ;
        RECT 4.255 -219.680 4.425 -218.460 ;
        RECT 4.745 -220.200 4.915 -218.640 ;
        RECT 5.345 -219.855 5.515 -218.640 ;
        RECT 5.835 -219.680 6.005 -218.460 ;
        RECT 6.325 -219.855 6.495 -218.640 ;
        RECT 6.885 -219.855 7.055 -218.095 ;
        RECT 5.345 -220.025 7.055 -219.855 ;
        RECT 7.235 -218.465 8.305 -218.295 ;
        RECT 7.235 -220.200 7.405 -218.465 ;
        RECT 8.135 -219.680 8.305 -218.465 ;
        RECT 9.115 -219.680 9.285 -218.095 ;
        RECT 9.550 -218.110 10.245 -217.840 ;
        RECT 10.640 -218.715 10.855 -217.020 ;
        RECT 11.060 -217.340 11.755 -217.070 ;
        RECT 12.190 -217.510 12.405 -216.555 ;
        RECT 12.700 -216.650 12.870 -215.655 ;
        RECT 16.245 -215.670 16.440 -215.055 ;
        RECT 22.250 -215.225 25.410 -215.055 ;
        RECT 16.755 -215.425 21.795 -215.245 ;
        RECT 15.120 -216.455 15.350 -215.775 ;
        RECT 15.145 -216.460 15.320 -216.455 ;
        RECT 11.690 -217.740 12.405 -217.510 ;
        RECT 10.665 -219.680 10.835 -218.715 ;
        RECT 12.190 -218.725 12.405 -217.740 ;
        RECT 12.625 -218.080 13.320 -217.810 ;
        RECT 15.145 -218.290 15.315 -216.460 ;
        RECT 16.265 -216.615 16.435 -215.670 ;
        RECT 16.255 -217.030 16.440 -216.615 ;
        RECT 16.755 -216.650 16.925 -215.425 ;
        RECT 18.335 -216.620 18.505 -215.610 ;
        RECT 18.825 -216.605 18.995 -215.610 ;
        RECT 20.145 -216.605 20.315 -215.610 ;
        RECT 18.320 -216.725 18.505 -216.620 ;
        RECT 17.725 -216.910 18.505 -216.725 ;
        RECT 18.815 -216.800 20.315 -216.605 ;
        RECT 17.725 -217.030 17.910 -216.910 ;
        RECT 16.255 -217.215 17.910 -217.030 ;
        RECT 20.635 -217.065 20.805 -215.610 ;
        RECT 21.615 -215.695 21.795 -215.425 ;
        RECT 21.615 -216.650 21.785 -215.695 ;
        RECT 22.105 -217.065 22.275 -215.610 ;
        RECT 23.165 -216.565 23.335 -215.610 ;
        RECT 23.630 -215.645 23.845 -215.225 ;
        RECT 23.140 -216.790 23.355 -216.565 ;
        RECT 23.655 -216.650 23.825 -215.645 ;
        RECT 24.710 -216.555 24.880 -215.610 ;
        RECT 25.175 -215.655 25.390 -215.225 ;
        RECT 22.660 -217.020 23.355 -216.790 ;
        RECT 19.470 -217.235 22.275 -217.065 ;
        RECT 19.470 -217.545 19.640 -217.235 ;
        RECT 16.260 -217.890 16.955 -217.620 ;
        RECT 18.910 -217.715 19.640 -217.545 ;
        RECT 18.910 -218.290 19.080 -217.715 ;
        RECT 20.005 -217.740 20.700 -217.470 ;
        RECT 15.145 -218.460 19.080 -218.290 ;
        RECT 19.385 -218.095 21.785 -217.925 ;
        RECT 12.210 -219.680 12.380 -218.725 ;
        RECT 3.765 -220.370 7.405 -220.200 ;
        RECT 16.265 -220.200 16.435 -218.640 ;
        RECT 16.755 -219.680 16.925 -218.460 ;
        RECT 17.245 -220.200 17.415 -218.640 ;
        RECT 17.845 -219.855 18.015 -218.640 ;
        RECT 18.335 -219.680 18.505 -218.460 ;
        RECT 18.825 -219.855 18.995 -218.640 ;
        RECT 19.385 -219.855 19.555 -218.095 ;
        RECT 17.845 -220.025 19.555 -219.855 ;
        RECT 19.735 -218.465 20.805 -218.295 ;
        RECT 19.735 -220.200 19.905 -218.465 ;
        RECT 20.635 -219.680 20.805 -218.465 ;
        RECT 21.615 -219.680 21.785 -218.095 ;
        RECT 22.050 -218.110 22.745 -217.840 ;
        RECT 23.140 -218.715 23.355 -217.020 ;
        RECT 24.690 -217.510 24.905 -216.555 ;
        RECT 25.200 -216.650 25.370 -215.655 ;
        RECT 31.245 -215.670 31.440 -215.055 ;
        RECT 31.755 -215.425 36.795 -215.245 ;
        RECT 37.170 -215.315 42.510 -215.055 ;
        RECT 44.840 -213.505 45.625 -213.305 ;
        RECT 29.645 -216.455 29.875 -215.775 ;
        RECT 24.190 -217.740 24.905 -217.510 ;
        RECT 23.165 -219.680 23.335 -218.715 ;
        RECT 24.690 -218.725 24.905 -217.740 ;
        RECT 25.125 -218.080 25.820 -217.810 ;
        RECT 29.675 -218.290 29.845 -216.455 ;
        RECT 31.265 -216.615 31.435 -215.670 ;
        RECT 31.255 -217.030 31.440 -216.615 ;
        RECT 31.755 -216.650 31.925 -215.425 ;
        RECT 33.335 -216.620 33.505 -215.610 ;
        RECT 33.825 -216.605 33.995 -215.610 ;
        RECT 35.145 -216.605 35.315 -215.610 ;
        RECT 33.320 -216.725 33.505 -216.620 ;
        RECT 32.725 -216.910 33.505 -216.725 ;
        RECT 33.815 -216.800 35.315 -216.605 ;
        RECT 32.725 -217.030 32.910 -216.910 ;
        RECT 31.255 -217.215 32.910 -217.030 ;
        RECT 35.635 -217.065 35.805 -215.610 ;
        RECT 36.615 -215.695 36.795 -215.425 ;
        RECT 36.615 -216.650 36.785 -215.695 ;
        RECT 37.105 -217.065 37.275 -215.610 ;
        RECT 38.165 -216.565 38.335 -215.610 ;
        RECT 38.630 -215.645 38.845 -215.315 ;
        RECT 38.140 -216.790 38.355 -216.565 ;
        RECT 38.655 -216.650 38.825 -215.645 ;
        RECT 39.710 -216.555 39.880 -215.610 ;
        RECT 40.175 -215.655 40.390 -215.315 ;
        RECT 37.660 -217.020 38.355 -216.790 ;
        RECT 34.470 -217.235 37.275 -217.065 ;
        RECT 34.470 -217.545 34.640 -217.235 ;
        RECT 31.260 -217.890 31.955 -217.620 ;
        RECT 33.910 -217.715 34.640 -217.545 ;
        RECT 33.910 -218.290 34.080 -217.715 ;
        RECT 35.005 -217.740 35.700 -217.470 ;
        RECT 29.675 -218.460 34.080 -218.290 ;
        RECT 34.385 -218.095 36.785 -217.925 ;
        RECT 24.710 -219.680 24.880 -218.725 ;
        RECT 16.265 -220.370 19.905 -220.200 ;
        RECT 31.265 -220.200 31.435 -218.640 ;
        RECT 31.755 -219.680 31.925 -218.460 ;
        RECT 32.245 -220.200 32.415 -218.640 ;
        RECT 32.845 -219.855 33.015 -218.640 ;
        RECT 33.335 -219.680 33.505 -218.460 ;
        RECT 33.825 -219.855 33.995 -218.640 ;
        RECT 34.385 -219.855 34.555 -218.095 ;
        RECT 32.845 -220.025 34.555 -219.855 ;
        RECT 34.735 -218.465 35.805 -218.295 ;
        RECT 34.735 -220.200 34.905 -218.465 ;
        RECT 35.635 -219.680 35.805 -218.465 ;
        RECT 36.615 -219.680 36.785 -218.095 ;
        RECT 37.050 -218.110 37.745 -217.840 ;
        RECT 38.140 -218.715 38.355 -217.020 ;
        RECT 39.690 -217.510 39.905 -216.555 ;
        RECT 40.200 -216.650 40.370 -215.655 ;
        RECT 39.190 -217.740 39.905 -217.510 ;
        RECT 38.165 -219.680 38.335 -218.715 ;
        RECT 39.690 -218.725 39.905 -217.740 ;
        RECT 40.125 -218.080 40.820 -217.810 ;
        RECT 39.710 -219.680 39.880 -218.725 ;
        RECT 31.265 -220.370 34.905 -220.200 ;
        RECT -36.555 -220.700 -35.740 -220.600 ;
        RECT -131.940 -221.800 -117.710 -220.870 ;
        RECT -95.030 -221.380 -35.740 -220.700 ;
        RECT 44.840 -221.160 45.110 -213.505 ;
        RECT 45.910 -215.025 46.180 -212.870 ;
        RECT 45.415 -215.295 46.180 -215.025 ;
        RECT 45.415 -221.160 45.685 -215.295 ;
        RECT 46.135 -220.685 46.405 -220.535 ;
        RECT 46.625 -220.685 46.895 -212.195 ;
        RECT 49.220 -218.880 50.525 -209.980 ;
        RECT 64.300 -211.140 67.440 -210.970 ;
        RECT 56.840 -211.255 57.010 -211.235 ;
        RECT 56.810 -212.520 57.040 -211.255 ;
        RECT 57.820 -212.195 57.990 -211.235 ;
        RECT 58.800 -212.195 58.970 -211.235 ;
        RECT 61.250 -211.255 61.420 -211.235 ;
        RECT 60.145 -212.165 60.430 -211.345 ;
        RECT 57.790 -212.520 58.020 -212.195 ;
        RECT 58.770 -212.520 59.000 -212.195 ;
        RECT 56.810 -212.560 59.000 -212.520 ;
        RECT 61.220 -212.520 61.450 -211.255 ;
        RECT 62.230 -212.195 62.400 -211.235 ;
        RECT 63.210 -212.195 63.380 -211.235 ;
        RECT 64.300 -211.365 64.480 -211.140 ;
        RECT 62.200 -212.520 62.430 -212.195 ;
        RECT 63.180 -212.520 63.410 -212.195 ;
        RECT 61.220 -212.560 63.410 -212.520 ;
        RECT 63.685 -212.440 64.055 -211.600 ;
        RECT 64.305 -211.735 64.475 -211.365 ;
        RECT 63.685 -212.560 64.050 -212.440 ;
        RECT 56.810 -212.670 59.150 -212.560 ;
        RECT 60.200 -212.650 61.040 -212.595 ;
        RECT 59.440 -212.670 59.740 -212.650 ;
        RECT 60.025 -212.670 61.040 -212.650 ;
        RECT 56.810 -212.750 61.040 -212.670 ;
        RECT 56.350 -213.930 56.520 -213.135 ;
        RECT 56.810 -213.215 57.040 -212.750 ;
        RECT 56.840 -213.675 57.010 -213.215 ;
        RECT 57.330 -213.930 57.500 -213.135 ;
        RECT 57.790 -213.215 58.020 -212.750 ;
        RECT 58.770 -212.880 61.040 -212.750 ;
        RECT 58.770 -212.910 59.150 -212.880 ;
        RECT 57.820 -213.675 57.990 -213.215 ;
        RECT 58.310 -213.930 58.480 -213.135 ;
        RECT 58.770 -213.215 59.000 -212.910 ;
        RECT 58.800 -213.675 58.970 -213.215 ;
        RECT 59.440 -213.310 59.740 -212.880 ;
        RECT 60.025 -212.940 61.040 -212.880 ;
        RECT 60.200 -212.965 61.040 -212.940 ;
        RECT 61.220 -212.750 64.050 -212.560 ;
        RECT 60.760 -213.930 60.930 -213.135 ;
        RECT 61.220 -213.215 61.450 -212.750 ;
        RECT 61.250 -213.675 61.420 -213.215 ;
        RECT 61.740 -213.930 61.910 -213.135 ;
        RECT 62.200 -213.215 62.430 -212.750 ;
        RECT 63.180 -212.910 64.050 -212.750 ;
        RECT 64.275 -212.470 64.510 -211.735 ;
        RECT 64.795 -211.770 64.965 -211.310 ;
        RECT 65.280 -211.415 65.490 -211.140 ;
        RECT 64.790 -212.030 64.970 -211.770 ;
        RECT 65.285 -211.850 65.455 -211.415 ;
        RECT 65.775 -211.760 65.945 -211.310 ;
        RECT 66.250 -211.420 66.460 -211.140 ;
        RECT 65.775 -211.850 65.960 -211.760 ;
        RECT 66.265 -211.850 66.435 -211.420 ;
        RECT 66.755 -211.760 66.925 -211.310 ;
        RECT 67.230 -211.395 67.440 -211.140 ;
        RECT 77.800 -211.140 80.940 -210.970 ;
        RECT 69.965 -211.255 70.135 -211.235 ;
        RECT 65.780 -212.030 65.960 -211.850 ;
        RECT 66.750 -212.030 66.930 -211.760 ;
        RECT 67.245 -211.850 67.415 -211.395 ;
        RECT 67.735 -211.810 67.905 -211.310 ;
        RECT 67.720 -212.030 67.930 -211.810 ;
        RECT 64.790 -212.200 67.930 -212.030 ;
        RECT 64.275 -212.840 65.135 -212.470 ;
        RECT 67.055 -212.640 67.930 -212.200 ;
        RECT 69.935 -212.520 70.165 -211.255 ;
        RECT 70.945 -212.195 71.115 -211.235 ;
        RECT 71.925 -212.195 72.095 -211.235 ;
        RECT 74.750 -211.255 74.920 -211.235 ;
        RECT 73.645 -211.735 73.930 -211.345 ;
        RECT 72.625 -211.960 73.930 -211.735 ;
        RECT 70.915 -212.520 71.145 -212.195 ;
        RECT 71.895 -212.520 72.125 -212.195 ;
        RECT 69.935 -212.560 72.125 -212.520 ;
        RECT 68.915 -212.640 69.755 -212.595 ;
        RECT 62.230 -213.675 62.400 -213.215 ;
        RECT 62.720 -213.930 62.890 -213.135 ;
        RECT 63.180 -213.215 63.410 -212.910 ;
        RECT 63.210 -213.675 63.380 -213.215 ;
        RECT 64.275 -213.515 64.510 -212.840 ;
        RECT 67.055 -212.925 69.755 -212.640 ;
        RECT 67.055 -213.035 67.930 -212.925 ;
        RECT 68.915 -212.965 69.755 -212.925 ;
        RECT 69.935 -212.630 72.275 -212.560 ;
        RECT 72.625 -212.630 72.850 -211.960 ;
        RECT 73.645 -212.165 73.930 -211.960 ;
        RECT 69.935 -212.750 72.850 -212.630 ;
        RECT 64.775 -213.205 67.930 -213.035 ;
        RECT 64.775 -213.410 64.980 -213.205 ;
        RECT 64.305 -213.865 64.475 -213.515 ;
        RECT 56.305 -214.270 63.385 -213.930 ;
        RECT 64.280 -214.155 64.500 -213.865 ;
        RECT 64.795 -213.925 64.965 -213.410 ;
        RECT 65.285 -213.810 65.455 -213.385 ;
        RECT 65.765 -213.450 65.970 -213.205 ;
        RECT 65.260 -214.155 65.480 -213.810 ;
        RECT 65.775 -213.925 65.945 -213.450 ;
        RECT 66.265 -213.810 66.435 -213.385 ;
        RECT 66.735 -213.450 66.940 -213.205 ;
        RECT 67.720 -213.240 67.930 -213.205 ;
        RECT 66.240 -214.155 66.460 -213.810 ;
        RECT 66.755 -213.925 66.925 -213.450 ;
        RECT 67.245 -213.865 67.415 -213.385 ;
        RECT 67.720 -213.405 67.925 -213.240 ;
        RECT 67.690 -213.455 67.925 -213.405 ;
        RECT 67.225 -214.155 67.445 -213.865 ;
        RECT 67.690 -214.065 67.920 -213.455 ;
        RECT 69.475 -213.930 69.645 -213.135 ;
        RECT 69.935 -213.215 70.165 -212.750 ;
        RECT 69.965 -213.675 70.135 -213.215 ;
        RECT 70.455 -213.930 70.625 -213.135 ;
        RECT 70.915 -213.215 71.145 -212.750 ;
        RECT 71.895 -212.855 72.850 -212.750 ;
        RECT 74.720 -212.520 74.950 -211.255 ;
        RECT 75.730 -212.195 75.900 -211.235 ;
        RECT 76.710 -212.195 76.880 -211.235 ;
        RECT 77.800 -211.365 77.980 -211.140 ;
        RECT 75.700 -212.520 75.930 -212.195 ;
        RECT 76.680 -212.520 76.910 -212.195 ;
        RECT 74.720 -212.560 76.910 -212.520 ;
        RECT 77.185 -212.440 77.555 -211.600 ;
        RECT 77.805 -211.735 77.975 -211.365 ;
        RECT 77.185 -212.560 77.550 -212.440 ;
        RECT 74.720 -212.750 77.550 -212.560 ;
        RECT 71.895 -212.910 72.275 -212.855 ;
        RECT 70.945 -213.675 71.115 -213.215 ;
        RECT 71.435 -213.930 71.605 -213.135 ;
        RECT 71.895 -213.215 72.125 -212.910 ;
        RECT 71.925 -213.675 72.095 -213.215 ;
        RECT 72.525 -213.430 72.825 -212.855 ;
        RECT 74.260 -213.930 74.430 -213.135 ;
        RECT 74.720 -213.215 74.950 -212.750 ;
        RECT 74.750 -213.675 74.920 -213.215 ;
        RECT 75.240 -213.930 75.410 -213.135 ;
        RECT 75.700 -213.215 75.930 -212.750 ;
        RECT 76.680 -212.910 77.550 -212.750 ;
        RECT 77.775 -212.470 78.010 -211.735 ;
        RECT 78.295 -211.770 78.465 -211.310 ;
        RECT 78.780 -211.415 78.990 -211.140 ;
        RECT 78.290 -212.030 78.470 -211.770 ;
        RECT 78.785 -211.850 78.955 -211.415 ;
        RECT 79.275 -211.760 79.445 -211.310 ;
        RECT 79.750 -211.420 79.960 -211.140 ;
        RECT 79.275 -211.850 79.460 -211.760 ;
        RECT 79.765 -211.850 79.935 -211.420 ;
        RECT 80.255 -211.760 80.425 -211.310 ;
        RECT 80.730 -211.395 80.940 -211.140 ;
        RECT 83.465 -211.255 83.635 -211.235 ;
        RECT 79.280 -212.030 79.460 -211.850 ;
        RECT 80.250 -212.030 80.430 -211.760 ;
        RECT 80.745 -211.850 80.915 -211.395 ;
        RECT 81.235 -211.810 81.405 -211.310 ;
        RECT 81.220 -212.030 81.430 -211.810 ;
        RECT 78.290 -212.200 81.430 -212.030 ;
        RECT 77.775 -212.840 78.635 -212.470 ;
        RECT 80.555 -212.625 81.430 -212.200 ;
        RECT 83.435 -212.520 83.665 -211.255 ;
        RECT 84.445 -212.195 84.615 -211.235 ;
        RECT 85.425 -212.195 85.595 -211.235 ;
        RECT 84.415 -212.520 84.645 -212.195 ;
        RECT 85.395 -212.520 85.625 -212.195 ;
        RECT 83.435 -212.560 85.625 -212.520 ;
        RECT 82.415 -212.625 83.255 -212.595 ;
        RECT 75.730 -213.675 75.900 -213.215 ;
        RECT 76.220 -213.930 76.390 -213.135 ;
        RECT 76.680 -213.215 76.910 -212.910 ;
        RECT 76.710 -213.675 76.880 -213.215 ;
        RECT 77.775 -213.515 78.010 -212.840 ;
        RECT 80.555 -212.890 83.255 -212.625 ;
        RECT 80.555 -213.035 81.430 -212.890 ;
        RECT 82.415 -212.965 83.255 -212.890 ;
        RECT 83.435 -212.605 85.775 -212.560 ;
        RECT 83.435 -212.615 86.185 -212.605 ;
        RECT 83.435 -212.750 86.190 -212.615 ;
        RECT 78.275 -213.205 81.430 -213.035 ;
        RECT 78.275 -213.410 78.480 -213.205 ;
        RECT 77.805 -213.865 77.975 -213.515 ;
        RECT 64.280 -214.325 67.445 -214.155 ;
        RECT 69.430 -214.270 76.885 -213.930 ;
        RECT 77.780 -214.155 78.000 -213.865 ;
        RECT 78.295 -213.925 78.465 -213.410 ;
        RECT 78.785 -213.810 78.955 -213.385 ;
        RECT 79.265 -213.450 79.470 -213.205 ;
        RECT 78.760 -214.155 78.980 -213.810 ;
        RECT 79.275 -213.925 79.445 -213.450 ;
        RECT 79.765 -213.810 79.935 -213.385 ;
        RECT 80.235 -213.450 80.440 -213.205 ;
        RECT 81.220 -213.240 81.430 -213.205 ;
        RECT 79.740 -214.155 79.960 -213.810 ;
        RECT 80.255 -213.925 80.425 -213.450 ;
        RECT 80.745 -213.865 80.915 -213.385 ;
        RECT 81.220 -213.455 81.425 -213.240 ;
        RECT 80.725 -214.155 80.945 -213.865 ;
        RECT 81.235 -213.925 81.405 -213.455 ;
        RECT 82.975 -213.930 83.145 -213.135 ;
        RECT 83.435 -213.215 83.665 -212.750 ;
        RECT 83.465 -213.675 83.635 -213.215 ;
        RECT 83.955 -213.930 84.125 -213.135 ;
        RECT 84.415 -213.215 84.645 -212.750 ;
        RECT 85.395 -212.800 86.190 -212.750 ;
        RECT 85.395 -212.910 85.775 -212.800 ;
        RECT 84.445 -213.675 84.615 -213.215 ;
        RECT 84.935 -213.930 85.105 -213.135 ;
        RECT 85.395 -213.215 85.625 -212.910 ;
        RECT 85.425 -213.675 85.595 -213.215 ;
        RECT 77.780 -214.325 80.945 -214.155 ;
        RECT 82.930 -214.270 85.600 -213.930 ;
        RECT 59.235 -214.505 59.895 -214.450 ;
        RECT 81.850 -214.505 82.510 -214.440 ;
        RECT 59.235 -214.700 84.540 -214.505 ;
        RECT 85.950 -214.590 86.190 -212.800 ;
        RECT 59.235 -214.750 59.895 -214.700 ;
        RECT 81.850 -214.740 82.510 -214.700 ;
        RECT 85.895 -215.275 86.195 -214.590 ;
        RECT 57.620 -215.395 58.280 -215.300 ;
        RECT 70.785 -215.395 71.470 -215.300 ;
        RECT 83.770 -215.395 84.455 -215.330 ;
        RECT 57.615 -215.590 84.540 -215.395 ;
        RECT 57.620 -215.600 59.445 -215.590 ;
        RECT 58.140 -218.880 59.445 -215.600 ;
        RECT 61.225 -215.945 64.390 -215.775 ;
        RECT 66.410 -215.830 66.965 -215.590 ;
        RECT 70.785 -215.600 71.470 -215.590 ;
        RECT 67.840 -215.830 70.440 -215.820 ;
        RECT 70.800 -215.830 71.355 -215.600 ;
        RECT 60.765 -216.645 60.935 -216.175 ;
        RECT 61.225 -216.235 61.445 -215.945 ;
        RECT 60.745 -216.860 60.950 -216.645 ;
        RECT 61.255 -216.715 61.425 -216.235 ;
        RECT 61.745 -216.650 61.915 -216.175 ;
        RECT 62.210 -216.290 62.430 -215.945 ;
        RECT 60.740 -216.895 60.950 -216.860 ;
        RECT 61.730 -216.895 61.935 -216.650 ;
        RECT 62.235 -216.715 62.405 -216.290 ;
        RECT 62.725 -216.650 62.895 -216.175 ;
        RECT 63.190 -216.290 63.410 -215.945 ;
        RECT 62.700 -216.895 62.905 -216.650 ;
        RECT 63.215 -216.715 63.385 -216.290 ;
        RECT 63.705 -216.690 63.875 -216.175 ;
        RECT 64.170 -216.235 64.390 -215.945 ;
        RECT 65.285 -216.160 72.140 -215.830 ;
        RECT 65.285 -216.170 67.955 -216.160 ;
        RECT 69.470 -216.170 72.140 -216.160 ;
        RECT 74.725 -215.945 77.890 -215.775 ;
        RECT 79.790 -215.830 80.345 -215.590 ;
        RECT 83.770 -215.630 84.455 -215.590 ;
        RECT 83.845 -215.830 84.400 -215.630 ;
        RECT 64.195 -216.585 64.365 -216.235 ;
        RECT 63.690 -216.895 63.895 -216.690 ;
        RECT 60.740 -217.055 63.895 -216.895 ;
        RECT 60.365 -217.065 63.895 -217.055 ;
        RECT 60.365 -217.355 61.615 -217.065 ;
        RECT 64.160 -217.260 64.395 -216.585 ;
        RECT 65.290 -216.885 65.460 -216.425 ;
        RECT 65.260 -217.190 65.490 -216.885 ;
        RECT 65.780 -216.965 65.950 -216.170 ;
        RECT 66.270 -216.885 66.440 -216.425 ;
        RECT 60.740 -217.900 61.615 -217.355 ;
        RECT 63.535 -217.630 64.395 -217.260 ;
        RECT 60.740 -218.070 63.880 -217.900 ;
        RECT 60.740 -218.290 60.950 -218.070 ;
        RECT 60.765 -218.790 60.935 -218.290 ;
        RECT 61.255 -218.705 61.425 -218.250 ;
        RECT 61.740 -218.340 61.920 -218.070 ;
        RECT 62.710 -218.250 62.890 -218.070 ;
        RECT 49.220 -220.185 59.445 -218.880 ;
        RECT 61.230 -218.960 61.440 -218.705 ;
        RECT 61.745 -218.790 61.915 -218.340 ;
        RECT 62.235 -218.680 62.405 -218.250 ;
        RECT 62.710 -218.340 62.895 -218.250 ;
        RECT 62.210 -218.960 62.420 -218.680 ;
        RECT 62.725 -218.790 62.895 -218.340 ;
        RECT 63.215 -218.685 63.385 -218.250 ;
        RECT 63.700 -218.330 63.880 -218.070 ;
        RECT 63.180 -218.960 63.390 -218.685 ;
        RECT 63.705 -218.790 63.875 -218.330 ;
        RECT 64.160 -218.365 64.395 -217.630 ;
        RECT 64.620 -217.350 65.490 -217.190 ;
        RECT 66.240 -217.350 66.470 -216.885 ;
        RECT 66.760 -216.965 66.930 -216.170 ;
        RECT 67.250 -216.885 67.420 -216.425 ;
        RECT 67.220 -217.350 67.450 -216.885 ;
        RECT 67.740 -216.965 67.910 -216.170 ;
        RECT 69.475 -216.885 69.645 -216.425 ;
        RECT 69.445 -217.190 69.675 -216.885 ;
        RECT 69.965 -216.965 70.135 -216.170 ;
        RECT 70.455 -216.885 70.625 -216.425 ;
        RECT 64.620 -217.540 67.450 -217.350 ;
        RECT 64.620 -217.660 64.985 -217.540 ;
        RECT 64.195 -218.735 64.365 -218.365 ;
        RECT 64.615 -218.500 64.985 -217.660 ;
        RECT 65.260 -217.580 67.450 -217.540 ;
        RECT 65.260 -217.905 65.490 -217.580 ;
        RECT 66.240 -217.905 66.470 -217.580 ;
        RECT 64.190 -218.960 64.370 -218.735 ;
        RECT 65.290 -218.865 65.460 -217.905 ;
        RECT 66.270 -218.865 66.440 -217.905 ;
        RECT 67.220 -218.845 67.450 -217.580 ;
        RECT 68.955 -217.350 69.675 -217.190 ;
        RECT 70.425 -217.350 70.655 -216.885 ;
        RECT 70.945 -216.965 71.115 -216.170 ;
        RECT 71.435 -216.885 71.605 -216.425 ;
        RECT 71.405 -217.350 71.635 -216.885 ;
        RECT 71.925 -216.965 72.095 -216.170 ;
        RECT 74.265 -216.645 74.435 -216.175 ;
        RECT 74.725 -216.235 74.945 -215.945 ;
        RECT 74.245 -216.860 74.450 -216.645 ;
        RECT 74.755 -216.715 74.925 -216.235 ;
        RECT 75.245 -216.650 75.415 -216.175 ;
        RECT 75.710 -216.290 75.930 -215.945 ;
        RECT 74.240 -216.895 74.450 -216.860 ;
        RECT 75.230 -216.895 75.435 -216.650 ;
        RECT 75.735 -216.715 75.905 -216.290 ;
        RECT 76.225 -216.650 76.395 -216.175 ;
        RECT 76.690 -216.290 76.910 -215.945 ;
        RECT 76.200 -216.895 76.405 -216.650 ;
        RECT 76.715 -216.715 76.885 -216.290 ;
        RECT 77.205 -216.690 77.375 -216.175 ;
        RECT 77.670 -216.235 77.890 -215.945 ;
        RECT 78.785 -216.170 85.640 -215.830 ;
        RECT 77.695 -216.585 77.865 -216.235 ;
        RECT 77.190 -216.895 77.395 -216.690 ;
        RECT 74.240 -217.065 77.395 -216.895 ;
        RECT 68.955 -217.540 71.635 -217.350 ;
        RECT 71.815 -217.170 72.655 -217.135 ;
        RECT 71.815 -217.470 72.765 -217.170 ;
        RECT 73.785 -217.365 75.115 -217.065 ;
        RECT 77.660 -217.260 77.895 -216.585 ;
        RECT 78.790 -216.885 78.960 -216.425 ;
        RECT 78.760 -217.190 78.990 -216.885 ;
        RECT 79.280 -216.965 79.450 -216.170 ;
        RECT 79.770 -216.885 79.940 -216.425 ;
        RECT 71.815 -217.505 72.655 -217.470 ;
        RECT 68.240 -218.185 68.525 -217.935 ;
        RECT 68.955 -218.185 69.265 -217.540 ;
        RECT 69.445 -217.580 71.635 -217.540 ;
        RECT 69.445 -217.905 69.675 -217.580 ;
        RECT 70.425 -217.905 70.655 -217.580 ;
        RECT 68.240 -218.495 69.265 -218.185 ;
        RECT 68.240 -218.755 68.525 -218.495 ;
        RECT 67.250 -218.865 67.420 -218.845 ;
        RECT 69.475 -218.865 69.645 -217.905 ;
        RECT 70.455 -218.865 70.625 -217.905 ;
        RECT 71.405 -218.845 71.635 -217.580 ;
        RECT 74.240 -217.900 75.115 -217.365 ;
        RECT 77.035 -217.630 77.895 -217.260 ;
        RECT 74.240 -218.070 77.380 -217.900 ;
        RECT 74.240 -218.290 74.450 -218.070 ;
        RECT 74.265 -218.790 74.435 -218.290 ;
        RECT 74.755 -218.705 74.925 -218.250 ;
        RECT 75.240 -218.340 75.420 -218.070 ;
        RECT 76.210 -218.250 76.390 -218.070 ;
        RECT 71.435 -218.865 71.605 -218.845 ;
        RECT 61.230 -219.130 64.370 -218.960 ;
        RECT 74.730 -218.960 74.940 -218.705 ;
        RECT 75.245 -218.790 75.415 -218.340 ;
        RECT 75.735 -218.680 75.905 -218.250 ;
        RECT 76.210 -218.340 76.395 -218.250 ;
        RECT 75.710 -218.960 75.920 -218.680 ;
        RECT 76.225 -218.790 76.395 -218.340 ;
        RECT 76.715 -218.685 76.885 -218.250 ;
        RECT 77.200 -218.330 77.380 -218.070 ;
        RECT 76.680 -218.960 76.890 -218.685 ;
        RECT 77.205 -218.790 77.375 -218.330 ;
        RECT 77.660 -218.365 77.895 -217.630 ;
        RECT 78.120 -217.350 78.990 -217.190 ;
        RECT 79.740 -217.350 79.970 -216.885 ;
        RECT 80.260 -216.965 80.430 -216.170 ;
        RECT 80.750 -216.885 80.920 -216.425 ;
        RECT 80.720 -217.350 80.950 -216.885 ;
        RECT 81.240 -216.965 81.410 -216.170 ;
        RECT 82.030 -217.135 82.330 -216.415 ;
        RECT 82.975 -216.885 83.145 -216.425 ;
        RECT 78.120 -217.540 80.950 -217.350 ;
        RECT 81.130 -217.445 82.330 -217.135 ;
        RECT 82.945 -217.190 83.175 -216.885 ;
        RECT 83.465 -216.965 83.635 -216.170 ;
        RECT 83.955 -216.885 84.125 -216.425 ;
        RECT 82.510 -217.350 83.175 -217.190 ;
        RECT 83.925 -217.350 84.155 -216.885 ;
        RECT 84.445 -216.965 84.615 -216.170 ;
        RECT 84.935 -216.885 85.105 -216.425 ;
        RECT 84.905 -217.350 85.135 -216.885 ;
        RECT 85.425 -216.965 85.595 -216.170 ;
        RECT 85.950 -217.135 86.190 -215.275 ;
        RECT 81.130 -217.450 82.145 -217.445 ;
        RECT 81.130 -217.505 81.970 -217.450 ;
        RECT 78.120 -217.660 78.485 -217.540 ;
        RECT 77.695 -218.735 77.865 -218.365 ;
        RECT 78.115 -218.500 78.485 -217.660 ;
        RECT 78.760 -217.580 80.950 -217.540 ;
        RECT 78.760 -217.905 78.990 -217.580 ;
        RECT 79.740 -217.905 79.970 -217.580 ;
        RECT 77.690 -218.960 77.870 -218.735 ;
        RECT 78.790 -218.865 78.960 -217.905 ;
        RECT 79.770 -218.865 79.940 -217.905 ;
        RECT 80.720 -218.845 80.950 -217.580 ;
        RECT 82.510 -217.540 85.135 -217.350 ;
        RECT 85.315 -217.355 86.190 -217.135 ;
        RECT 85.315 -217.505 86.155 -217.355 ;
        RECT 81.740 -218.190 82.025 -217.935 ;
        RECT 82.510 -218.190 82.740 -217.540 ;
        RECT 82.945 -217.580 85.135 -217.540 ;
        RECT 82.945 -217.905 83.175 -217.580 ;
        RECT 83.925 -217.905 84.155 -217.580 ;
        RECT 81.740 -218.435 82.740 -218.190 ;
        RECT 81.740 -218.755 82.025 -218.435 ;
        RECT 80.750 -218.865 80.920 -218.845 ;
        RECT 82.975 -218.865 83.145 -217.905 ;
        RECT 83.955 -218.865 84.125 -217.905 ;
        RECT 84.905 -218.845 85.135 -217.580 ;
        RECT 132.935 -218.640 133.665 -199.890 ;
        RECT 136.915 -200.730 137.295 -199.890 ;
        RECT 136.915 -201.110 137.625 -200.730 ;
        RECT 137.245 -203.055 137.625 -201.110 ;
        RECT 142.290 -200.940 145.615 -200.800 ;
        RECT 142.290 -201.230 147.465 -200.940 ;
        RECT 151.335 -201.225 151.795 -200.800 ;
        RECT 142.290 -201.635 142.720 -201.230 ;
        RECT 143.590 -201.415 143.765 -201.230 ;
        RECT 145.215 -201.245 147.465 -201.230 ;
        RECT 138.030 -202.065 142.720 -201.635 ;
        RECT 137.245 -203.515 137.920 -203.055 ;
        RECT 138.730 -203.345 138.900 -202.065 ;
        RECT 139.220 -203.345 139.390 -202.305 ;
        RECT 139.710 -203.345 139.880 -202.065 ;
        RECT 140.200 -203.175 140.370 -202.305 ;
        RECT 143.105 -202.955 143.275 -201.415 ;
        RECT 143.595 -202.955 143.765 -201.415 ;
        RECT 144.085 -202.955 144.255 -201.415 ;
        RECT 144.575 -202.955 144.745 -201.415 ;
        RECT 145.065 -202.955 145.235 -201.415 ;
        RECT 142.945 -203.170 143.300 -203.165 ;
        RECT 145.005 -203.170 145.375 -203.140 ;
        RECT 142.945 -203.175 145.375 -203.170 ;
        RECT 140.200 -203.345 145.375 -203.175 ;
        RECT 147.160 -203.280 147.465 -201.245 ;
        RECT 140.205 -203.365 145.375 -203.345 ;
        RECT 140.205 -203.375 142.950 -203.365 ;
        RECT 138.140 -203.515 138.505 -203.485 ;
        RECT 145.005 -203.495 145.375 -203.365 ;
        RECT 137.245 -203.600 138.505 -203.515 ;
        RECT 137.270 -203.720 138.505 -203.600 ;
        RECT 142.680 -203.655 143.355 -203.615 ;
        RECT 142.580 -203.665 143.355 -203.655 ;
        RECT 137.270 -203.805 137.920 -203.720 ;
        RECT 138.140 -203.785 138.505 -203.720 ;
        RECT 141.545 -203.845 143.355 -203.665 ;
        RECT 145.940 -203.710 149.865 -203.280 ;
        RECT 142.580 -203.855 143.355 -203.845 ;
        RECT 142.680 -203.885 143.355 -203.855 ;
        RECT 143.595 -203.770 145.690 -203.730 ;
        RECT 143.595 -203.920 145.745 -203.770 ;
        RECT 138.730 -204.995 138.900 -203.955 ;
        RECT 139.710 -204.995 139.880 -203.955 ;
        RECT 140.690 -204.995 140.860 -203.955 ;
        RECT 143.595 -205.640 143.765 -203.920 ;
        RECT 144.575 -205.640 144.745 -203.920 ;
        RECT 145.440 -204.665 145.745 -203.920 ;
        RECT 146.640 -204.490 146.810 -203.710 ;
        RECT 147.130 -204.490 147.300 -203.950 ;
        RECT 147.620 -204.490 147.790 -203.710 ;
        RECT 148.110 -204.490 148.280 -203.950 ;
        RECT 146.050 -204.665 146.415 -204.635 ;
        RECT 145.440 -204.730 146.415 -204.665 ;
        RECT 145.550 -204.870 146.415 -204.730 ;
        RECT 146.050 -204.935 146.415 -204.870 ;
        RECT 148.600 -204.785 150.460 -204.435 ;
        RECT 146.640 -205.645 146.810 -205.105 ;
        RECT 147.620 -205.645 147.790 -205.105 ;
        RECT 148.600 -205.645 148.770 -204.785 ;
        RECT 146.870 -207.985 148.070 -207.815 ;
        RECT 138.600 -210.320 138.770 -208.600 ;
        RECT 139.580 -210.320 139.750 -208.600 ;
        RECT 141.645 -209.135 141.815 -208.595 ;
        RECT 142.625 -209.135 142.795 -208.595 ;
        RECT 141.055 -209.370 141.420 -209.305 ;
        RECT 140.555 -209.510 141.420 -209.370 ;
        RECT 140.445 -209.575 141.420 -209.510 ;
        RECT 140.445 -210.320 140.750 -209.575 ;
        RECT 141.055 -209.605 141.420 -209.575 ;
        RECT 143.605 -209.455 143.775 -208.595 ;
        RECT 138.600 -210.470 140.750 -210.320 ;
        RECT 138.600 -210.510 140.695 -210.470 ;
        RECT 141.645 -210.530 141.815 -209.750 ;
        RECT 142.135 -210.290 142.305 -209.750 ;
        RECT 142.625 -210.530 142.795 -209.750 ;
        RECT 143.115 -210.290 143.285 -209.750 ;
        RECT 143.605 -209.805 144.995 -209.455 ;
        RECT 136.820 -210.875 137.955 -210.865 ;
        RECT 140.010 -210.875 140.380 -210.745 ;
        RECT 136.820 -211.065 140.380 -210.875 ;
        RECT 140.945 -210.960 144.020 -210.530 ;
        RECT 137.950 -211.070 140.380 -211.065 ;
        RECT 137.950 -211.075 138.305 -211.070 ;
        RECT 140.010 -211.100 140.380 -211.070 ;
        RECT 138.110 -212.825 138.280 -211.285 ;
        RECT 138.600 -212.825 138.770 -211.285 ;
        RECT 139.090 -212.825 139.260 -211.285 ;
        RECT 139.580 -212.825 139.750 -211.285 ;
        RECT 140.070 -212.825 140.240 -211.285 ;
        RECT 138.595 -213.085 138.770 -212.825 ;
        RECT 142.165 -212.995 142.470 -210.960 ;
        RECT 144.615 -211.780 144.965 -209.805 ;
        RECT 145.835 -211.075 146.005 -208.155 ;
        RECT 146.870 -208.195 147.080 -207.985 ;
        RECT 145.815 -211.370 146.025 -211.075 ;
        RECT 146.890 -211.105 147.060 -208.195 ;
        RECT 147.380 -211.095 147.550 -208.155 ;
        RECT 147.860 -208.205 148.070 -207.985 ;
        RECT 146.875 -211.370 147.085 -211.105 ;
        RECT 145.815 -211.550 147.085 -211.370 ;
        RECT 147.360 -211.365 147.570 -211.095 ;
        RECT 147.870 -211.195 148.040 -208.205 ;
        RECT 148.930 -211.125 149.100 -208.155 ;
        RECT 147.360 -211.560 148.065 -211.365 ;
        RECT 147.850 -211.620 148.065 -211.560 ;
        RECT 146.640 -211.780 147.415 -211.730 ;
        RECT 144.615 -211.960 147.415 -211.780 ;
        RECT 144.615 -211.970 144.965 -211.960 ;
        RECT 146.640 -212.005 147.415 -211.960 ;
        RECT 147.850 -211.895 148.755 -211.620 ;
        RECT 147.850 -212.245 148.065 -211.895 ;
        RECT 145.290 -212.315 146.065 -212.270 ;
        RECT 145.105 -212.485 146.065 -212.315 ;
        RECT 145.290 -212.545 146.065 -212.485 ;
        RECT 146.295 -212.445 148.065 -212.245 ;
        RECT 148.925 -212.345 149.140 -211.125 ;
        RECT 150.110 -211.470 150.460 -204.785 ;
        RECT 151.450 -211.100 151.665 -201.225 ;
        RECT 153.085 -203.340 153.465 -199.820 ;
        RECT 154.595 -199.600 163.530 -199.410 ;
        RECT 175.835 -198.835 179.495 -198.105 ;
        RECT 184.405 -197.565 184.710 -196.090 ;
        RECT 188.075 -196.975 188.245 -195.505 ;
        RECT 188.535 -195.585 188.760 -195.235 ;
        RECT 190.495 -195.335 195.115 -195.135 ;
        RECT 190.735 -195.350 195.115 -195.335 ;
        RECT 188.040 -197.565 188.275 -196.975 ;
        RECT 188.565 -197.045 188.735 -195.585 ;
        RECT 189.055 -196.970 189.225 -195.505 ;
        RECT 190.265 -196.920 190.435 -195.505 ;
        RECT 190.735 -195.550 190.955 -195.350 ;
        RECT 196.105 -195.460 196.500 -195.110 ;
        RECT 189.020 -197.565 189.255 -196.970 ;
        RECT 190.230 -197.565 190.465 -196.920 ;
        RECT 190.755 -197.045 190.925 -195.550 ;
        RECT 197.545 -196.670 197.715 -195.215 ;
        RECT 197.535 -197.225 197.720 -196.670 ;
        RECT 198.035 -196.755 198.205 -193.530 ;
        RECT 199.180 -193.880 199.370 -193.530 ;
        RECT 200.380 -193.720 200.550 -193.325 ;
        RECT 201.755 -193.370 202.445 -193.325 ;
        RECT 199.130 -194.570 199.400 -193.880 ;
        RECT 199.895 -193.890 200.550 -193.720 ;
        RECT 200.880 -193.805 201.570 -193.535 ;
        RECT 202.805 -193.880 203.075 -193.190 ;
        RECT 203.265 -193.195 203.435 -192.975 ;
        RECT 203.265 -193.465 204.095 -193.195 ;
        RECT 199.895 -196.755 200.065 -193.890 ;
        RECT 203.265 -194.040 203.435 -193.465 ;
        RECT 203.695 -194.040 203.965 -193.955 ;
        RECT 200.385 -194.235 201.180 -194.060 ;
        RECT 203.265 -194.065 203.965 -194.040 ;
        RECT 203.125 -194.210 203.965 -194.065 ;
        RECT 200.385 -196.755 200.555 -194.235 ;
        RECT 201.010 -196.755 201.180 -194.235 ;
        RECT 201.500 -196.670 201.670 -194.215 ;
        RECT 202.150 -196.665 202.320 -194.215 ;
        RECT 194.850 -197.245 197.905 -197.225 ;
        RECT 201.495 -197.245 201.680 -196.670 ;
        RECT 202.135 -197.245 202.320 -196.665 ;
        RECT 202.640 -196.755 202.810 -194.215 ;
        RECT 203.125 -194.235 203.435 -194.210 ;
        RECT 203.130 -196.755 203.300 -194.235 ;
        RECT 203.695 -194.250 203.965 -194.210 ;
        RECT 204.270 -194.800 204.460 -192.335 ;
        RECT 225.155 -193.305 225.325 -191.585 ;
        RECT 226.135 -193.305 226.305 -191.585 ;
        RECT 228.200 -192.120 228.370 -191.580 ;
        RECT 229.180 -192.120 229.350 -191.580 ;
        RECT 227.610 -192.355 227.975 -192.290 ;
        RECT 227.110 -192.495 227.975 -192.355 ;
        RECT 227.000 -192.560 227.975 -192.495 ;
        RECT 227.000 -193.305 227.305 -192.560 ;
        RECT 227.610 -192.590 227.975 -192.560 ;
        RECT 230.160 -192.440 230.330 -191.580 ;
        RECT 225.155 -193.455 227.305 -193.305 ;
        RECT 225.155 -193.495 227.250 -193.455 ;
        RECT 228.200 -193.515 228.370 -192.735 ;
        RECT 228.690 -193.275 228.860 -192.735 ;
        RECT 229.180 -193.515 229.350 -192.735 ;
        RECT 229.670 -193.275 229.840 -192.735 ;
        RECT 230.160 -192.790 231.550 -192.440 ;
        RECT 223.375 -193.860 224.510 -193.850 ;
        RECT 226.565 -193.860 226.935 -193.730 ;
        RECT 223.375 -194.050 226.935 -193.860 ;
        RECT 227.500 -193.945 230.575 -193.515 ;
        RECT 204.270 -194.990 205.730 -194.800 ;
        RECT 203.780 -196.660 203.950 -195.215 ;
        RECT 204.270 -195.240 204.460 -194.990 ;
        RECT 203.770 -197.245 203.955 -196.660 ;
        RECT 204.270 -196.755 204.440 -195.240 ;
        RECT 194.850 -197.565 204.520 -197.245 ;
        RECT 184.405 -197.790 204.520 -197.565 ;
        RECT 184.405 -198.130 195.415 -197.790 ;
        RECT 197.155 -198.050 204.520 -197.790 ;
        RECT 154.595 -201.490 154.785 -199.600 ;
        RECT 160.630 -201.095 163.955 -200.955 ;
        RECT 160.630 -201.385 165.805 -201.095 ;
        RECT 154.480 -201.760 154.845 -201.490 ;
        RECT 160.630 -201.790 161.060 -201.385 ;
        RECT 161.930 -201.570 162.105 -201.385 ;
        RECT 163.555 -201.400 165.805 -201.385 ;
        RECT 156.370 -202.220 161.060 -201.790 ;
        RECT 155.610 -203.340 156.260 -203.210 ;
        RECT 153.085 -203.670 156.260 -203.340 ;
        RECT 157.070 -203.500 157.240 -202.220 ;
        RECT 157.560 -203.500 157.730 -202.460 ;
        RECT 158.050 -203.500 158.220 -202.220 ;
        RECT 158.540 -203.330 158.710 -202.460 ;
        RECT 161.445 -203.110 161.615 -201.570 ;
        RECT 161.935 -203.110 162.105 -201.570 ;
        RECT 162.425 -203.110 162.595 -201.570 ;
        RECT 162.915 -203.110 163.085 -201.570 ;
        RECT 163.405 -203.110 163.575 -201.570 ;
        RECT 161.285 -203.325 161.640 -203.320 ;
        RECT 163.345 -203.325 163.715 -203.295 ;
        RECT 161.285 -203.330 163.715 -203.325 ;
        RECT 158.540 -203.500 163.715 -203.330 ;
        RECT 165.500 -203.435 165.805 -201.400 ;
        RECT 158.545 -203.520 163.715 -203.500 ;
        RECT 158.545 -203.530 161.290 -203.520 ;
        RECT 156.480 -203.670 156.845 -203.640 ;
        RECT 163.345 -203.650 163.715 -203.520 ;
        RECT 153.085 -203.720 156.845 -203.670 ;
        RECT 155.610 -203.875 156.845 -203.720 ;
        RECT 161.020 -203.810 161.695 -203.770 ;
        RECT 160.920 -203.820 161.695 -203.810 ;
        RECT 155.610 -203.960 156.260 -203.875 ;
        RECT 156.480 -203.940 156.845 -203.875 ;
        RECT 155.745 -204.210 156.125 -203.960 ;
        RECT 159.885 -204.000 161.695 -203.820 ;
        RECT 164.280 -203.865 168.205 -203.435 ;
        RECT 160.920 -204.010 161.695 -204.000 ;
        RECT 161.020 -204.040 161.695 -204.010 ;
        RECT 161.935 -203.925 164.030 -203.885 ;
        RECT 161.935 -204.075 164.085 -203.925 ;
        RECT 157.070 -205.150 157.240 -204.110 ;
        RECT 158.050 -205.150 158.220 -204.110 ;
        RECT 159.030 -205.150 159.200 -204.110 ;
        RECT 161.935 -205.795 162.105 -204.075 ;
        RECT 162.915 -205.795 163.085 -204.075 ;
        RECT 163.780 -204.820 164.085 -204.075 ;
        RECT 164.980 -204.645 165.150 -203.865 ;
        RECT 165.470 -204.645 165.640 -204.105 ;
        RECT 165.960 -204.645 166.130 -203.865 ;
        RECT 166.450 -204.645 166.620 -204.105 ;
        RECT 164.390 -204.820 164.755 -204.790 ;
        RECT 163.780 -204.885 164.755 -204.820 ;
        RECT 163.890 -205.025 164.755 -204.885 ;
        RECT 164.390 -205.090 164.755 -205.025 ;
        RECT 166.940 -204.940 168.800 -204.590 ;
        RECT 164.980 -205.800 165.150 -205.260 ;
        RECT 165.960 -205.800 166.130 -205.260 ;
        RECT 166.940 -205.800 167.110 -204.940 ;
        RECT 165.210 -208.140 166.410 -207.970 ;
        RECT 156.940 -210.475 157.110 -208.755 ;
        RECT 157.920 -210.475 158.090 -208.755 ;
        RECT 159.985 -209.290 160.155 -208.750 ;
        RECT 160.965 -209.290 161.135 -208.750 ;
        RECT 159.395 -209.525 159.760 -209.460 ;
        RECT 158.895 -209.665 159.760 -209.525 ;
        RECT 158.785 -209.730 159.760 -209.665 ;
        RECT 158.785 -210.475 159.090 -209.730 ;
        RECT 159.395 -209.760 159.760 -209.730 ;
        RECT 161.945 -209.610 162.115 -208.750 ;
        RECT 156.940 -210.625 159.090 -210.475 ;
        RECT 156.940 -210.665 159.035 -210.625 ;
        RECT 159.985 -210.685 160.155 -209.905 ;
        RECT 160.475 -210.445 160.645 -209.905 ;
        RECT 160.965 -210.685 161.135 -209.905 ;
        RECT 161.455 -210.445 161.625 -209.905 ;
        RECT 161.945 -209.960 163.335 -209.610 ;
        RECT 155.160 -211.030 156.295 -211.020 ;
        RECT 158.350 -211.030 158.720 -210.900 ;
        RECT 151.450 -211.315 152.875 -211.100 ;
        RECT 155.160 -211.220 158.720 -211.030 ;
        RECT 159.285 -211.115 162.360 -210.685 ;
        RECT 156.290 -211.225 158.720 -211.220 ;
        RECT 156.290 -211.230 156.645 -211.225 ;
        RECT 158.350 -211.255 158.720 -211.225 ;
        RECT 150.055 -211.830 150.580 -211.470 ;
        RECT 152.660 -212.345 152.875 -211.315 ;
        RECT 140.220 -213.085 142.470 -212.995 ;
        RECT 138.010 -213.300 142.470 -213.085 ;
        RECT 138.010 -213.390 140.255 -213.300 ;
        RECT 142.165 -214.775 142.470 -213.300 ;
        RECT 145.835 -214.185 146.005 -212.715 ;
        RECT 146.295 -212.795 146.520 -212.445 ;
        RECT 148.255 -212.545 152.875 -212.345 ;
        RECT 148.495 -212.560 152.875 -212.545 ;
        RECT 145.800 -214.775 146.035 -214.185 ;
        RECT 146.325 -214.255 146.495 -212.795 ;
        RECT 146.815 -214.180 146.985 -212.715 ;
        RECT 148.025 -214.130 148.195 -212.715 ;
        RECT 148.495 -212.760 148.715 -212.560 ;
        RECT 146.780 -214.775 147.015 -214.180 ;
        RECT 147.990 -214.775 148.225 -214.130 ;
        RECT 148.515 -214.255 148.685 -212.760 ;
        RECT 156.450 -212.980 156.620 -211.440 ;
        RECT 156.940 -212.980 157.110 -211.440 ;
        RECT 157.430 -212.980 157.600 -211.440 ;
        RECT 157.920 -212.980 158.090 -211.440 ;
        RECT 158.410 -212.980 158.580 -211.440 ;
        RECT 156.935 -213.240 157.110 -212.980 ;
        RECT 160.505 -213.150 160.810 -211.115 ;
        RECT 162.955 -211.935 163.305 -209.960 ;
        RECT 164.175 -211.230 164.345 -208.310 ;
        RECT 165.210 -208.350 165.420 -208.140 ;
        RECT 164.155 -211.525 164.365 -211.230 ;
        RECT 165.230 -211.260 165.400 -208.350 ;
        RECT 165.720 -211.250 165.890 -208.310 ;
        RECT 166.200 -208.360 166.410 -208.140 ;
        RECT 165.215 -211.525 165.425 -211.260 ;
        RECT 164.155 -211.705 165.425 -211.525 ;
        RECT 165.700 -211.520 165.910 -211.250 ;
        RECT 166.210 -211.350 166.380 -208.360 ;
        RECT 167.270 -211.280 167.440 -208.310 ;
        RECT 165.700 -211.715 166.405 -211.520 ;
        RECT 166.190 -211.775 166.405 -211.715 ;
        RECT 164.980 -211.935 165.755 -211.885 ;
        RECT 162.955 -212.115 165.755 -211.935 ;
        RECT 162.955 -212.125 163.305 -212.115 ;
        RECT 164.980 -212.160 165.755 -212.115 ;
        RECT 166.190 -212.050 167.095 -211.775 ;
        RECT 166.190 -212.400 166.405 -212.050 ;
        RECT 163.630 -212.470 164.405 -212.425 ;
        RECT 163.445 -212.640 164.405 -212.470 ;
        RECT 163.630 -212.700 164.405 -212.640 ;
        RECT 164.635 -212.600 166.405 -212.400 ;
        RECT 167.265 -212.500 167.480 -211.280 ;
        RECT 168.450 -211.625 168.800 -204.940 ;
        RECT 168.395 -211.985 168.920 -211.625 ;
        RECT 170.925 -212.500 172.040 -212.050 ;
        RECT 158.560 -213.240 160.810 -213.150 ;
        RECT 156.350 -213.455 160.810 -213.240 ;
        RECT 156.350 -213.545 158.595 -213.455 ;
        RECT 142.165 -215.340 149.550 -214.775 ;
        RECT 160.505 -214.930 160.810 -213.455 ;
        RECT 164.175 -214.340 164.345 -212.870 ;
        RECT 164.635 -212.950 164.860 -212.600 ;
        RECT 166.595 -212.700 172.605 -212.500 ;
        RECT 166.835 -212.715 172.605 -212.700 ;
        RECT 164.140 -214.930 164.375 -214.340 ;
        RECT 164.665 -214.410 164.835 -212.950 ;
        RECT 165.155 -214.335 165.325 -212.870 ;
        RECT 166.365 -214.285 166.535 -212.870 ;
        RECT 166.835 -212.915 167.055 -212.715 ;
        RECT 170.925 -212.900 172.040 -212.715 ;
        RECT 165.120 -214.930 165.355 -214.335 ;
        RECT 166.330 -214.930 166.565 -214.285 ;
        RECT 166.855 -214.410 167.025 -212.915 ;
        RECT 160.505 -215.495 167.890 -214.930 ;
        RECT 123.605 -218.650 133.665 -218.640 ;
        RECT 84.935 -218.865 85.105 -218.845 ;
        RECT 74.730 -219.130 77.870 -218.960 ;
        RECT 123.605 -219.490 133.760 -218.650 ;
        RECT 175.835 -218.750 176.565 -198.835 ;
        RECT 179.115 -199.495 179.495 -198.835 ;
        RECT 205.540 -199.465 205.730 -194.990 ;
        RECT 223.430 -198.740 223.810 -194.050 ;
        RECT 224.505 -194.055 226.935 -194.050 ;
        RECT 224.505 -194.060 224.860 -194.055 ;
        RECT 226.565 -194.085 226.935 -194.055 ;
        RECT 224.665 -195.810 224.835 -194.270 ;
        RECT 225.155 -195.810 225.325 -194.270 ;
        RECT 225.645 -195.810 225.815 -194.270 ;
        RECT 226.135 -195.810 226.305 -194.270 ;
        RECT 226.625 -195.810 226.795 -194.270 ;
        RECT 225.150 -196.070 225.325 -195.810 ;
        RECT 228.720 -195.980 229.025 -193.945 ;
        RECT 231.170 -194.765 231.520 -192.790 ;
        RECT 232.390 -194.060 232.560 -191.140 ;
        RECT 233.425 -191.180 233.635 -190.970 ;
        RECT 232.370 -194.355 232.580 -194.060 ;
        RECT 233.445 -194.090 233.615 -191.180 ;
        RECT 233.935 -194.080 234.105 -191.140 ;
        RECT 234.415 -191.190 234.625 -190.970 ;
        RECT 233.430 -194.355 233.640 -194.090 ;
        RECT 232.370 -194.535 233.640 -194.355 ;
        RECT 233.915 -194.350 234.125 -194.080 ;
        RECT 234.425 -194.180 234.595 -191.190 ;
        RECT 235.485 -194.110 235.655 -191.140 ;
        RECT 233.915 -194.545 234.620 -194.350 ;
        RECT 234.405 -194.605 234.620 -194.545 ;
        RECT 233.195 -194.765 233.970 -194.715 ;
        RECT 231.170 -194.945 233.970 -194.765 ;
        RECT 231.170 -194.955 231.520 -194.945 ;
        RECT 233.195 -194.990 233.970 -194.945 ;
        RECT 234.405 -194.880 235.310 -194.605 ;
        RECT 234.405 -195.230 234.620 -194.880 ;
        RECT 231.845 -195.300 232.620 -195.255 ;
        RECT 231.660 -195.470 232.620 -195.300 ;
        RECT 231.845 -195.530 232.620 -195.470 ;
        RECT 232.850 -195.430 234.620 -195.230 ;
        RECT 235.480 -195.330 235.695 -194.110 ;
        RECT 236.665 -194.455 237.015 -187.770 ;
        RECT 271.275 -187.810 271.445 -186.770 ;
        RECT 272.255 -187.810 272.425 -186.770 ;
        RECT 273.235 -187.810 273.405 -186.770 ;
        RECT 276.140 -188.455 276.310 -186.735 ;
        RECT 277.120 -188.455 277.290 -186.735 ;
        RECT 277.985 -187.480 278.290 -186.735 ;
        RECT 279.185 -187.305 279.355 -186.525 ;
        RECT 279.675 -187.305 279.845 -186.765 ;
        RECT 280.165 -187.305 280.335 -186.525 ;
        RECT 280.655 -187.305 280.825 -186.765 ;
        RECT 278.595 -187.480 278.960 -187.450 ;
        RECT 277.985 -187.545 278.960 -187.480 ;
        RECT 278.095 -187.685 278.960 -187.545 ;
        RECT 278.595 -187.750 278.960 -187.685 ;
        RECT 281.145 -187.600 283.005 -187.250 ;
        RECT 315.045 -187.480 315.215 -186.440 ;
        RECT 316.025 -187.480 316.195 -186.440 ;
        RECT 317.005 -187.480 317.175 -186.440 ;
        RECT 279.185 -188.460 279.355 -187.920 ;
        RECT 280.165 -188.460 280.335 -187.920 ;
        RECT 281.145 -188.460 281.315 -187.600 ;
        RECT 243.245 -190.250 244.850 -190.080 ;
        RECT 242.350 -192.930 242.520 -190.430 ;
        RECT 242.345 -193.160 242.520 -192.930 ;
        RECT 243.245 -193.160 243.445 -190.250 ;
        RECT 243.690 -190.450 243.865 -190.250 ;
        RECT 243.695 -192.970 243.865 -190.450 ;
        RECT 244.185 -192.935 244.355 -190.430 ;
        RECT 244.675 -190.445 244.850 -190.250 ;
        RECT 242.345 -193.360 243.445 -193.160 ;
        RECT 244.170 -193.535 244.360 -192.935 ;
        RECT 244.675 -192.970 244.845 -190.445 ;
        RECT 245.325 -193.350 245.495 -190.430 ;
        RECT 246.955 -193.000 247.125 -190.430 ;
        RECT 248.095 -191.880 248.265 -190.430 ;
        RECT 279.415 -190.800 280.615 -190.630 ;
        RECT 248.090 -192.345 248.275 -191.880 ;
        RECT 248.090 -192.530 248.775 -192.345 ;
        RECT 246.955 -193.170 247.750 -193.000 ;
        RECT 246.070 -193.350 246.760 -193.295 ;
        RECT 242.350 -193.725 244.360 -193.535 ;
        RECT 244.695 -193.520 246.760 -193.350 ;
        RECT 241.165 -193.780 241.855 -193.730 ;
        RECT 239.215 -193.950 241.855 -193.780 ;
        RECT 236.610 -194.815 237.135 -194.455 ;
        RECT 239.215 -195.330 239.430 -193.950 ;
        RECT 241.165 -194.000 241.855 -193.950 ;
        RECT 241.445 -194.455 242.135 -194.410 ;
        RECT 240.395 -194.625 242.135 -194.455 ;
        RECT 240.395 -195.260 240.755 -194.625 ;
        RECT 241.445 -194.680 242.135 -194.625 ;
        RECT 240.395 -195.305 240.815 -195.260 ;
        RECT 226.775 -196.070 229.025 -195.980 ;
        RECT 224.565 -196.285 229.025 -196.070 ;
        RECT 224.565 -196.375 226.810 -196.285 ;
        RECT 228.720 -197.760 229.025 -196.285 ;
        RECT 232.390 -197.170 232.560 -195.700 ;
        RECT 232.850 -195.780 233.075 -195.430 ;
        RECT 234.810 -195.530 239.430 -195.330 ;
        RECT 235.050 -195.545 239.430 -195.530 ;
        RECT 232.355 -197.760 232.590 -197.170 ;
        RECT 232.880 -197.240 233.050 -195.780 ;
        RECT 233.370 -197.165 233.540 -195.700 ;
        RECT 234.580 -197.115 234.750 -195.700 ;
        RECT 235.050 -195.745 235.270 -195.545 ;
        RECT 240.420 -195.655 240.815 -195.305 ;
        RECT 233.335 -197.760 233.570 -197.165 ;
        RECT 234.545 -197.760 234.780 -197.115 ;
        RECT 235.070 -197.240 235.240 -195.745 ;
        RECT 241.860 -196.865 242.030 -195.410 ;
        RECT 241.850 -197.420 242.035 -196.865 ;
        RECT 242.350 -196.950 242.520 -193.725 ;
        RECT 243.495 -194.075 243.685 -193.725 ;
        RECT 244.695 -193.915 244.865 -193.520 ;
        RECT 246.070 -193.565 246.760 -193.520 ;
        RECT 243.445 -194.765 243.715 -194.075 ;
        RECT 244.210 -194.085 244.865 -193.915 ;
        RECT 245.195 -194.000 245.885 -193.730 ;
        RECT 247.120 -194.075 247.390 -193.385 ;
        RECT 247.580 -193.390 247.750 -193.170 ;
        RECT 247.580 -193.660 248.410 -193.390 ;
        RECT 244.210 -196.950 244.380 -194.085 ;
        RECT 247.580 -194.235 247.750 -193.660 ;
        RECT 248.010 -194.235 248.280 -194.150 ;
        RECT 244.700 -194.430 245.495 -194.255 ;
        RECT 247.580 -194.260 248.280 -194.235 ;
        RECT 247.440 -194.405 248.280 -194.260 ;
        RECT 244.700 -196.950 244.870 -194.430 ;
        RECT 245.325 -196.950 245.495 -194.430 ;
        RECT 245.815 -196.865 245.985 -194.410 ;
        RECT 246.465 -196.860 246.635 -194.410 ;
        RECT 239.165 -197.440 242.220 -197.420 ;
        RECT 245.810 -197.440 245.995 -196.865 ;
        RECT 246.450 -197.440 246.635 -196.860 ;
        RECT 246.955 -196.950 247.125 -194.410 ;
        RECT 247.440 -194.430 247.750 -194.405 ;
        RECT 247.445 -196.950 247.615 -194.430 ;
        RECT 248.010 -194.445 248.280 -194.405 ;
        RECT 248.585 -194.995 248.775 -192.530 ;
        RECT 271.145 -193.135 271.315 -191.415 ;
        RECT 272.125 -193.135 272.295 -191.415 ;
        RECT 274.190 -191.950 274.360 -191.410 ;
        RECT 275.170 -191.950 275.340 -191.410 ;
        RECT 273.600 -192.185 273.965 -192.120 ;
        RECT 273.100 -192.325 273.965 -192.185 ;
        RECT 272.990 -192.390 273.965 -192.325 ;
        RECT 272.990 -193.135 273.295 -192.390 ;
        RECT 273.600 -192.420 273.965 -192.390 ;
        RECT 276.150 -192.270 276.320 -191.410 ;
        RECT 271.145 -193.285 273.295 -193.135 ;
        RECT 271.145 -193.325 273.240 -193.285 ;
        RECT 274.190 -193.345 274.360 -192.565 ;
        RECT 274.680 -193.105 274.850 -192.565 ;
        RECT 275.170 -193.345 275.340 -192.565 ;
        RECT 275.660 -193.105 275.830 -192.565 ;
        RECT 276.150 -192.620 277.540 -192.270 ;
        RECT 269.365 -193.690 270.500 -193.680 ;
        RECT 272.555 -193.690 272.925 -193.560 ;
        RECT 269.365 -193.880 272.925 -193.690 ;
        RECT 273.490 -193.775 276.565 -193.345 ;
        RECT 248.585 -195.185 250.045 -194.995 ;
        RECT 248.095 -196.855 248.265 -195.410 ;
        RECT 248.585 -195.435 248.775 -195.185 ;
        RECT 248.085 -197.440 248.270 -196.855 ;
        RECT 248.585 -196.950 248.755 -195.435 ;
        RECT 239.165 -197.760 248.835 -197.440 ;
        RECT 228.720 -197.985 248.835 -197.760 ;
        RECT 228.720 -198.325 239.730 -197.985 ;
        RECT 241.470 -198.245 248.835 -197.985 ;
        RECT 179.115 -199.875 195.665 -199.495 ;
        RECT 179.115 -200.785 179.495 -199.875 ;
        RECT 179.115 -201.165 179.825 -200.785 ;
        RECT 179.445 -203.110 179.825 -201.165 ;
        RECT 184.490 -200.995 187.815 -200.855 ;
        RECT 184.490 -201.285 189.665 -200.995 ;
        RECT 193.535 -201.280 193.995 -200.855 ;
        RECT 184.490 -201.690 184.920 -201.285 ;
        RECT 185.790 -201.470 185.965 -201.285 ;
        RECT 187.415 -201.300 189.665 -201.285 ;
        RECT 180.230 -202.120 184.920 -201.690 ;
        RECT 179.445 -203.570 180.120 -203.110 ;
        RECT 180.930 -203.400 181.100 -202.120 ;
        RECT 181.420 -203.400 181.590 -202.360 ;
        RECT 181.910 -203.400 182.080 -202.120 ;
        RECT 182.400 -203.230 182.570 -202.360 ;
        RECT 185.305 -203.010 185.475 -201.470 ;
        RECT 185.795 -203.010 185.965 -201.470 ;
        RECT 186.285 -203.010 186.455 -201.470 ;
        RECT 186.775 -203.010 186.945 -201.470 ;
        RECT 187.265 -203.010 187.435 -201.470 ;
        RECT 185.145 -203.225 185.500 -203.220 ;
        RECT 187.205 -203.225 187.575 -203.195 ;
        RECT 185.145 -203.230 187.575 -203.225 ;
        RECT 182.400 -203.400 187.575 -203.230 ;
        RECT 189.360 -203.335 189.665 -201.300 ;
        RECT 182.405 -203.420 187.575 -203.400 ;
        RECT 182.405 -203.430 185.150 -203.420 ;
        RECT 180.340 -203.570 180.705 -203.540 ;
        RECT 187.205 -203.550 187.575 -203.420 ;
        RECT 179.445 -203.655 180.705 -203.570 ;
        RECT 179.470 -203.775 180.705 -203.655 ;
        RECT 184.880 -203.710 185.555 -203.670 ;
        RECT 184.780 -203.720 185.555 -203.710 ;
        RECT 179.470 -203.860 180.120 -203.775 ;
        RECT 180.340 -203.840 180.705 -203.775 ;
        RECT 183.745 -203.900 185.555 -203.720 ;
        RECT 188.140 -203.765 192.065 -203.335 ;
        RECT 184.780 -203.910 185.555 -203.900 ;
        RECT 184.880 -203.940 185.555 -203.910 ;
        RECT 185.795 -203.825 187.890 -203.785 ;
        RECT 185.795 -203.975 187.945 -203.825 ;
        RECT 180.930 -205.050 181.100 -204.010 ;
        RECT 181.910 -205.050 182.080 -204.010 ;
        RECT 182.890 -205.050 183.060 -204.010 ;
        RECT 185.795 -205.695 185.965 -203.975 ;
        RECT 186.775 -205.695 186.945 -203.975 ;
        RECT 187.640 -204.720 187.945 -203.975 ;
        RECT 188.840 -204.545 189.010 -203.765 ;
        RECT 189.330 -204.545 189.500 -204.005 ;
        RECT 189.820 -204.545 189.990 -203.765 ;
        RECT 190.310 -204.545 190.480 -204.005 ;
        RECT 188.250 -204.720 188.615 -204.690 ;
        RECT 187.640 -204.785 188.615 -204.720 ;
        RECT 187.750 -204.925 188.615 -204.785 ;
        RECT 188.250 -204.990 188.615 -204.925 ;
        RECT 190.800 -204.840 192.660 -204.490 ;
        RECT 188.840 -205.700 189.010 -205.160 ;
        RECT 189.820 -205.700 189.990 -205.160 ;
        RECT 190.800 -205.700 190.970 -204.840 ;
        RECT 189.070 -208.040 190.270 -207.870 ;
        RECT 180.800 -210.375 180.970 -208.655 ;
        RECT 181.780 -210.375 181.950 -208.655 ;
        RECT 183.845 -209.190 184.015 -208.650 ;
        RECT 184.825 -209.190 184.995 -208.650 ;
        RECT 183.255 -209.425 183.620 -209.360 ;
        RECT 182.755 -209.565 183.620 -209.425 ;
        RECT 182.645 -209.630 183.620 -209.565 ;
        RECT 182.645 -210.375 182.950 -209.630 ;
        RECT 183.255 -209.660 183.620 -209.630 ;
        RECT 185.805 -209.510 185.975 -208.650 ;
        RECT 180.800 -210.525 182.950 -210.375 ;
        RECT 180.800 -210.565 182.895 -210.525 ;
        RECT 183.845 -210.585 184.015 -209.805 ;
        RECT 184.335 -210.345 184.505 -209.805 ;
        RECT 184.825 -210.585 184.995 -209.805 ;
        RECT 185.315 -210.345 185.485 -209.805 ;
        RECT 185.805 -209.860 187.195 -209.510 ;
        RECT 179.020 -210.930 180.155 -210.920 ;
        RECT 182.210 -210.930 182.580 -210.800 ;
        RECT 179.020 -211.120 182.580 -210.930 ;
        RECT 183.145 -211.015 186.220 -210.585 ;
        RECT 180.150 -211.125 182.580 -211.120 ;
        RECT 180.150 -211.130 180.505 -211.125 ;
        RECT 182.210 -211.155 182.580 -211.125 ;
        RECT 180.310 -212.880 180.480 -211.340 ;
        RECT 180.800 -212.880 180.970 -211.340 ;
        RECT 181.290 -212.880 181.460 -211.340 ;
        RECT 181.780 -212.880 181.950 -211.340 ;
        RECT 182.270 -212.880 182.440 -211.340 ;
        RECT 180.795 -213.140 180.970 -212.880 ;
        RECT 184.365 -213.050 184.670 -211.015 ;
        RECT 186.815 -211.835 187.165 -209.860 ;
        RECT 188.035 -211.130 188.205 -208.210 ;
        RECT 189.070 -208.250 189.280 -208.040 ;
        RECT 188.015 -211.425 188.225 -211.130 ;
        RECT 189.090 -211.160 189.260 -208.250 ;
        RECT 189.580 -211.150 189.750 -208.210 ;
        RECT 190.060 -208.260 190.270 -208.040 ;
        RECT 189.075 -211.425 189.285 -211.160 ;
        RECT 188.015 -211.605 189.285 -211.425 ;
        RECT 189.560 -211.420 189.770 -211.150 ;
        RECT 190.070 -211.250 190.240 -208.260 ;
        RECT 191.130 -211.180 191.300 -208.210 ;
        RECT 189.560 -211.615 190.265 -211.420 ;
        RECT 190.050 -211.675 190.265 -211.615 ;
        RECT 188.840 -211.835 189.615 -211.785 ;
        RECT 186.815 -212.015 189.615 -211.835 ;
        RECT 186.815 -212.025 187.165 -212.015 ;
        RECT 188.840 -212.060 189.615 -212.015 ;
        RECT 190.050 -211.950 190.955 -211.675 ;
        RECT 190.050 -212.300 190.265 -211.950 ;
        RECT 187.490 -212.370 188.265 -212.325 ;
        RECT 187.305 -212.540 188.265 -212.370 ;
        RECT 187.490 -212.600 188.265 -212.540 ;
        RECT 188.495 -212.500 190.265 -212.300 ;
        RECT 191.125 -212.400 191.340 -211.180 ;
        RECT 192.310 -211.525 192.660 -204.840 ;
        RECT 193.650 -211.155 193.865 -201.280 ;
        RECT 195.285 -203.395 195.665 -199.875 ;
        RECT 196.795 -199.655 205.730 -199.465 ;
        RECT 220.180 -199.470 223.810 -198.740 ;
        RECT 196.795 -201.545 196.985 -199.655 ;
        RECT 202.830 -201.150 206.155 -201.010 ;
        RECT 202.830 -201.440 208.005 -201.150 ;
        RECT 196.680 -201.815 197.045 -201.545 ;
        RECT 202.830 -201.845 203.260 -201.440 ;
        RECT 204.130 -201.625 204.305 -201.440 ;
        RECT 205.755 -201.455 208.005 -201.440 ;
        RECT 198.570 -202.275 203.260 -201.845 ;
        RECT 197.810 -203.395 198.460 -203.265 ;
        RECT 195.285 -203.725 198.460 -203.395 ;
        RECT 199.270 -203.555 199.440 -202.275 ;
        RECT 199.760 -203.555 199.930 -202.515 ;
        RECT 200.250 -203.555 200.420 -202.275 ;
        RECT 200.740 -203.385 200.910 -202.515 ;
        RECT 203.645 -203.165 203.815 -201.625 ;
        RECT 204.135 -203.165 204.305 -201.625 ;
        RECT 204.625 -203.165 204.795 -201.625 ;
        RECT 205.115 -203.165 205.285 -201.625 ;
        RECT 205.605 -203.165 205.775 -201.625 ;
        RECT 203.485 -203.380 203.840 -203.375 ;
        RECT 205.545 -203.380 205.915 -203.350 ;
        RECT 203.485 -203.385 205.915 -203.380 ;
        RECT 200.740 -203.555 205.915 -203.385 ;
        RECT 207.700 -203.490 208.005 -201.455 ;
        RECT 200.745 -203.575 205.915 -203.555 ;
        RECT 200.745 -203.585 203.490 -203.575 ;
        RECT 198.680 -203.725 199.045 -203.695 ;
        RECT 205.545 -203.705 205.915 -203.575 ;
        RECT 195.285 -203.775 199.045 -203.725 ;
        RECT 197.810 -203.930 199.045 -203.775 ;
        RECT 203.220 -203.865 203.895 -203.825 ;
        RECT 203.120 -203.875 203.895 -203.865 ;
        RECT 197.810 -204.015 198.460 -203.930 ;
        RECT 198.680 -203.995 199.045 -203.930 ;
        RECT 197.945 -204.265 198.325 -204.015 ;
        RECT 202.085 -204.055 203.895 -203.875 ;
        RECT 206.480 -203.920 210.405 -203.490 ;
        RECT 203.120 -204.065 203.895 -204.055 ;
        RECT 203.220 -204.095 203.895 -204.065 ;
        RECT 204.135 -203.980 206.230 -203.940 ;
        RECT 204.135 -204.130 206.285 -203.980 ;
        RECT 199.270 -205.205 199.440 -204.165 ;
        RECT 200.250 -205.205 200.420 -204.165 ;
        RECT 201.230 -205.205 201.400 -204.165 ;
        RECT 204.135 -205.850 204.305 -204.130 ;
        RECT 205.115 -205.850 205.285 -204.130 ;
        RECT 205.980 -204.875 206.285 -204.130 ;
        RECT 207.180 -204.700 207.350 -203.920 ;
        RECT 207.670 -204.700 207.840 -204.160 ;
        RECT 208.160 -204.700 208.330 -203.920 ;
        RECT 208.650 -204.700 208.820 -204.160 ;
        RECT 206.590 -204.875 206.955 -204.845 ;
        RECT 205.980 -204.940 206.955 -204.875 ;
        RECT 206.090 -205.080 206.955 -204.940 ;
        RECT 206.590 -205.145 206.955 -205.080 ;
        RECT 209.140 -204.995 211.000 -204.645 ;
        RECT 207.180 -205.855 207.350 -205.315 ;
        RECT 208.160 -205.855 208.330 -205.315 ;
        RECT 209.140 -205.855 209.310 -204.995 ;
        RECT 207.410 -208.195 208.610 -208.025 ;
        RECT 199.140 -210.530 199.310 -208.810 ;
        RECT 200.120 -210.530 200.290 -208.810 ;
        RECT 202.185 -209.345 202.355 -208.805 ;
        RECT 203.165 -209.345 203.335 -208.805 ;
        RECT 201.595 -209.580 201.960 -209.515 ;
        RECT 201.095 -209.720 201.960 -209.580 ;
        RECT 200.985 -209.785 201.960 -209.720 ;
        RECT 200.985 -210.530 201.290 -209.785 ;
        RECT 201.595 -209.815 201.960 -209.785 ;
        RECT 204.145 -209.665 204.315 -208.805 ;
        RECT 199.140 -210.680 201.290 -210.530 ;
        RECT 199.140 -210.720 201.235 -210.680 ;
        RECT 202.185 -210.740 202.355 -209.960 ;
        RECT 202.675 -210.500 202.845 -209.960 ;
        RECT 203.165 -210.740 203.335 -209.960 ;
        RECT 203.655 -210.500 203.825 -209.960 ;
        RECT 204.145 -210.015 205.535 -209.665 ;
        RECT 197.360 -211.085 198.495 -211.075 ;
        RECT 200.550 -211.085 200.920 -210.955 ;
        RECT 193.650 -211.370 195.075 -211.155 ;
        RECT 197.360 -211.275 200.920 -211.085 ;
        RECT 201.485 -211.170 204.560 -210.740 ;
        RECT 198.490 -211.280 200.920 -211.275 ;
        RECT 198.490 -211.285 198.845 -211.280 ;
        RECT 200.550 -211.310 200.920 -211.280 ;
        RECT 192.255 -211.885 192.780 -211.525 ;
        RECT 194.860 -212.400 195.075 -211.370 ;
        RECT 182.420 -213.140 184.670 -213.050 ;
        RECT 180.210 -213.355 184.670 -213.140 ;
        RECT 180.210 -213.445 182.455 -213.355 ;
        RECT 184.365 -214.830 184.670 -213.355 ;
        RECT 188.035 -214.240 188.205 -212.770 ;
        RECT 188.495 -212.850 188.720 -212.500 ;
        RECT 190.455 -212.600 195.075 -212.400 ;
        RECT 190.695 -212.615 195.075 -212.600 ;
        RECT 188.000 -214.830 188.235 -214.240 ;
        RECT 188.525 -214.310 188.695 -212.850 ;
        RECT 189.015 -214.235 189.185 -212.770 ;
        RECT 190.225 -214.185 190.395 -212.770 ;
        RECT 190.695 -212.815 190.915 -212.615 ;
        RECT 188.980 -214.830 189.215 -214.235 ;
        RECT 190.190 -214.830 190.425 -214.185 ;
        RECT 190.715 -214.310 190.885 -212.815 ;
        RECT 198.650 -213.035 198.820 -211.495 ;
        RECT 199.140 -213.035 199.310 -211.495 ;
        RECT 199.630 -213.035 199.800 -211.495 ;
        RECT 200.120 -213.035 200.290 -211.495 ;
        RECT 200.610 -213.035 200.780 -211.495 ;
        RECT 199.135 -213.295 199.310 -213.035 ;
        RECT 202.705 -213.205 203.010 -211.170 ;
        RECT 205.155 -211.990 205.505 -210.015 ;
        RECT 206.375 -211.285 206.545 -208.365 ;
        RECT 207.410 -208.405 207.620 -208.195 ;
        RECT 206.355 -211.580 206.565 -211.285 ;
        RECT 207.430 -211.315 207.600 -208.405 ;
        RECT 207.920 -211.305 208.090 -208.365 ;
        RECT 208.400 -208.415 208.610 -208.195 ;
        RECT 207.415 -211.580 207.625 -211.315 ;
        RECT 206.355 -211.760 207.625 -211.580 ;
        RECT 207.900 -211.575 208.110 -211.305 ;
        RECT 208.410 -211.405 208.580 -208.415 ;
        RECT 209.470 -211.335 209.640 -208.365 ;
        RECT 207.900 -211.770 208.605 -211.575 ;
        RECT 208.390 -211.830 208.605 -211.770 ;
        RECT 207.180 -211.990 207.955 -211.940 ;
        RECT 205.155 -212.170 207.955 -211.990 ;
        RECT 205.155 -212.180 205.505 -212.170 ;
        RECT 207.180 -212.215 207.955 -212.170 ;
        RECT 208.390 -212.105 209.295 -211.830 ;
        RECT 208.390 -212.455 208.605 -212.105 ;
        RECT 205.830 -212.525 206.605 -212.480 ;
        RECT 205.645 -212.695 206.605 -212.525 ;
        RECT 205.830 -212.755 206.605 -212.695 ;
        RECT 206.835 -212.655 208.605 -212.455 ;
        RECT 209.465 -212.555 209.680 -211.335 ;
        RECT 210.650 -211.680 211.000 -204.995 ;
        RECT 210.595 -212.040 211.120 -211.680 ;
        RECT 213.170 -212.555 214.855 -211.740 ;
        RECT 200.760 -213.295 203.010 -213.205 ;
        RECT 198.550 -213.510 203.010 -213.295 ;
        RECT 198.550 -213.600 200.795 -213.510 ;
        RECT 184.365 -215.395 191.750 -214.830 ;
        RECT 202.705 -214.985 203.010 -213.510 ;
        RECT 206.375 -214.395 206.545 -212.925 ;
        RECT 206.835 -213.005 207.060 -212.655 ;
        RECT 208.795 -212.755 214.855 -212.555 ;
        RECT 209.035 -212.770 214.855 -212.755 ;
        RECT 206.340 -214.985 206.575 -214.395 ;
        RECT 206.865 -214.465 207.035 -213.005 ;
        RECT 207.355 -214.390 207.525 -212.925 ;
        RECT 208.565 -214.340 208.735 -212.925 ;
        RECT 209.035 -212.970 209.255 -212.770 ;
        RECT 207.320 -214.985 207.555 -214.390 ;
        RECT 208.530 -214.985 208.765 -214.340 ;
        RECT 209.055 -214.465 209.225 -212.970 ;
        RECT 213.170 -213.395 214.855 -212.770 ;
        RECT 202.705 -215.550 210.090 -214.985 ;
        RECT 175.720 -219.485 176.735 -218.750 ;
        RECT 123.605 -219.495 133.380 -219.490 ;
        RECT 211.375 -219.655 212.960 -218.200 ;
        RECT 220.180 -219.475 220.910 -199.470 ;
        RECT 223.430 -199.690 223.810 -199.470 ;
        RECT 249.855 -199.660 250.045 -195.185 ;
        RECT 269.420 -198.235 269.800 -193.880 ;
        RECT 270.495 -193.885 272.925 -193.880 ;
        RECT 270.495 -193.890 270.850 -193.885 ;
        RECT 272.555 -193.915 272.925 -193.885 ;
        RECT 270.655 -195.640 270.825 -194.100 ;
        RECT 271.145 -195.640 271.315 -194.100 ;
        RECT 271.635 -195.640 271.805 -194.100 ;
        RECT 272.125 -195.640 272.295 -194.100 ;
        RECT 272.615 -195.640 272.785 -194.100 ;
        RECT 271.140 -195.900 271.315 -195.640 ;
        RECT 274.710 -195.810 275.015 -193.775 ;
        RECT 277.160 -194.595 277.510 -192.620 ;
        RECT 278.380 -193.890 278.550 -190.970 ;
        RECT 279.415 -191.010 279.625 -190.800 ;
        RECT 278.360 -194.185 278.570 -193.890 ;
        RECT 279.435 -193.920 279.605 -191.010 ;
        RECT 279.925 -193.910 280.095 -190.970 ;
        RECT 280.405 -191.020 280.615 -190.800 ;
        RECT 279.420 -194.185 279.630 -193.920 ;
        RECT 278.360 -194.365 279.630 -194.185 ;
        RECT 279.905 -194.180 280.115 -193.910 ;
        RECT 280.415 -194.010 280.585 -191.020 ;
        RECT 281.475 -193.940 281.645 -190.970 ;
        RECT 279.905 -194.375 280.610 -194.180 ;
        RECT 280.395 -194.435 280.610 -194.375 ;
        RECT 279.185 -194.595 279.960 -194.545 ;
        RECT 277.160 -194.775 279.960 -194.595 ;
        RECT 277.160 -194.785 277.510 -194.775 ;
        RECT 279.185 -194.820 279.960 -194.775 ;
        RECT 280.395 -194.710 281.300 -194.435 ;
        RECT 280.395 -195.060 280.610 -194.710 ;
        RECT 277.835 -195.130 278.610 -195.085 ;
        RECT 277.650 -195.300 278.610 -195.130 ;
        RECT 277.835 -195.360 278.610 -195.300 ;
        RECT 278.840 -195.260 280.610 -195.060 ;
        RECT 281.470 -195.160 281.685 -193.940 ;
        RECT 282.655 -194.285 283.005 -187.600 ;
        RECT 319.910 -188.125 320.080 -186.405 ;
        RECT 320.890 -188.125 321.060 -186.405 ;
        RECT 321.755 -187.150 322.060 -186.405 ;
        RECT 322.955 -186.975 323.125 -186.195 ;
        RECT 323.445 -186.975 323.615 -186.435 ;
        RECT 323.935 -186.975 324.105 -186.195 ;
        RECT 359.350 -186.205 360.000 -186.120 ;
        RECT 360.220 -186.185 360.585 -186.120 ;
        RECT 363.625 -186.245 365.435 -186.065 ;
        RECT 368.020 -186.110 371.945 -185.680 ;
        RECT 406.170 -185.725 406.820 -185.265 ;
        RECT 407.630 -185.555 407.800 -184.275 ;
        RECT 408.120 -185.555 408.290 -184.515 ;
        RECT 408.610 -185.555 408.780 -184.275 ;
        RECT 409.100 -185.385 409.270 -184.515 ;
        RECT 412.005 -185.165 412.175 -183.625 ;
        RECT 412.495 -185.165 412.665 -183.625 ;
        RECT 412.985 -185.165 413.155 -183.625 ;
        RECT 413.475 -185.165 413.645 -183.625 ;
        RECT 413.965 -185.165 414.135 -183.625 ;
        RECT 411.845 -185.380 412.200 -185.375 ;
        RECT 413.905 -185.380 414.275 -185.350 ;
        RECT 411.845 -185.385 414.275 -185.380 ;
        RECT 409.100 -185.555 414.275 -185.385 ;
        RECT 416.060 -185.490 416.365 -183.455 ;
        RECT 409.105 -185.575 414.275 -185.555 ;
        RECT 409.105 -185.585 411.850 -185.575 ;
        RECT 407.040 -185.725 407.405 -185.695 ;
        RECT 413.905 -185.705 414.275 -185.575 ;
        RECT 406.170 -185.930 407.405 -185.725 ;
        RECT 411.580 -185.865 412.255 -185.825 ;
        RECT 411.480 -185.875 412.255 -185.865 ;
        RECT 406.170 -186.015 406.820 -185.930 ;
        RECT 407.040 -185.995 407.405 -185.930 ;
        RECT 410.445 -186.055 412.255 -185.875 ;
        RECT 414.840 -185.920 418.765 -185.490 ;
        RECT 411.480 -186.065 412.255 -186.055 ;
        RECT 411.580 -186.095 412.255 -186.065 ;
        RECT 412.495 -185.980 414.590 -185.940 ;
        RECT 364.660 -186.255 365.435 -186.245 ;
        RECT 364.760 -186.285 365.435 -186.255 ;
        RECT 365.675 -186.170 367.770 -186.130 ;
        RECT 365.675 -186.320 367.825 -186.170 ;
        RECT 324.425 -186.975 324.595 -186.435 ;
        RECT 322.365 -187.150 322.730 -187.120 ;
        RECT 321.755 -187.215 322.730 -187.150 ;
        RECT 321.865 -187.355 322.730 -187.215 ;
        RECT 322.365 -187.420 322.730 -187.355 ;
        RECT 324.915 -187.270 326.775 -186.920 ;
        RECT 322.955 -188.130 323.125 -187.590 ;
        RECT 323.935 -188.130 324.105 -187.590 ;
        RECT 324.915 -188.130 325.085 -187.270 ;
        RECT 289.235 -190.080 290.840 -189.910 ;
        RECT 288.340 -192.760 288.510 -190.260 ;
        RECT 288.335 -192.990 288.510 -192.760 ;
        RECT 289.235 -192.990 289.435 -190.080 ;
        RECT 289.680 -190.280 289.855 -190.080 ;
        RECT 289.685 -192.800 289.855 -190.280 ;
        RECT 290.175 -192.765 290.345 -190.260 ;
        RECT 290.665 -190.275 290.840 -190.080 ;
        RECT 288.335 -193.190 289.435 -192.990 ;
        RECT 290.160 -193.365 290.350 -192.765 ;
        RECT 290.665 -192.800 290.835 -190.275 ;
        RECT 291.315 -193.180 291.485 -190.260 ;
        RECT 292.945 -192.830 293.115 -190.260 ;
        RECT 294.085 -191.710 294.255 -190.260 ;
        RECT 323.185 -190.470 324.385 -190.300 ;
        RECT 294.080 -192.175 294.265 -191.710 ;
        RECT 294.080 -192.360 294.765 -192.175 ;
        RECT 292.945 -193.000 293.740 -192.830 ;
        RECT 292.060 -193.180 292.750 -193.125 ;
        RECT 288.340 -193.555 290.350 -193.365 ;
        RECT 290.685 -193.350 292.750 -193.180 ;
        RECT 287.155 -193.610 287.845 -193.560 ;
        RECT 285.205 -193.780 287.845 -193.610 ;
        RECT 282.600 -194.645 283.125 -194.285 ;
        RECT 285.205 -195.160 285.420 -193.780 ;
        RECT 287.155 -193.830 287.845 -193.780 ;
        RECT 287.435 -194.285 288.125 -194.240 ;
        RECT 286.385 -194.455 288.125 -194.285 ;
        RECT 286.385 -195.090 286.745 -194.455 ;
        RECT 287.435 -194.510 288.125 -194.455 ;
        RECT 286.385 -195.135 286.805 -195.090 ;
        RECT 272.765 -195.900 275.015 -195.810 ;
        RECT 270.555 -196.115 275.015 -195.900 ;
        RECT 270.555 -196.205 272.800 -196.115 ;
        RECT 274.710 -197.590 275.015 -196.115 ;
        RECT 278.380 -197.000 278.550 -195.530 ;
        RECT 278.840 -195.610 279.065 -195.260 ;
        RECT 280.800 -195.360 285.420 -195.160 ;
        RECT 281.040 -195.375 285.420 -195.360 ;
        RECT 278.345 -197.590 278.580 -197.000 ;
        RECT 278.870 -197.070 279.040 -195.610 ;
        RECT 279.360 -196.995 279.530 -195.530 ;
        RECT 280.570 -196.945 280.740 -195.530 ;
        RECT 281.040 -195.575 281.260 -195.375 ;
        RECT 286.410 -195.485 286.805 -195.135 ;
        RECT 279.325 -197.590 279.560 -196.995 ;
        RECT 280.535 -197.590 280.770 -196.945 ;
        RECT 281.060 -197.070 281.230 -195.575 ;
        RECT 287.850 -196.695 288.020 -195.240 ;
        RECT 287.840 -197.250 288.025 -196.695 ;
        RECT 288.340 -196.780 288.510 -193.555 ;
        RECT 289.485 -193.905 289.675 -193.555 ;
        RECT 290.685 -193.745 290.855 -193.350 ;
        RECT 292.060 -193.395 292.750 -193.350 ;
        RECT 289.435 -194.595 289.705 -193.905 ;
        RECT 290.200 -193.915 290.855 -193.745 ;
        RECT 291.185 -193.830 291.875 -193.560 ;
        RECT 293.110 -193.905 293.380 -193.215 ;
        RECT 293.570 -193.220 293.740 -193.000 ;
        RECT 293.570 -193.490 294.400 -193.220 ;
        RECT 290.200 -196.780 290.370 -193.915 ;
        RECT 293.570 -194.065 293.740 -193.490 ;
        RECT 294.000 -194.065 294.270 -193.980 ;
        RECT 290.690 -194.260 291.485 -194.085 ;
        RECT 293.570 -194.090 294.270 -194.065 ;
        RECT 293.430 -194.235 294.270 -194.090 ;
        RECT 290.690 -196.780 290.860 -194.260 ;
        RECT 291.315 -196.780 291.485 -194.260 ;
        RECT 291.805 -196.695 291.975 -194.240 ;
        RECT 292.455 -196.690 292.625 -194.240 ;
        RECT 285.155 -197.270 288.210 -197.250 ;
        RECT 291.800 -197.270 291.985 -196.695 ;
        RECT 292.440 -197.270 292.625 -196.690 ;
        RECT 292.945 -196.780 293.115 -194.240 ;
        RECT 293.430 -194.260 293.740 -194.235 ;
        RECT 293.435 -196.780 293.605 -194.260 ;
        RECT 294.000 -194.275 294.270 -194.235 ;
        RECT 294.575 -194.825 294.765 -192.360 ;
        RECT 314.915 -192.805 315.085 -191.085 ;
        RECT 315.895 -192.805 316.065 -191.085 ;
        RECT 317.960 -191.620 318.130 -191.080 ;
        RECT 318.940 -191.620 319.110 -191.080 ;
        RECT 317.370 -191.855 317.735 -191.790 ;
        RECT 316.870 -191.995 317.735 -191.855 ;
        RECT 316.760 -192.060 317.735 -191.995 ;
        RECT 316.760 -192.805 317.065 -192.060 ;
        RECT 317.370 -192.090 317.735 -192.060 ;
        RECT 319.920 -191.940 320.090 -191.080 ;
        RECT 314.915 -192.955 317.065 -192.805 ;
        RECT 314.915 -192.995 317.010 -192.955 ;
        RECT 317.960 -193.015 318.130 -192.235 ;
        RECT 318.450 -192.775 318.620 -192.235 ;
        RECT 318.940 -193.015 319.110 -192.235 ;
        RECT 319.430 -192.775 319.600 -192.235 ;
        RECT 319.920 -192.290 321.310 -191.940 ;
        RECT 313.135 -193.360 314.270 -193.350 ;
        RECT 316.325 -193.360 316.695 -193.230 ;
        RECT 313.135 -193.550 316.695 -193.360 ;
        RECT 317.260 -193.445 320.335 -193.015 ;
        RECT 294.575 -195.015 296.035 -194.825 ;
        RECT 294.085 -196.685 294.255 -195.240 ;
        RECT 294.575 -195.265 294.765 -195.015 ;
        RECT 294.075 -197.270 294.260 -196.685 ;
        RECT 294.575 -196.780 294.745 -195.265 ;
        RECT 285.155 -197.590 294.825 -197.270 ;
        RECT 274.710 -197.815 294.825 -197.590 ;
        RECT 274.710 -198.155 285.720 -197.815 ;
        RECT 287.460 -198.075 294.825 -197.815 ;
        RECT 223.430 -200.070 239.980 -199.690 ;
        RECT 223.430 -200.980 223.810 -200.070 ;
        RECT 223.430 -201.360 224.140 -200.980 ;
        RECT 223.760 -203.305 224.140 -201.360 ;
        RECT 228.805 -201.190 232.130 -201.050 ;
        RECT 228.805 -201.480 233.980 -201.190 ;
        RECT 237.850 -201.475 238.310 -201.050 ;
        RECT 228.805 -201.885 229.235 -201.480 ;
        RECT 230.105 -201.665 230.280 -201.480 ;
        RECT 231.730 -201.495 233.980 -201.480 ;
        RECT 224.545 -202.315 229.235 -201.885 ;
        RECT 223.760 -203.765 224.435 -203.305 ;
        RECT 225.245 -203.595 225.415 -202.315 ;
        RECT 225.735 -203.595 225.905 -202.555 ;
        RECT 226.225 -203.595 226.395 -202.315 ;
        RECT 226.715 -203.425 226.885 -202.555 ;
        RECT 229.620 -203.205 229.790 -201.665 ;
        RECT 230.110 -203.205 230.280 -201.665 ;
        RECT 230.600 -203.205 230.770 -201.665 ;
        RECT 231.090 -203.205 231.260 -201.665 ;
        RECT 231.580 -203.205 231.750 -201.665 ;
        RECT 229.460 -203.420 229.815 -203.415 ;
        RECT 231.520 -203.420 231.890 -203.390 ;
        RECT 229.460 -203.425 231.890 -203.420 ;
        RECT 226.715 -203.595 231.890 -203.425 ;
        RECT 233.675 -203.530 233.980 -201.495 ;
        RECT 226.720 -203.615 231.890 -203.595 ;
        RECT 226.720 -203.625 229.465 -203.615 ;
        RECT 224.655 -203.765 225.020 -203.735 ;
        RECT 231.520 -203.745 231.890 -203.615 ;
        RECT 223.760 -203.850 225.020 -203.765 ;
        RECT 223.785 -203.970 225.020 -203.850 ;
        RECT 229.195 -203.905 229.870 -203.865 ;
        RECT 229.095 -203.915 229.870 -203.905 ;
        RECT 223.785 -204.055 224.435 -203.970 ;
        RECT 224.655 -204.035 225.020 -203.970 ;
        RECT 228.060 -204.095 229.870 -203.915 ;
        RECT 232.455 -203.960 236.380 -203.530 ;
        RECT 229.095 -204.105 229.870 -204.095 ;
        RECT 229.195 -204.135 229.870 -204.105 ;
        RECT 230.110 -204.020 232.205 -203.980 ;
        RECT 230.110 -204.170 232.260 -204.020 ;
        RECT 225.245 -205.245 225.415 -204.205 ;
        RECT 226.225 -205.245 226.395 -204.205 ;
        RECT 227.205 -205.245 227.375 -204.205 ;
        RECT 230.110 -205.890 230.280 -204.170 ;
        RECT 231.090 -205.890 231.260 -204.170 ;
        RECT 231.955 -204.915 232.260 -204.170 ;
        RECT 233.155 -204.740 233.325 -203.960 ;
        RECT 233.645 -204.740 233.815 -204.200 ;
        RECT 234.135 -204.740 234.305 -203.960 ;
        RECT 234.625 -204.740 234.795 -204.200 ;
        RECT 232.565 -204.915 232.930 -204.885 ;
        RECT 231.955 -204.980 232.930 -204.915 ;
        RECT 232.065 -205.120 232.930 -204.980 ;
        RECT 232.565 -205.185 232.930 -205.120 ;
        RECT 235.115 -205.035 236.975 -204.685 ;
        RECT 233.155 -205.895 233.325 -205.355 ;
        RECT 234.135 -205.895 234.305 -205.355 ;
        RECT 235.115 -205.895 235.285 -205.035 ;
        RECT 233.385 -208.235 234.585 -208.065 ;
        RECT 225.115 -210.570 225.285 -208.850 ;
        RECT 226.095 -210.570 226.265 -208.850 ;
        RECT 228.160 -209.385 228.330 -208.845 ;
        RECT 229.140 -209.385 229.310 -208.845 ;
        RECT 227.570 -209.620 227.935 -209.555 ;
        RECT 227.070 -209.760 227.935 -209.620 ;
        RECT 226.960 -209.825 227.935 -209.760 ;
        RECT 226.960 -210.570 227.265 -209.825 ;
        RECT 227.570 -209.855 227.935 -209.825 ;
        RECT 230.120 -209.705 230.290 -208.845 ;
        RECT 225.115 -210.720 227.265 -210.570 ;
        RECT 225.115 -210.760 227.210 -210.720 ;
        RECT 228.160 -210.780 228.330 -210.000 ;
        RECT 228.650 -210.540 228.820 -210.000 ;
        RECT 229.140 -210.780 229.310 -210.000 ;
        RECT 229.630 -210.540 229.800 -210.000 ;
        RECT 230.120 -210.055 231.510 -209.705 ;
        RECT 223.335 -211.125 224.470 -211.115 ;
        RECT 226.525 -211.125 226.895 -210.995 ;
        RECT 223.335 -211.315 226.895 -211.125 ;
        RECT 227.460 -211.210 230.535 -210.780 ;
        RECT 224.465 -211.320 226.895 -211.315 ;
        RECT 224.465 -211.325 224.820 -211.320 ;
        RECT 226.525 -211.350 226.895 -211.320 ;
        RECT 224.625 -213.075 224.795 -211.535 ;
        RECT 225.115 -213.075 225.285 -211.535 ;
        RECT 225.605 -213.075 225.775 -211.535 ;
        RECT 226.095 -213.075 226.265 -211.535 ;
        RECT 226.585 -213.075 226.755 -211.535 ;
        RECT 225.110 -213.335 225.285 -213.075 ;
        RECT 228.680 -213.245 228.985 -211.210 ;
        RECT 231.130 -212.030 231.480 -210.055 ;
        RECT 232.350 -211.325 232.520 -208.405 ;
        RECT 233.385 -208.445 233.595 -208.235 ;
        RECT 232.330 -211.620 232.540 -211.325 ;
        RECT 233.405 -211.355 233.575 -208.445 ;
        RECT 233.895 -211.345 234.065 -208.405 ;
        RECT 234.375 -208.455 234.585 -208.235 ;
        RECT 233.390 -211.620 233.600 -211.355 ;
        RECT 232.330 -211.800 233.600 -211.620 ;
        RECT 233.875 -211.615 234.085 -211.345 ;
        RECT 234.385 -211.445 234.555 -208.455 ;
        RECT 235.445 -211.375 235.615 -208.405 ;
        RECT 233.875 -211.810 234.580 -211.615 ;
        RECT 234.365 -211.870 234.580 -211.810 ;
        RECT 233.155 -212.030 233.930 -211.980 ;
        RECT 231.130 -212.210 233.930 -212.030 ;
        RECT 231.130 -212.220 231.480 -212.210 ;
        RECT 233.155 -212.255 233.930 -212.210 ;
        RECT 234.365 -212.145 235.270 -211.870 ;
        RECT 234.365 -212.495 234.580 -212.145 ;
        RECT 231.805 -212.565 232.580 -212.520 ;
        RECT 231.620 -212.735 232.580 -212.565 ;
        RECT 231.805 -212.795 232.580 -212.735 ;
        RECT 232.810 -212.695 234.580 -212.495 ;
        RECT 235.440 -212.595 235.655 -211.375 ;
        RECT 236.625 -211.720 236.975 -205.035 ;
        RECT 237.965 -211.350 238.180 -201.475 ;
        RECT 239.600 -203.590 239.980 -200.070 ;
        RECT 241.110 -199.850 250.045 -199.660 ;
        RECT 265.865 -199.040 269.800 -198.235 ;
        RECT 241.110 -201.740 241.300 -199.850 ;
        RECT 247.145 -201.345 250.470 -201.205 ;
        RECT 247.145 -201.635 252.320 -201.345 ;
        RECT 240.995 -202.010 241.360 -201.740 ;
        RECT 247.145 -202.040 247.575 -201.635 ;
        RECT 248.445 -201.820 248.620 -201.635 ;
        RECT 250.070 -201.650 252.320 -201.635 ;
        RECT 242.885 -202.470 247.575 -202.040 ;
        RECT 242.125 -203.590 242.775 -203.460 ;
        RECT 239.600 -203.920 242.775 -203.590 ;
        RECT 243.585 -203.750 243.755 -202.470 ;
        RECT 244.075 -203.750 244.245 -202.710 ;
        RECT 244.565 -203.750 244.735 -202.470 ;
        RECT 245.055 -203.580 245.225 -202.710 ;
        RECT 247.960 -203.360 248.130 -201.820 ;
        RECT 248.450 -203.360 248.620 -201.820 ;
        RECT 248.940 -203.360 249.110 -201.820 ;
        RECT 249.430 -203.360 249.600 -201.820 ;
        RECT 249.920 -203.360 250.090 -201.820 ;
        RECT 247.800 -203.575 248.155 -203.570 ;
        RECT 249.860 -203.575 250.230 -203.545 ;
        RECT 247.800 -203.580 250.230 -203.575 ;
        RECT 245.055 -203.750 250.230 -203.580 ;
        RECT 252.015 -203.685 252.320 -201.650 ;
        RECT 245.060 -203.770 250.230 -203.750 ;
        RECT 245.060 -203.780 247.805 -203.770 ;
        RECT 242.995 -203.920 243.360 -203.890 ;
        RECT 249.860 -203.900 250.230 -203.770 ;
        RECT 239.600 -203.970 243.360 -203.920 ;
        RECT 242.125 -204.125 243.360 -203.970 ;
        RECT 247.535 -204.060 248.210 -204.020 ;
        RECT 247.435 -204.070 248.210 -204.060 ;
        RECT 242.125 -204.210 242.775 -204.125 ;
        RECT 242.995 -204.190 243.360 -204.125 ;
        RECT 242.260 -204.460 242.640 -204.210 ;
        RECT 246.400 -204.250 248.210 -204.070 ;
        RECT 250.795 -204.115 254.720 -203.685 ;
        RECT 247.435 -204.260 248.210 -204.250 ;
        RECT 247.535 -204.290 248.210 -204.260 ;
        RECT 248.450 -204.175 250.545 -204.135 ;
        RECT 248.450 -204.325 250.600 -204.175 ;
        RECT 243.585 -205.400 243.755 -204.360 ;
        RECT 244.565 -205.400 244.735 -204.360 ;
        RECT 245.545 -205.400 245.715 -204.360 ;
        RECT 248.450 -206.045 248.620 -204.325 ;
        RECT 249.430 -206.045 249.600 -204.325 ;
        RECT 250.295 -205.070 250.600 -204.325 ;
        RECT 251.495 -204.895 251.665 -204.115 ;
        RECT 251.985 -204.895 252.155 -204.355 ;
        RECT 252.475 -204.895 252.645 -204.115 ;
        RECT 252.965 -204.895 253.135 -204.355 ;
        RECT 250.905 -205.070 251.270 -205.040 ;
        RECT 250.295 -205.135 251.270 -205.070 ;
        RECT 250.405 -205.275 251.270 -205.135 ;
        RECT 250.905 -205.340 251.270 -205.275 ;
        RECT 253.455 -205.190 255.315 -204.840 ;
        RECT 251.495 -206.050 251.665 -205.510 ;
        RECT 252.475 -206.050 252.645 -205.510 ;
        RECT 253.455 -206.050 253.625 -205.190 ;
        RECT 251.725 -208.390 252.925 -208.220 ;
        RECT 243.455 -210.725 243.625 -209.005 ;
        RECT 244.435 -210.725 244.605 -209.005 ;
        RECT 246.500 -209.540 246.670 -209.000 ;
        RECT 247.480 -209.540 247.650 -209.000 ;
        RECT 245.910 -209.775 246.275 -209.710 ;
        RECT 245.410 -209.915 246.275 -209.775 ;
        RECT 245.300 -209.980 246.275 -209.915 ;
        RECT 245.300 -210.725 245.605 -209.980 ;
        RECT 245.910 -210.010 246.275 -209.980 ;
        RECT 248.460 -209.860 248.630 -209.000 ;
        RECT 243.455 -210.875 245.605 -210.725 ;
        RECT 243.455 -210.915 245.550 -210.875 ;
        RECT 246.500 -210.935 246.670 -210.155 ;
        RECT 246.990 -210.695 247.160 -210.155 ;
        RECT 247.480 -210.935 247.650 -210.155 ;
        RECT 247.970 -210.695 248.140 -210.155 ;
        RECT 248.460 -210.210 249.850 -209.860 ;
        RECT 241.675 -211.280 242.810 -211.270 ;
        RECT 244.865 -211.280 245.235 -211.150 ;
        RECT 237.965 -211.565 239.390 -211.350 ;
        RECT 241.675 -211.470 245.235 -211.280 ;
        RECT 245.800 -211.365 248.875 -210.935 ;
        RECT 242.805 -211.475 245.235 -211.470 ;
        RECT 242.805 -211.480 243.160 -211.475 ;
        RECT 244.865 -211.505 245.235 -211.475 ;
        RECT 236.570 -212.080 237.095 -211.720 ;
        RECT 239.175 -212.595 239.390 -211.565 ;
        RECT 226.735 -213.335 228.985 -213.245 ;
        RECT 224.525 -213.550 228.985 -213.335 ;
        RECT 224.525 -213.640 226.770 -213.550 ;
        RECT 228.680 -215.025 228.985 -213.550 ;
        RECT 232.350 -214.435 232.520 -212.965 ;
        RECT 232.810 -213.045 233.035 -212.695 ;
        RECT 234.770 -212.795 239.390 -212.595 ;
        RECT 235.010 -212.810 239.390 -212.795 ;
        RECT 232.315 -215.025 232.550 -214.435 ;
        RECT 232.840 -214.505 233.010 -213.045 ;
        RECT 233.330 -214.430 233.500 -212.965 ;
        RECT 234.540 -214.380 234.710 -212.965 ;
        RECT 235.010 -213.010 235.230 -212.810 ;
        RECT 233.295 -215.025 233.530 -214.430 ;
        RECT 234.505 -215.025 234.740 -214.380 ;
        RECT 235.030 -214.505 235.200 -213.010 ;
        RECT 242.965 -213.230 243.135 -211.690 ;
        RECT 243.455 -213.230 243.625 -211.690 ;
        RECT 243.945 -213.230 244.115 -211.690 ;
        RECT 244.435 -213.230 244.605 -211.690 ;
        RECT 244.925 -213.230 245.095 -211.690 ;
        RECT 243.450 -213.490 243.625 -213.230 ;
        RECT 247.020 -213.400 247.325 -211.365 ;
        RECT 249.470 -212.185 249.820 -210.210 ;
        RECT 250.690 -211.480 250.860 -208.560 ;
        RECT 251.725 -208.600 251.935 -208.390 ;
        RECT 250.670 -211.775 250.880 -211.480 ;
        RECT 251.745 -211.510 251.915 -208.600 ;
        RECT 252.235 -211.500 252.405 -208.560 ;
        RECT 252.715 -208.610 252.925 -208.390 ;
        RECT 251.730 -211.775 251.940 -211.510 ;
        RECT 250.670 -211.955 251.940 -211.775 ;
        RECT 252.215 -211.770 252.425 -211.500 ;
        RECT 252.725 -211.600 252.895 -208.610 ;
        RECT 253.785 -211.530 253.955 -208.560 ;
        RECT 252.215 -211.965 252.920 -211.770 ;
        RECT 252.705 -212.025 252.920 -211.965 ;
        RECT 251.495 -212.185 252.270 -212.135 ;
        RECT 249.470 -212.365 252.270 -212.185 ;
        RECT 249.470 -212.375 249.820 -212.365 ;
        RECT 251.495 -212.410 252.270 -212.365 ;
        RECT 252.705 -212.300 253.610 -212.025 ;
        RECT 252.705 -212.650 252.920 -212.300 ;
        RECT 250.145 -212.720 250.920 -212.675 ;
        RECT 249.960 -212.890 250.920 -212.720 ;
        RECT 250.145 -212.950 250.920 -212.890 ;
        RECT 251.150 -212.850 252.920 -212.650 ;
        RECT 253.780 -212.750 253.995 -211.530 ;
        RECT 254.965 -211.875 255.315 -205.190 ;
        RECT 254.910 -212.235 255.435 -211.875 ;
        RECT 257.560 -212.750 258.630 -212.175 ;
        RECT 245.075 -213.490 247.325 -213.400 ;
        RECT 242.865 -213.705 247.325 -213.490 ;
        RECT 242.865 -213.795 245.110 -213.705 ;
        RECT 228.680 -215.590 236.065 -215.025 ;
        RECT 247.020 -215.180 247.325 -213.705 ;
        RECT 250.690 -214.590 250.860 -213.120 ;
        RECT 251.150 -213.200 251.375 -212.850 ;
        RECT 253.110 -212.950 259.120 -212.750 ;
        RECT 253.350 -212.965 259.120 -212.950 ;
        RECT 250.655 -215.180 250.890 -214.590 ;
        RECT 251.180 -214.660 251.350 -213.200 ;
        RECT 251.670 -214.585 251.840 -213.120 ;
        RECT 252.880 -214.535 253.050 -213.120 ;
        RECT 253.350 -213.165 253.570 -212.965 ;
        RECT 251.635 -215.180 251.870 -214.585 ;
        RECT 252.845 -215.180 253.080 -214.535 ;
        RECT 253.370 -214.660 253.540 -213.165 ;
        RECT 257.560 -213.275 258.630 -212.965 ;
        RECT 247.020 -215.745 254.405 -215.180 ;
        RECT 265.865 -218.645 266.670 -199.040 ;
        RECT 269.420 -199.520 269.800 -199.040 ;
        RECT 295.845 -199.490 296.035 -195.015 ;
        RECT 313.190 -198.370 313.570 -193.550 ;
        RECT 314.265 -193.555 316.695 -193.550 ;
        RECT 314.265 -193.560 314.620 -193.555 ;
        RECT 316.325 -193.585 316.695 -193.555 ;
        RECT 314.425 -195.310 314.595 -193.770 ;
        RECT 314.915 -195.310 315.085 -193.770 ;
        RECT 315.405 -195.310 315.575 -193.770 ;
        RECT 315.895 -195.310 316.065 -193.770 ;
        RECT 316.385 -195.310 316.555 -193.770 ;
        RECT 314.910 -195.570 315.085 -195.310 ;
        RECT 318.480 -195.480 318.785 -193.445 ;
        RECT 320.930 -194.265 321.280 -192.290 ;
        RECT 322.150 -193.560 322.320 -190.640 ;
        RECT 323.185 -190.680 323.395 -190.470 ;
        RECT 322.130 -193.855 322.340 -193.560 ;
        RECT 323.205 -193.590 323.375 -190.680 ;
        RECT 323.695 -193.580 323.865 -190.640 ;
        RECT 324.175 -190.690 324.385 -190.470 ;
        RECT 323.190 -193.855 323.400 -193.590 ;
        RECT 322.130 -194.035 323.400 -193.855 ;
        RECT 323.675 -193.850 323.885 -193.580 ;
        RECT 324.185 -193.680 324.355 -190.690 ;
        RECT 325.245 -193.610 325.415 -190.640 ;
        RECT 323.675 -194.045 324.380 -193.850 ;
        RECT 324.165 -194.105 324.380 -194.045 ;
        RECT 322.955 -194.265 323.730 -194.215 ;
        RECT 320.930 -194.445 323.730 -194.265 ;
        RECT 320.930 -194.455 321.280 -194.445 ;
        RECT 322.955 -194.490 323.730 -194.445 ;
        RECT 324.165 -194.380 325.070 -194.105 ;
        RECT 324.165 -194.730 324.380 -194.380 ;
        RECT 321.605 -194.800 322.380 -194.755 ;
        RECT 321.420 -194.970 322.380 -194.800 ;
        RECT 321.605 -195.030 322.380 -194.970 ;
        RECT 322.610 -194.930 324.380 -194.730 ;
        RECT 325.240 -194.830 325.455 -193.610 ;
        RECT 326.425 -193.955 326.775 -187.270 ;
        RECT 360.810 -187.395 360.980 -186.355 ;
        RECT 361.790 -187.395 361.960 -186.355 ;
        RECT 362.770 -187.395 362.940 -186.355 ;
        RECT 365.675 -188.040 365.845 -186.320 ;
        RECT 366.655 -188.040 366.825 -186.320 ;
        RECT 367.520 -187.065 367.825 -186.320 ;
        RECT 368.720 -186.890 368.890 -186.110 ;
        RECT 369.210 -186.890 369.380 -186.350 ;
        RECT 369.700 -186.890 369.870 -186.110 ;
        RECT 412.495 -186.130 414.645 -185.980 ;
        RECT 370.190 -186.890 370.360 -186.350 ;
        RECT 368.130 -187.065 368.495 -187.035 ;
        RECT 367.520 -187.130 368.495 -187.065 ;
        RECT 367.630 -187.270 368.495 -187.130 ;
        RECT 368.130 -187.335 368.495 -187.270 ;
        RECT 370.680 -187.185 372.540 -186.835 ;
        RECT 368.720 -188.045 368.890 -187.505 ;
        RECT 369.700 -188.045 369.870 -187.505 ;
        RECT 370.680 -188.045 370.850 -187.185 ;
        RECT 333.005 -189.750 334.610 -189.580 ;
        RECT 332.110 -192.430 332.280 -189.930 ;
        RECT 332.105 -192.660 332.280 -192.430 ;
        RECT 333.005 -192.660 333.205 -189.750 ;
        RECT 333.450 -189.950 333.625 -189.750 ;
        RECT 333.455 -192.470 333.625 -189.950 ;
        RECT 333.945 -192.435 334.115 -189.930 ;
        RECT 334.435 -189.945 334.610 -189.750 ;
        RECT 332.105 -192.860 333.205 -192.660 ;
        RECT 333.930 -193.035 334.120 -192.435 ;
        RECT 334.435 -192.470 334.605 -189.945 ;
        RECT 335.085 -192.850 335.255 -189.930 ;
        RECT 336.715 -192.500 336.885 -189.930 ;
        RECT 337.855 -191.380 338.025 -189.930 ;
        RECT 368.950 -190.385 370.150 -190.215 ;
        RECT 337.850 -191.845 338.035 -191.380 ;
        RECT 337.850 -192.030 338.535 -191.845 ;
        RECT 336.715 -192.670 337.510 -192.500 ;
        RECT 335.830 -192.850 336.520 -192.795 ;
        RECT 332.110 -193.225 334.120 -193.035 ;
        RECT 334.455 -193.020 336.520 -192.850 ;
        RECT 330.925 -193.280 331.615 -193.230 ;
        RECT 328.975 -193.450 331.615 -193.280 ;
        RECT 326.370 -194.315 326.895 -193.955 ;
        RECT 328.975 -194.830 329.190 -193.450 ;
        RECT 330.925 -193.500 331.615 -193.450 ;
        RECT 331.205 -193.955 331.895 -193.910 ;
        RECT 330.155 -194.125 331.895 -193.955 ;
        RECT 330.155 -194.760 330.515 -194.125 ;
        RECT 331.205 -194.180 331.895 -194.125 ;
        RECT 330.155 -194.805 330.575 -194.760 ;
        RECT 316.535 -195.570 318.785 -195.480 ;
        RECT 314.325 -195.785 318.785 -195.570 ;
        RECT 314.325 -195.875 316.570 -195.785 ;
        RECT 318.480 -197.260 318.785 -195.785 ;
        RECT 322.150 -196.670 322.320 -195.200 ;
        RECT 322.610 -195.280 322.835 -194.930 ;
        RECT 324.570 -195.030 329.190 -194.830 ;
        RECT 324.810 -195.045 329.190 -195.030 ;
        RECT 322.115 -197.260 322.350 -196.670 ;
        RECT 322.640 -196.740 322.810 -195.280 ;
        RECT 323.130 -196.665 323.300 -195.200 ;
        RECT 324.340 -196.615 324.510 -195.200 ;
        RECT 324.810 -195.245 325.030 -195.045 ;
        RECT 330.180 -195.155 330.575 -194.805 ;
        RECT 323.095 -197.260 323.330 -196.665 ;
        RECT 324.305 -197.260 324.540 -196.615 ;
        RECT 324.830 -196.740 325.000 -195.245 ;
        RECT 331.620 -196.365 331.790 -194.910 ;
        RECT 331.610 -196.920 331.795 -196.365 ;
        RECT 332.110 -196.450 332.280 -193.225 ;
        RECT 333.255 -193.575 333.445 -193.225 ;
        RECT 334.455 -193.415 334.625 -193.020 ;
        RECT 335.830 -193.065 336.520 -193.020 ;
        RECT 333.205 -194.265 333.475 -193.575 ;
        RECT 333.970 -193.585 334.625 -193.415 ;
        RECT 334.955 -193.500 335.645 -193.230 ;
        RECT 336.880 -193.575 337.150 -192.885 ;
        RECT 337.340 -192.890 337.510 -192.670 ;
        RECT 337.340 -193.160 338.170 -192.890 ;
        RECT 333.970 -196.450 334.140 -193.585 ;
        RECT 337.340 -193.735 337.510 -193.160 ;
        RECT 337.770 -193.735 338.040 -193.650 ;
        RECT 334.460 -193.930 335.255 -193.755 ;
        RECT 337.340 -193.760 338.040 -193.735 ;
        RECT 337.200 -193.905 338.040 -193.760 ;
        RECT 334.460 -196.450 334.630 -193.930 ;
        RECT 335.085 -196.450 335.255 -193.930 ;
        RECT 335.575 -196.365 335.745 -193.910 ;
        RECT 336.225 -196.360 336.395 -193.910 ;
        RECT 328.925 -196.940 331.980 -196.920 ;
        RECT 335.570 -196.940 335.755 -196.365 ;
        RECT 336.210 -196.940 336.395 -196.360 ;
        RECT 336.715 -196.450 336.885 -193.910 ;
        RECT 337.200 -193.930 337.510 -193.905 ;
        RECT 337.205 -196.450 337.375 -193.930 ;
        RECT 337.770 -193.945 338.040 -193.905 ;
        RECT 338.345 -194.495 338.535 -192.030 ;
        RECT 360.680 -192.720 360.850 -191.000 ;
        RECT 361.660 -192.720 361.830 -191.000 ;
        RECT 363.725 -191.535 363.895 -190.995 ;
        RECT 364.705 -191.535 364.875 -190.995 ;
        RECT 363.135 -191.770 363.500 -191.705 ;
        RECT 362.635 -191.910 363.500 -191.770 ;
        RECT 362.525 -191.975 363.500 -191.910 ;
        RECT 362.525 -192.720 362.830 -191.975 ;
        RECT 363.135 -192.005 363.500 -191.975 ;
        RECT 365.685 -191.855 365.855 -190.995 ;
        RECT 360.680 -192.870 362.830 -192.720 ;
        RECT 360.680 -192.910 362.775 -192.870 ;
        RECT 363.725 -192.930 363.895 -192.150 ;
        RECT 364.215 -192.690 364.385 -192.150 ;
        RECT 364.705 -192.930 364.875 -192.150 ;
        RECT 365.195 -192.690 365.365 -192.150 ;
        RECT 365.685 -192.205 367.075 -191.855 ;
        RECT 358.900 -193.275 360.035 -193.265 ;
        RECT 362.090 -193.275 362.460 -193.145 ;
        RECT 358.900 -193.465 362.460 -193.275 ;
        RECT 363.025 -193.360 366.100 -192.930 ;
        RECT 338.345 -194.685 339.805 -194.495 ;
        RECT 337.855 -196.355 338.025 -194.910 ;
        RECT 338.345 -194.935 338.535 -194.685 ;
        RECT 337.845 -196.940 338.030 -196.355 ;
        RECT 338.345 -196.450 338.515 -194.935 ;
        RECT 328.925 -197.260 338.595 -196.940 ;
        RECT 318.480 -197.485 338.595 -197.260 ;
        RECT 318.480 -197.825 329.490 -197.485 ;
        RECT 331.230 -197.745 338.595 -197.485 ;
        RECT 269.420 -199.900 285.970 -199.520 ;
        RECT 269.420 -200.810 269.800 -199.900 ;
        RECT 269.420 -201.190 270.130 -200.810 ;
        RECT 269.750 -203.135 270.130 -201.190 ;
        RECT 274.795 -201.020 278.120 -200.880 ;
        RECT 274.795 -201.310 279.970 -201.020 ;
        RECT 283.840 -201.305 284.300 -200.880 ;
        RECT 274.795 -201.715 275.225 -201.310 ;
        RECT 276.095 -201.495 276.270 -201.310 ;
        RECT 277.720 -201.325 279.970 -201.310 ;
        RECT 270.535 -202.145 275.225 -201.715 ;
        RECT 269.750 -203.595 270.425 -203.135 ;
        RECT 271.235 -203.425 271.405 -202.145 ;
        RECT 271.725 -203.425 271.895 -202.385 ;
        RECT 272.215 -203.425 272.385 -202.145 ;
        RECT 272.705 -203.255 272.875 -202.385 ;
        RECT 275.610 -203.035 275.780 -201.495 ;
        RECT 276.100 -203.035 276.270 -201.495 ;
        RECT 276.590 -203.035 276.760 -201.495 ;
        RECT 277.080 -203.035 277.250 -201.495 ;
        RECT 277.570 -203.035 277.740 -201.495 ;
        RECT 275.450 -203.250 275.805 -203.245 ;
        RECT 277.510 -203.250 277.880 -203.220 ;
        RECT 275.450 -203.255 277.880 -203.250 ;
        RECT 272.705 -203.425 277.880 -203.255 ;
        RECT 279.665 -203.360 279.970 -201.325 ;
        RECT 272.710 -203.445 277.880 -203.425 ;
        RECT 272.710 -203.455 275.455 -203.445 ;
        RECT 270.645 -203.595 271.010 -203.565 ;
        RECT 277.510 -203.575 277.880 -203.445 ;
        RECT 269.750 -203.680 271.010 -203.595 ;
        RECT 269.775 -203.800 271.010 -203.680 ;
        RECT 275.185 -203.735 275.860 -203.695 ;
        RECT 275.085 -203.745 275.860 -203.735 ;
        RECT 269.775 -203.885 270.425 -203.800 ;
        RECT 270.645 -203.865 271.010 -203.800 ;
        RECT 274.050 -203.925 275.860 -203.745 ;
        RECT 278.445 -203.790 282.370 -203.360 ;
        RECT 275.085 -203.935 275.860 -203.925 ;
        RECT 275.185 -203.965 275.860 -203.935 ;
        RECT 276.100 -203.850 278.195 -203.810 ;
        RECT 276.100 -204.000 278.250 -203.850 ;
        RECT 271.235 -205.075 271.405 -204.035 ;
        RECT 272.215 -205.075 272.385 -204.035 ;
        RECT 273.195 -205.075 273.365 -204.035 ;
        RECT 276.100 -205.720 276.270 -204.000 ;
        RECT 277.080 -205.720 277.250 -204.000 ;
        RECT 277.945 -204.745 278.250 -204.000 ;
        RECT 279.145 -204.570 279.315 -203.790 ;
        RECT 279.635 -204.570 279.805 -204.030 ;
        RECT 280.125 -204.570 280.295 -203.790 ;
        RECT 280.615 -204.570 280.785 -204.030 ;
        RECT 278.555 -204.745 278.920 -204.715 ;
        RECT 277.945 -204.810 278.920 -204.745 ;
        RECT 278.055 -204.950 278.920 -204.810 ;
        RECT 278.555 -205.015 278.920 -204.950 ;
        RECT 281.105 -204.865 282.965 -204.515 ;
        RECT 279.145 -205.725 279.315 -205.185 ;
        RECT 280.125 -205.725 280.295 -205.185 ;
        RECT 281.105 -205.725 281.275 -204.865 ;
        RECT 279.375 -208.065 280.575 -207.895 ;
        RECT 271.105 -210.400 271.275 -208.680 ;
        RECT 272.085 -210.400 272.255 -208.680 ;
        RECT 274.150 -209.215 274.320 -208.675 ;
        RECT 275.130 -209.215 275.300 -208.675 ;
        RECT 273.560 -209.450 273.925 -209.385 ;
        RECT 273.060 -209.590 273.925 -209.450 ;
        RECT 272.950 -209.655 273.925 -209.590 ;
        RECT 272.950 -210.400 273.255 -209.655 ;
        RECT 273.560 -209.685 273.925 -209.655 ;
        RECT 276.110 -209.535 276.280 -208.675 ;
        RECT 271.105 -210.550 273.255 -210.400 ;
        RECT 271.105 -210.590 273.200 -210.550 ;
        RECT 274.150 -210.610 274.320 -209.830 ;
        RECT 274.640 -210.370 274.810 -209.830 ;
        RECT 275.130 -210.610 275.300 -209.830 ;
        RECT 275.620 -210.370 275.790 -209.830 ;
        RECT 276.110 -209.885 277.500 -209.535 ;
        RECT 269.325 -210.955 270.460 -210.945 ;
        RECT 272.515 -210.955 272.885 -210.825 ;
        RECT 269.325 -211.145 272.885 -210.955 ;
        RECT 273.450 -211.040 276.525 -210.610 ;
        RECT 270.455 -211.150 272.885 -211.145 ;
        RECT 270.455 -211.155 270.810 -211.150 ;
        RECT 272.515 -211.180 272.885 -211.150 ;
        RECT 270.615 -212.905 270.785 -211.365 ;
        RECT 271.105 -212.905 271.275 -211.365 ;
        RECT 271.595 -212.905 271.765 -211.365 ;
        RECT 272.085 -212.905 272.255 -211.365 ;
        RECT 272.575 -212.905 272.745 -211.365 ;
        RECT 271.100 -213.165 271.275 -212.905 ;
        RECT 274.670 -213.075 274.975 -211.040 ;
        RECT 277.120 -211.860 277.470 -209.885 ;
        RECT 278.340 -211.155 278.510 -208.235 ;
        RECT 279.375 -208.275 279.585 -208.065 ;
        RECT 278.320 -211.450 278.530 -211.155 ;
        RECT 279.395 -211.185 279.565 -208.275 ;
        RECT 279.885 -211.175 280.055 -208.235 ;
        RECT 280.365 -208.285 280.575 -208.065 ;
        RECT 279.380 -211.450 279.590 -211.185 ;
        RECT 278.320 -211.630 279.590 -211.450 ;
        RECT 279.865 -211.445 280.075 -211.175 ;
        RECT 280.375 -211.275 280.545 -208.285 ;
        RECT 281.435 -211.205 281.605 -208.235 ;
        RECT 279.865 -211.640 280.570 -211.445 ;
        RECT 280.355 -211.700 280.570 -211.640 ;
        RECT 279.145 -211.860 279.920 -211.810 ;
        RECT 277.120 -212.040 279.920 -211.860 ;
        RECT 277.120 -212.050 277.470 -212.040 ;
        RECT 279.145 -212.085 279.920 -212.040 ;
        RECT 280.355 -211.975 281.260 -211.700 ;
        RECT 280.355 -212.325 280.570 -211.975 ;
        RECT 277.795 -212.395 278.570 -212.350 ;
        RECT 277.610 -212.565 278.570 -212.395 ;
        RECT 277.795 -212.625 278.570 -212.565 ;
        RECT 278.800 -212.525 280.570 -212.325 ;
        RECT 281.430 -212.425 281.645 -211.205 ;
        RECT 282.615 -211.550 282.965 -204.865 ;
        RECT 283.955 -211.180 284.170 -201.305 ;
        RECT 285.590 -203.420 285.970 -199.900 ;
        RECT 287.100 -199.680 296.035 -199.490 ;
        RECT 309.625 -199.190 313.570 -198.370 ;
        RECT 339.615 -199.160 339.805 -194.685 ;
        RECT 358.955 -198.575 359.335 -193.465 ;
        RECT 360.030 -193.470 362.460 -193.465 ;
        RECT 360.030 -193.475 360.385 -193.470 ;
        RECT 362.090 -193.500 362.460 -193.470 ;
        RECT 360.190 -195.225 360.360 -193.685 ;
        RECT 360.680 -195.225 360.850 -193.685 ;
        RECT 361.170 -195.225 361.340 -193.685 ;
        RECT 361.660 -195.225 361.830 -193.685 ;
        RECT 362.150 -195.225 362.320 -193.685 ;
        RECT 360.675 -195.485 360.850 -195.225 ;
        RECT 364.245 -195.395 364.550 -193.360 ;
        RECT 366.695 -194.180 367.045 -192.205 ;
        RECT 367.915 -193.475 368.085 -190.555 ;
        RECT 368.950 -190.595 369.160 -190.385 ;
        RECT 367.895 -193.770 368.105 -193.475 ;
        RECT 368.970 -193.505 369.140 -190.595 ;
        RECT 369.460 -193.495 369.630 -190.555 ;
        RECT 369.940 -190.605 370.150 -190.385 ;
        RECT 368.955 -193.770 369.165 -193.505 ;
        RECT 367.895 -193.950 369.165 -193.770 ;
        RECT 369.440 -193.765 369.650 -193.495 ;
        RECT 369.950 -193.595 370.120 -190.605 ;
        RECT 371.010 -193.525 371.180 -190.555 ;
        RECT 369.440 -193.960 370.145 -193.765 ;
        RECT 369.930 -194.020 370.145 -193.960 ;
        RECT 368.720 -194.180 369.495 -194.130 ;
        RECT 366.695 -194.360 369.495 -194.180 ;
        RECT 366.695 -194.370 367.045 -194.360 ;
        RECT 368.720 -194.405 369.495 -194.360 ;
        RECT 369.930 -194.295 370.835 -194.020 ;
        RECT 369.930 -194.645 370.145 -194.295 ;
        RECT 367.370 -194.715 368.145 -194.670 ;
        RECT 367.185 -194.885 368.145 -194.715 ;
        RECT 367.370 -194.945 368.145 -194.885 ;
        RECT 368.375 -194.845 370.145 -194.645 ;
        RECT 371.005 -194.745 371.220 -193.525 ;
        RECT 372.190 -193.870 372.540 -187.185 ;
        RECT 407.630 -187.205 407.800 -186.165 ;
        RECT 408.610 -187.205 408.780 -186.165 ;
        RECT 409.590 -187.205 409.760 -186.165 ;
        RECT 412.495 -187.850 412.665 -186.130 ;
        RECT 413.475 -187.850 413.645 -186.130 ;
        RECT 414.340 -186.875 414.645 -186.130 ;
        RECT 415.540 -186.700 415.710 -185.920 ;
        RECT 416.030 -186.700 416.200 -186.160 ;
        RECT 416.520 -186.700 416.690 -185.920 ;
        RECT 417.010 -186.700 417.180 -186.160 ;
        RECT 414.950 -186.875 415.315 -186.845 ;
        RECT 414.340 -186.940 415.315 -186.875 ;
        RECT 414.450 -187.080 415.315 -186.940 ;
        RECT 414.950 -187.145 415.315 -187.080 ;
        RECT 417.500 -186.995 419.360 -186.645 ;
        RECT 415.540 -187.855 415.710 -187.315 ;
        RECT 416.520 -187.855 416.690 -187.315 ;
        RECT 417.500 -187.855 417.670 -186.995 ;
        RECT 378.770 -189.665 380.375 -189.495 ;
        RECT 377.875 -192.345 378.045 -189.845 ;
        RECT 377.870 -192.575 378.045 -192.345 ;
        RECT 378.770 -192.575 378.970 -189.665 ;
        RECT 379.215 -189.865 379.390 -189.665 ;
        RECT 379.220 -192.385 379.390 -189.865 ;
        RECT 379.710 -192.350 379.880 -189.845 ;
        RECT 380.200 -189.860 380.375 -189.665 ;
        RECT 377.870 -192.775 378.970 -192.575 ;
        RECT 379.695 -192.950 379.885 -192.350 ;
        RECT 380.200 -192.385 380.370 -189.860 ;
        RECT 380.850 -192.765 381.020 -189.845 ;
        RECT 382.480 -192.415 382.650 -189.845 ;
        RECT 383.620 -191.295 383.790 -189.845 ;
        RECT 415.770 -190.195 416.970 -190.025 ;
        RECT 383.615 -191.760 383.800 -191.295 ;
        RECT 383.615 -191.945 384.300 -191.760 ;
        RECT 382.480 -192.585 383.275 -192.415 ;
        RECT 381.595 -192.765 382.285 -192.710 ;
        RECT 377.875 -193.140 379.885 -192.950 ;
        RECT 380.220 -192.935 382.285 -192.765 ;
        RECT 376.690 -193.195 377.380 -193.145 ;
        RECT 374.740 -193.365 377.380 -193.195 ;
        RECT 372.135 -194.230 372.660 -193.870 ;
        RECT 374.740 -194.745 374.955 -193.365 ;
        RECT 376.690 -193.415 377.380 -193.365 ;
        RECT 376.970 -193.870 377.660 -193.825 ;
        RECT 375.920 -194.040 377.660 -193.870 ;
        RECT 375.920 -194.675 376.280 -194.040 ;
        RECT 376.970 -194.095 377.660 -194.040 ;
        RECT 375.920 -194.720 376.340 -194.675 ;
        RECT 362.300 -195.485 364.550 -195.395 ;
        RECT 360.090 -195.700 364.550 -195.485 ;
        RECT 360.090 -195.790 362.335 -195.700 ;
        RECT 364.245 -197.175 364.550 -195.700 ;
        RECT 367.915 -196.585 368.085 -195.115 ;
        RECT 368.375 -195.195 368.600 -194.845 ;
        RECT 370.335 -194.945 374.955 -194.745 ;
        RECT 370.575 -194.960 374.955 -194.945 ;
        RECT 367.880 -197.175 368.115 -196.585 ;
        RECT 368.405 -196.655 368.575 -195.195 ;
        RECT 368.895 -196.580 369.065 -195.115 ;
        RECT 370.105 -196.530 370.275 -195.115 ;
        RECT 370.575 -195.160 370.795 -194.960 ;
        RECT 375.945 -195.070 376.340 -194.720 ;
        RECT 368.860 -197.175 369.095 -196.580 ;
        RECT 370.070 -197.175 370.305 -196.530 ;
        RECT 370.595 -196.655 370.765 -195.160 ;
        RECT 377.385 -196.280 377.555 -194.825 ;
        RECT 377.375 -196.835 377.560 -196.280 ;
        RECT 377.875 -196.365 378.045 -193.140 ;
        RECT 379.020 -193.490 379.210 -193.140 ;
        RECT 380.220 -193.330 380.390 -192.935 ;
        RECT 381.595 -192.980 382.285 -192.935 ;
        RECT 378.970 -194.180 379.240 -193.490 ;
        RECT 379.735 -193.500 380.390 -193.330 ;
        RECT 380.720 -193.415 381.410 -193.145 ;
        RECT 382.645 -193.490 382.915 -192.800 ;
        RECT 383.105 -192.805 383.275 -192.585 ;
        RECT 383.105 -193.075 383.935 -192.805 ;
        RECT 379.735 -196.365 379.905 -193.500 ;
        RECT 383.105 -193.650 383.275 -193.075 ;
        RECT 383.535 -193.650 383.805 -193.565 ;
        RECT 380.225 -193.845 381.020 -193.670 ;
        RECT 383.105 -193.675 383.805 -193.650 ;
        RECT 382.965 -193.820 383.805 -193.675 ;
        RECT 380.225 -196.365 380.395 -193.845 ;
        RECT 380.850 -196.365 381.020 -193.845 ;
        RECT 381.340 -196.280 381.510 -193.825 ;
        RECT 381.990 -196.275 382.160 -193.825 ;
        RECT 374.690 -196.855 377.745 -196.835 ;
        RECT 381.335 -196.855 381.520 -196.280 ;
        RECT 381.975 -196.855 382.160 -196.275 ;
        RECT 382.480 -196.365 382.650 -193.825 ;
        RECT 382.965 -193.845 383.275 -193.820 ;
        RECT 382.970 -196.365 383.140 -193.845 ;
        RECT 383.535 -193.860 383.805 -193.820 ;
        RECT 384.110 -194.410 384.300 -191.945 ;
        RECT 407.500 -192.530 407.670 -190.810 ;
        RECT 408.480 -192.530 408.650 -190.810 ;
        RECT 410.545 -191.345 410.715 -190.805 ;
        RECT 411.525 -191.345 411.695 -190.805 ;
        RECT 409.955 -191.580 410.320 -191.515 ;
        RECT 409.455 -191.720 410.320 -191.580 ;
        RECT 409.345 -191.785 410.320 -191.720 ;
        RECT 409.345 -192.530 409.650 -191.785 ;
        RECT 409.955 -191.815 410.320 -191.785 ;
        RECT 412.505 -191.665 412.675 -190.805 ;
        RECT 407.500 -192.680 409.650 -192.530 ;
        RECT 407.500 -192.720 409.595 -192.680 ;
        RECT 410.545 -192.740 410.715 -191.960 ;
        RECT 411.035 -192.500 411.205 -191.960 ;
        RECT 411.525 -192.740 411.695 -191.960 ;
        RECT 412.015 -192.500 412.185 -191.960 ;
        RECT 412.505 -192.015 413.895 -191.665 ;
        RECT 405.720 -193.085 406.855 -193.075 ;
        RECT 408.910 -193.085 409.280 -192.955 ;
        RECT 405.720 -193.275 409.280 -193.085 ;
        RECT 409.845 -193.170 412.920 -192.740 ;
        RECT 384.110 -194.600 385.570 -194.410 ;
        RECT 383.620 -196.270 383.790 -194.825 ;
        RECT 384.110 -194.850 384.300 -194.600 ;
        RECT 383.610 -196.855 383.795 -196.270 ;
        RECT 384.110 -196.365 384.280 -194.850 ;
        RECT 374.690 -197.175 384.360 -196.855 ;
        RECT 364.245 -197.400 384.360 -197.175 ;
        RECT 364.245 -197.740 375.255 -197.400 ;
        RECT 376.995 -197.660 384.360 -197.400 ;
        RECT 309.625 -199.455 329.740 -199.190 ;
        RECT 287.100 -201.570 287.290 -199.680 ;
        RECT 293.135 -201.175 296.460 -201.035 ;
        RECT 293.135 -201.465 298.310 -201.175 ;
        RECT 286.985 -201.840 287.350 -201.570 ;
        RECT 293.135 -201.870 293.565 -201.465 ;
        RECT 294.435 -201.650 294.610 -201.465 ;
        RECT 296.060 -201.480 298.310 -201.465 ;
        RECT 288.875 -202.300 293.565 -201.870 ;
        RECT 288.115 -203.420 288.765 -203.290 ;
        RECT 285.590 -203.750 288.765 -203.420 ;
        RECT 289.575 -203.580 289.745 -202.300 ;
        RECT 290.065 -203.580 290.235 -202.540 ;
        RECT 290.555 -203.580 290.725 -202.300 ;
        RECT 291.045 -203.410 291.215 -202.540 ;
        RECT 293.950 -203.190 294.120 -201.650 ;
        RECT 294.440 -203.190 294.610 -201.650 ;
        RECT 294.930 -203.190 295.100 -201.650 ;
        RECT 295.420 -203.190 295.590 -201.650 ;
        RECT 295.910 -203.190 296.080 -201.650 ;
        RECT 293.790 -203.405 294.145 -203.400 ;
        RECT 295.850 -203.405 296.220 -203.375 ;
        RECT 293.790 -203.410 296.220 -203.405 ;
        RECT 291.045 -203.580 296.220 -203.410 ;
        RECT 298.005 -203.515 298.310 -201.480 ;
        RECT 291.050 -203.600 296.220 -203.580 ;
        RECT 291.050 -203.610 293.795 -203.600 ;
        RECT 288.985 -203.750 289.350 -203.720 ;
        RECT 295.850 -203.730 296.220 -203.600 ;
        RECT 285.590 -203.800 289.350 -203.750 ;
        RECT 288.115 -203.955 289.350 -203.800 ;
        RECT 293.525 -203.890 294.200 -203.850 ;
        RECT 293.425 -203.900 294.200 -203.890 ;
        RECT 288.115 -204.040 288.765 -203.955 ;
        RECT 288.985 -204.020 289.350 -203.955 ;
        RECT 288.250 -204.290 288.630 -204.040 ;
        RECT 292.390 -204.080 294.200 -203.900 ;
        RECT 296.785 -203.945 300.710 -203.515 ;
        RECT 293.425 -204.090 294.200 -204.080 ;
        RECT 293.525 -204.120 294.200 -204.090 ;
        RECT 294.440 -204.005 296.535 -203.965 ;
        RECT 294.440 -204.155 296.590 -204.005 ;
        RECT 289.575 -205.230 289.745 -204.190 ;
        RECT 290.555 -205.230 290.725 -204.190 ;
        RECT 291.535 -205.230 291.705 -204.190 ;
        RECT 294.440 -205.875 294.610 -204.155 ;
        RECT 295.420 -205.875 295.590 -204.155 ;
        RECT 296.285 -204.900 296.590 -204.155 ;
        RECT 297.485 -204.725 297.655 -203.945 ;
        RECT 297.975 -204.725 298.145 -204.185 ;
        RECT 298.465 -204.725 298.635 -203.945 ;
        RECT 298.955 -204.725 299.125 -204.185 ;
        RECT 296.895 -204.900 297.260 -204.870 ;
        RECT 296.285 -204.965 297.260 -204.900 ;
        RECT 296.395 -205.105 297.260 -204.965 ;
        RECT 296.895 -205.170 297.260 -205.105 ;
        RECT 299.445 -205.020 301.305 -204.670 ;
        RECT 297.485 -205.880 297.655 -205.340 ;
        RECT 298.465 -205.880 298.635 -205.340 ;
        RECT 299.445 -205.880 299.615 -205.020 ;
        RECT 297.715 -208.220 298.915 -208.050 ;
        RECT 289.445 -210.555 289.615 -208.835 ;
        RECT 290.425 -210.555 290.595 -208.835 ;
        RECT 292.490 -209.370 292.660 -208.830 ;
        RECT 293.470 -209.370 293.640 -208.830 ;
        RECT 291.900 -209.605 292.265 -209.540 ;
        RECT 291.400 -209.745 292.265 -209.605 ;
        RECT 291.290 -209.810 292.265 -209.745 ;
        RECT 291.290 -210.555 291.595 -209.810 ;
        RECT 291.900 -209.840 292.265 -209.810 ;
        RECT 294.450 -209.690 294.620 -208.830 ;
        RECT 289.445 -210.705 291.595 -210.555 ;
        RECT 289.445 -210.745 291.540 -210.705 ;
        RECT 292.490 -210.765 292.660 -209.985 ;
        RECT 292.980 -210.525 293.150 -209.985 ;
        RECT 293.470 -210.765 293.640 -209.985 ;
        RECT 293.960 -210.525 294.130 -209.985 ;
        RECT 294.450 -210.040 295.840 -209.690 ;
        RECT 287.665 -211.110 288.800 -211.100 ;
        RECT 290.855 -211.110 291.225 -210.980 ;
        RECT 283.955 -211.395 285.380 -211.180 ;
        RECT 287.665 -211.300 291.225 -211.110 ;
        RECT 291.790 -211.195 294.865 -210.765 ;
        RECT 288.795 -211.305 291.225 -211.300 ;
        RECT 288.795 -211.310 289.150 -211.305 ;
        RECT 290.855 -211.335 291.225 -211.305 ;
        RECT 282.560 -211.910 283.085 -211.550 ;
        RECT 285.165 -212.425 285.380 -211.395 ;
        RECT 272.725 -213.165 274.975 -213.075 ;
        RECT 270.515 -213.380 274.975 -213.165 ;
        RECT 270.515 -213.470 272.760 -213.380 ;
        RECT 274.670 -214.855 274.975 -213.380 ;
        RECT 278.340 -214.265 278.510 -212.795 ;
        RECT 278.800 -212.875 279.025 -212.525 ;
        RECT 280.760 -212.625 285.380 -212.425 ;
        RECT 281.000 -212.640 285.380 -212.625 ;
        RECT 278.305 -214.855 278.540 -214.265 ;
        RECT 278.830 -214.335 279.000 -212.875 ;
        RECT 279.320 -214.260 279.490 -212.795 ;
        RECT 280.530 -214.210 280.700 -212.795 ;
        RECT 281.000 -212.840 281.220 -212.640 ;
        RECT 279.285 -214.855 279.520 -214.260 ;
        RECT 280.495 -214.855 280.730 -214.210 ;
        RECT 281.020 -214.335 281.190 -212.840 ;
        RECT 288.955 -213.060 289.125 -211.520 ;
        RECT 289.445 -213.060 289.615 -211.520 ;
        RECT 289.935 -213.060 290.105 -211.520 ;
        RECT 290.425 -213.060 290.595 -211.520 ;
        RECT 290.915 -213.060 291.085 -211.520 ;
        RECT 289.440 -213.320 289.615 -213.060 ;
        RECT 293.010 -213.230 293.315 -211.195 ;
        RECT 295.460 -212.015 295.810 -210.040 ;
        RECT 296.680 -211.310 296.850 -208.390 ;
        RECT 297.715 -208.430 297.925 -208.220 ;
        RECT 296.660 -211.605 296.870 -211.310 ;
        RECT 297.735 -211.340 297.905 -208.430 ;
        RECT 298.225 -211.330 298.395 -208.390 ;
        RECT 298.705 -208.440 298.915 -208.220 ;
        RECT 297.720 -211.605 297.930 -211.340 ;
        RECT 296.660 -211.785 297.930 -211.605 ;
        RECT 298.205 -211.600 298.415 -211.330 ;
        RECT 298.715 -211.430 298.885 -208.440 ;
        RECT 299.775 -211.360 299.945 -208.390 ;
        RECT 298.205 -211.795 298.910 -211.600 ;
        RECT 298.695 -211.855 298.910 -211.795 ;
        RECT 297.485 -212.015 298.260 -211.965 ;
        RECT 295.460 -212.195 298.260 -212.015 ;
        RECT 295.460 -212.205 295.810 -212.195 ;
        RECT 297.485 -212.240 298.260 -212.195 ;
        RECT 298.695 -212.130 299.600 -211.855 ;
        RECT 298.695 -212.480 298.910 -212.130 ;
        RECT 296.135 -212.550 296.910 -212.505 ;
        RECT 295.950 -212.720 296.910 -212.550 ;
        RECT 296.135 -212.780 296.910 -212.720 ;
        RECT 297.140 -212.680 298.910 -212.480 ;
        RECT 299.770 -212.580 299.985 -211.360 ;
        RECT 300.955 -211.705 301.305 -205.020 ;
        RECT 300.900 -212.065 301.425 -211.705 ;
        RECT 303.190 -212.580 304.650 -211.735 ;
        RECT 291.065 -213.320 293.315 -213.230 ;
        RECT 288.855 -213.535 293.315 -213.320 ;
        RECT 288.855 -213.625 291.100 -213.535 ;
        RECT 274.670 -215.420 282.055 -214.855 ;
        RECT 293.010 -215.010 293.315 -213.535 ;
        RECT 296.680 -214.420 296.850 -212.950 ;
        RECT 297.140 -213.030 297.365 -212.680 ;
        RECT 299.100 -212.780 305.110 -212.580 ;
        RECT 299.340 -212.795 305.110 -212.780 ;
        RECT 296.645 -215.010 296.880 -214.420 ;
        RECT 297.170 -214.490 297.340 -213.030 ;
        RECT 297.660 -214.415 297.830 -212.950 ;
        RECT 298.870 -214.365 299.040 -212.950 ;
        RECT 299.340 -212.995 299.560 -212.795 ;
        RECT 297.625 -215.010 297.860 -214.415 ;
        RECT 298.835 -215.010 299.070 -214.365 ;
        RECT 299.360 -214.490 299.530 -212.995 ;
        RECT 303.190 -213.230 304.650 -212.795 ;
        RECT 293.010 -215.575 300.395 -215.010 ;
        RECT 265.775 -219.480 266.745 -218.645 ;
        RECT 46.135 -220.955 46.895 -220.685 ;
        RECT 46.135 -221.160 46.405 -220.955 ;
        RECT -95.030 -221.385 -94.340 -221.380 ;
        RECT -111.060 -221.610 -110.270 -221.445 ;
        RECT -36.555 -221.475 -35.740 -221.380 ;
        RECT -95.720 -221.610 -95.035 -221.585 ;
        RECT -111.060 -221.870 -95.035 -221.610 ;
        RECT -111.060 -222.025 -110.270 -221.870 ;
        RECT -95.720 -221.875 -95.035 -221.870 ;
        RECT 211.460 -223.555 212.790 -219.655 ;
        RECT 309.625 -222.305 310.710 -199.455 ;
        RECT 313.190 -199.570 329.740 -199.455 ;
        RECT 313.190 -200.480 313.570 -199.570 ;
        RECT 313.190 -200.860 313.900 -200.480 ;
        RECT 313.520 -202.805 313.900 -200.860 ;
        RECT 318.565 -200.690 321.890 -200.550 ;
        RECT 318.565 -200.980 323.740 -200.690 ;
        RECT 327.610 -200.975 328.070 -200.550 ;
        RECT 318.565 -201.385 318.995 -200.980 ;
        RECT 319.865 -201.165 320.040 -200.980 ;
        RECT 321.490 -200.995 323.740 -200.980 ;
        RECT 314.305 -201.815 318.995 -201.385 ;
        RECT 313.520 -203.265 314.195 -202.805 ;
        RECT 315.005 -203.095 315.175 -201.815 ;
        RECT 315.495 -203.095 315.665 -202.055 ;
        RECT 315.985 -203.095 316.155 -201.815 ;
        RECT 316.475 -202.925 316.645 -202.055 ;
        RECT 319.380 -202.705 319.550 -201.165 ;
        RECT 319.870 -202.705 320.040 -201.165 ;
        RECT 320.360 -202.705 320.530 -201.165 ;
        RECT 320.850 -202.705 321.020 -201.165 ;
        RECT 321.340 -202.705 321.510 -201.165 ;
        RECT 319.220 -202.920 319.575 -202.915 ;
        RECT 321.280 -202.920 321.650 -202.890 ;
        RECT 319.220 -202.925 321.650 -202.920 ;
        RECT 316.475 -203.095 321.650 -202.925 ;
        RECT 323.435 -203.030 323.740 -200.995 ;
        RECT 316.480 -203.115 321.650 -203.095 ;
        RECT 316.480 -203.125 319.225 -203.115 ;
        RECT 314.415 -203.265 314.780 -203.235 ;
        RECT 321.280 -203.245 321.650 -203.115 ;
        RECT 313.520 -203.350 314.780 -203.265 ;
        RECT 313.545 -203.470 314.780 -203.350 ;
        RECT 318.955 -203.405 319.630 -203.365 ;
        RECT 318.855 -203.415 319.630 -203.405 ;
        RECT 313.545 -203.555 314.195 -203.470 ;
        RECT 314.415 -203.535 314.780 -203.470 ;
        RECT 317.820 -203.595 319.630 -203.415 ;
        RECT 322.215 -203.460 326.140 -203.030 ;
        RECT 318.855 -203.605 319.630 -203.595 ;
        RECT 318.955 -203.635 319.630 -203.605 ;
        RECT 319.870 -203.520 321.965 -203.480 ;
        RECT 319.870 -203.670 322.020 -203.520 ;
        RECT 315.005 -204.745 315.175 -203.705 ;
        RECT 315.985 -204.745 316.155 -203.705 ;
        RECT 316.965 -204.745 317.135 -203.705 ;
        RECT 319.870 -205.390 320.040 -203.670 ;
        RECT 320.850 -205.390 321.020 -203.670 ;
        RECT 321.715 -204.415 322.020 -203.670 ;
        RECT 322.915 -204.240 323.085 -203.460 ;
        RECT 323.405 -204.240 323.575 -203.700 ;
        RECT 323.895 -204.240 324.065 -203.460 ;
        RECT 324.385 -204.240 324.555 -203.700 ;
        RECT 322.325 -204.415 322.690 -204.385 ;
        RECT 321.715 -204.480 322.690 -204.415 ;
        RECT 321.825 -204.620 322.690 -204.480 ;
        RECT 322.325 -204.685 322.690 -204.620 ;
        RECT 324.875 -204.535 326.735 -204.185 ;
        RECT 322.915 -205.395 323.085 -204.855 ;
        RECT 323.895 -205.395 324.065 -204.855 ;
        RECT 324.875 -205.395 325.045 -204.535 ;
        RECT 323.145 -207.735 324.345 -207.565 ;
        RECT 314.875 -210.070 315.045 -208.350 ;
        RECT 315.855 -210.070 316.025 -208.350 ;
        RECT 317.920 -208.885 318.090 -208.345 ;
        RECT 318.900 -208.885 319.070 -208.345 ;
        RECT 317.330 -209.120 317.695 -209.055 ;
        RECT 316.830 -209.260 317.695 -209.120 ;
        RECT 316.720 -209.325 317.695 -209.260 ;
        RECT 316.720 -210.070 317.025 -209.325 ;
        RECT 317.330 -209.355 317.695 -209.325 ;
        RECT 319.880 -209.205 320.050 -208.345 ;
        RECT 313.960 -210.135 314.635 -210.105 ;
        RECT 313.860 -210.145 314.635 -210.135 ;
        RECT 311.220 -210.325 314.635 -210.145 ;
        RECT 314.875 -210.220 317.025 -210.070 ;
        RECT 314.875 -210.260 316.970 -210.220 ;
        RECT 317.920 -210.280 318.090 -209.500 ;
        RECT 318.410 -210.040 318.580 -209.500 ;
        RECT 318.900 -210.280 319.070 -209.500 ;
        RECT 319.390 -210.040 319.560 -209.500 ;
        RECT 319.880 -209.555 321.270 -209.205 ;
        RECT 312.135 -215.460 312.815 -210.325 ;
        RECT 313.860 -210.335 314.635 -210.325 ;
        RECT 313.960 -210.375 314.635 -210.335 ;
        RECT 313.095 -210.625 314.230 -210.615 ;
        RECT 316.285 -210.625 316.655 -210.495 ;
        RECT 313.095 -210.815 316.655 -210.625 ;
        RECT 317.220 -210.710 320.295 -210.280 ;
        RECT 314.225 -210.820 316.655 -210.815 ;
        RECT 314.225 -210.825 314.580 -210.820 ;
        RECT 316.285 -210.850 316.655 -210.820 ;
        RECT 314.385 -212.575 314.555 -211.035 ;
        RECT 314.875 -212.575 315.045 -211.035 ;
        RECT 315.365 -212.575 315.535 -211.035 ;
        RECT 315.855 -212.575 316.025 -211.035 ;
        RECT 316.345 -212.575 316.515 -211.035 ;
        RECT 314.870 -212.835 315.045 -212.575 ;
        RECT 318.440 -212.745 318.745 -210.710 ;
        RECT 320.890 -211.530 321.240 -209.555 ;
        RECT 322.110 -210.825 322.280 -207.905 ;
        RECT 323.145 -207.945 323.355 -207.735 ;
        RECT 322.090 -211.120 322.300 -210.825 ;
        RECT 323.165 -210.855 323.335 -207.945 ;
        RECT 323.655 -210.845 323.825 -207.905 ;
        RECT 324.135 -207.955 324.345 -207.735 ;
        RECT 323.150 -211.120 323.360 -210.855 ;
        RECT 322.090 -211.300 323.360 -211.120 ;
        RECT 323.635 -211.115 323.845 -210.845 ;
        RECT 324.145 -210.945 324.315 -207.955 ;
        RECT 325.205 -210.875 325.375 -207.905 ;
        RECT 323.635 -211.310 324.340 -211.115 ;
        RECT 324.125 -211.370 324.340 -211.310 ;
        RECT 322.915 -211.530 323.690 -211.480 ;
        RECT 320.890 -211.710 323.690 -211.530 ;
        RECT 320.890 -211.720 321.240 -211.710 ;
        RECT 322.915 -211.755 323.690 -211.710 ;
        RECT 324.125 -211.645 325.030 -211.370 ;
        RECT 324.125 -211.995 324.340 -211.645 ;
        RECT 321.565 -212.065 322.340 -212.020 ;
        RECT 321.380 -212.235 322.340 -212.065 ;
        RECT 321.565 -212.295 322.340 -212.235 ;
        RECT 322.570 -212.195 324.340 -211.995 ;
        RECT 325.200 -212.095 325.415 -210.875 ;
        RECT 326.385 -211.220 326.735 -204.535 ;
        RECT 327.725 -210.850 327.940 -200.975 ;
        RECT 329.360 -203.090 329.740 -199.570 ;
        RECT 330.870 -199.350 339.805 -199.160 ;
        RECT 355.580 -199.105 359.335 -198.575 ;
        RECT 385.380 -199.075 385.570 -194.600 ;
        RECT 405.775 -198.180 406.155 -193.275 ;
        RECT 406.850 -193.280 409.280 -193.275 ;
        RECT 406.850 -193.285 407.205 -193.280 ;
        RECT 408.910 -193.310 409.280 -193.280 ;
        RECT 407.010 -195.035 407.180 -193.495 ;
        RECT 407.500 -195.035 407.670 -193.495 ;
        RECT 407.990 -195.035 408.160 -193.495 ;
        RECT 408.480 -195.035 408.650 -193.495 ;
        RECT 408.970 -195.035 409.140 -193.495 ;
        RECT 407.495 -195.295 407.670 -195.035 ;
        RECT 411.065 -195.205 411.370 -193.170 ;
        RECT 413.515 -193.990 413.865 -192.015 ;
        RECT 414.735 -193.285 414.905 -190.365 ;
        RECT 415.770 -190.405 415.980 -190.195 ;
        RECT 414.715 -193.580 414.925 -193.285 ;
        RECT 415.790 -193.315 415.960 -190.405 ;
        RECT 416.280 -193.305 416.450 -190.365 ;
        RECT 416.760 -190.415 416.970 -190.195 ;
        RECT 415.775 -193.580 415.985 -193.315 ;
        RECT 414.715 -193.760 415.985 -193.580 ;
        RECT 416.260 -193.575 416.470 -193.305 ;
        RECT 416.770 -193.405 416.940 -190.415 ;
        RECT 417.830 -193.335 418.000 -190.365 ;
        RECT 416.260 -193.770 416.965 -193.575 ;
        RECT 416.750 -193.830 416.965 -193.770 ;
        RECT 415.540 -193.990 416.315 -193.940 ;
        RECT 413.515 -194.170 416.315 -193.990 ;
        RECT 413.515 -194.180 413.865 -194.170 ;
        RECT 415.540 -194.215 416.315 -194.170 ;
        RECT 416.750 -194.105 417.655 -193.830 ;
        RECT 416.750 -194.455 416.965 -194.105 ;
        RECT 414.190 -194.525 414.965 -194.480 ;
        RECT 414.005 -194.695 414.965 -194.525 ;
        RECT 414.190 -194.755 414.965 -194.695 ;
        RECT 415.195 -194.655 416.965 -194.455 ;
        RECT 417.825 -194.555 418.040 -193.335 ;
        RECT 419.010 -193.680 419.360 -186.995 ;
        RECT 425.590 -189.475 427.195 -189.305 ;
        RECT 424.695 -192.155 424.865 -189.655 ;
        RECT 424.690 -192.385 424.865 -192.155 ;
        RECT 425.590 -192.385 425.790 -189.475 ;
        RECT 426.035 -189.675 426.210 -189.475 ;
        RECT 426.040 -192.195 426.210 -189.675 ;
        RECT 426.530 -192.160 426.700 -189.655 ;
        RECT 427.020 -189.670 427.195 -189.475 ;
        RECT 424.690 -192.585 425.790 -192.385 ;
        RECT 426.515 -192.760 426.705 -192.160 ;
        RECT 427.020 -192.195 427.190 -189.670 ;
        RECT 427.670 -192.575 427.840 -189.655 ;
        RECT 429.300 -192.225 429.470 -189.655 ;
        RECT 430.440 -191.105 430.610 -189.655 ;
        RECT 430.435 -191.570 430.620 -191.105 ;
        RECT 430.435 -191.755 431.120 -191.570 ;
        RECT 429.300 -192.395 430.095 -192.225 ;
        RECT 428.415 -192.575 429.105 -192.520 ;
        RECT 424.695 -192.950 426.705 -192.760 ;
        RECT 427.040 -192.745 429.105 -192.575 ;
        RECT 423.510 -193.005 424.200 -192.955 ;
        RECT 421.560 -193.175 424.200 -193.005 ;
        RECT 418.955 -194.040 419.480 -193.680 ;
        RECT 421.560 -194.555 421.775 -193.175 ;
        RECT 423.510 -193.225 424.200 -193.175 ;
        RECT 423.790 -193.680 424.480 -193.635 ;
        RECT 422.740 -193.850 424.480 -193.680 ;
        RECT 422.740 -194.485 423.100 -193.850 ;
        RECT 423.790 -193.905 424.480 -193.850 ;
        RECT 422.740 -194.530 423.160 -194.485 ;
        RECT 409.120 -195.295 411.370 -195.205 ;
        RECT 406.910 -195.510 411.370 -195.295 ;
        RECT 406.910 -195.600 409.155 -195.510 ;
        RECT 411.065 -196.985 411.370 -195.510 ;
        RECT 414.735 -196.395 414.905 -194.925 ;
        RECT 415.195 -195.005 415.420 -194.655 ;
        RECT 417.155 -194.755 421.775 -194.555 ;
        RECT 417.395 -194.770 421.775 -194.755 ;
        RECT 414.700 -196.985 414.935 -196.395 ;
        RECT 415.225 -196.465 415.395 -195.005 ;
        RECT 415.715 -196.390 415.885 -194.925 ;
        RECT 416.925 -196.340 417.095 -194.925 ;
        RECT 417.395 -194.970 417.615 -194.770 ;
        RECT 422.765 -194.880 423.160 -194.530 ;
        RECT 415.680 -196.985 415.915 -196.390 ;
        RECT 416.890 -196.985 417.125 -196.340 ;
        RECT 417.415 -196.465 417.585 -194.970 ;
        RECT 424.205 -196.090 424.375 -194.635 ;
        RECT 424.195 -196.645 424.380 -196.090 ;
        RECT 424.695 -196.175 424.865 -192.950 ;
        RECT 425.840 -193.300 426.030 -192.950 ;
        RECT 427.040 -193.140 427.210 -192.745 ;
        RECT 428.415 -192.790 429.105 -192.745 ;
        RECT 425.790 -193.990 426.060 -193.300 ;
        RECT 426.555 -193.310 427.210 -193.140 ;
        RECT 427.540 -193.225 428.230 -192.955 ;
        RECT 429.465 -193.300 429.735 -192.610 ;
        RECT 429.925 -192.615 430.095 -192.395 ;
        RECT 429.925 -192.885 430.755 -192.615 ;
        RECT 426.555 -196.175 426.725 -193.310 ;
        RECT 429.925 -193.460 430.095 -192.885 ;
        RECT 430.355 -193.460 430.625 -193.375 ;
        RECT 427.045 -193.655 427.840 -193.480 ;
        RECT 429.925 -193.485 430.625 -193.460 ;
        RECT 429.785 -193.630 430.625 -193.485 ;
        RECT 427.045 -196.175 427.215 -193.655 ;
        RECT 427.670 -196.175 427.840 -193.655 ;
        RECT 428.160 -196.090 428.330 -193.635 ;
        RECT 428.810 -196.085 428.980 -193.635 ;
        RECT 421.510 -196.665 424.565 -196.645 ;
        RECT 428.155 -196.665 428.340 -196.090 ;
        RECT 428.795 -196.665 428.980 -196.085 ;
        RECT 429.300 -196.175 429.470 -193.635 ;
        RECT 429.785 -193.655 430.095 -193.630 ;
        RECT 429.790 -196.175 429.960 -193.655 ;
        RECT 430.355 -193.670 430.625 -193.630 ;
        RECT 430.930 -194.220 431.120 -191.755 ;
        RECT 430.930 -194.410 432.390 -194.220 ;
        RECT 430.440 -196.080 430.610 -194.635 ;
        RECT 430.930 -194.660 431.120 -194.410 ;
        RECT 430.430 -196.665 430.615 -196.080 ;
        RECT 430.930 -196.175 431.100 -194.660 ;
        RECT 421.510 -196.985 431.180 -196.665 ;
        RECT 411.065 -197.210 431.180 -196.985 ;
        RECT 411.065 -197.550 422.075 -197.210 ;
        RECT 423.815 -197.470 431.180 -197.210 ;
        RECT 330.870 -201.240 331.060 -199.350 ;
        RECT 355.580 -199.425 375.505 -199.105 ;
        RECT 336.905 -200.845 340.230 -200.705 ;
        RECT 336.905 -201.135 342.080 -200.845 ;
        RECT 330.755 -201.510 331.120 -201.240 ;
        RECT 336.905 -201.540 337.335 -201.135 ;
        RECT 338.205 -201.320 338.380 -201.135 ;
        RECT 339.830 -201.150 342.080 -201.135 ;
        RECT 332.645 -201.970 337.335 -201.540 ;
        RECT 331.885 -203.090 332.535 -202.960 ;
        RECT 329.360 -203.420 332.535 -203.090 ;
        RECT 333.345 -203.250 333.515 -201.970 ;
        RECT 333.835 -203.250 334.005 -202.210 ;
        RECT 334.325 -203.250 334.495 -201.970 ;
        RECT 334.815 -203.080 334.985 -202.210 ;
        RECT 337.720 -202.860 337.890 -201.320 ;
        RECT 338.210 -202.860 338.380 -201.320 ;
        RECT 338.700 -202.860 338.870 -201.320 ;
        RECT 339.190 -202.860 339.360 -201.320 ;
        RECT 339.680 -202.860 339.850 -201.320 ;
        RECT 337.560 -203.075 337.915 -203.070 ;
        RECT 339.620 -203.075 339.990 -203.045 ;
        RECT 337.560 -203.080 339.990 -203.075 ;
        RECT 334.815 -203.250 339.990 -203.080 ;
        RECT 341.775 -203.185 342.080 -201.150 ;
        RECT 334.820 -203.270 339.990 -203.250 ;
        RECT 334.820 -203.280 337.565 -203.270 ;
        RECT 332.755 -203.420 333.120 -203.390 ;
        RECT 339.620 -203.400 339.990 -203.270 ;
        RECT 329.360 -203.470 333.120 -203.420 ;
        RECT 331.885 -203.625 333.120 -203.470 ;
        RECT 337.295 -203.560 337.970 -203.520 ;
        RECT 337.195 -203.570 337.970 -203.560 ;
        RECT 331.885 -203.710 332.535 -203.625 ;
        RECT 332.755 -203.690 333.120 -203.625 ;
        RECT 332.020 -203.960 332.400 -203.710 ;
        RECT 336.160 -203.750 337.970 -203.570 ;
        RECT 340.555 -203.615 344.480 -203.185 ;
        RECT 337.195 -203.760 337.970 -203.750 ;
        RECT 337.295 -203.790 337.970 -203.760 ;
        RECT 338.210 -203.675 340.305 -203.635 ;
        RECT 338.210 -203.825 340.360 -203.675 ;
        RECT 333.345 -204.900 333.515 -203.860 ;
        RECT 334.325 -204.900 334.495 -203.860 ;
        RECT 335.305 -204.900 335.475 -203.860 ;
        RECT 338.210 -205.545 338.380 -203.825 ;
        RECT 339.190 -205.545 339.360 -203.825 ;
        RECT 340.055 -204.570 340.360 -203.825 ;
        RECT 341.255 -204.395 341.425 -203.615 ;
        RECT 341.745 -204.395 341.915 -203.855 ;
        RECT 342.235 -204.395 342.405 -203.615 ;
        RECT 342.725 -204.395 342.895 -203.855 ;
        RECT 340.665 -204.570 341.030 -204.540 ;
        RECT 340.055 -204.635 341.030 -204.570 ;
        RECT 340.165 -204.775 341.030 -204.635 ;
        RECT 340.665 -204.840 341.030 -204.775 ;
        RECT 343.215 -204.690 345.075 -204.340 ;
        RECT 341.255 -205.550 341.425 -205.010 ;
        RECT 342.235 -205.550 342.405 -205.010 ;
        RECT 343.215 -205.550 343.385 -204.690 ;
        RECT 341.485 -207.890 342.685 -207.720 ;
        RECT 333.215 -210.225 333.385 -208.505 ;
        RECT 334.195 -210.225 334.365 -208.505 ;
        RECT 336.260 -209.040 336.430 -208.500 ;
        RECT 337.240 -209.040 337.410 -208.500 ;
        RECT 335.670 -209.275 336.035 -209.210 ;
        RECT 335.170 -209.415 336.035 -209.275 ;
        RECT 335.060 -209.480 336.035 -209.415 ;
        RECT 335.060 -210.225 335.365 -209.480 ;
        RECT 335.670 -209.510 336.035 -209.480 ;
        RECT 338.220 -209.360 338.390 -208.500 ;
        RECT 332.300 -210.290 332.975 -210.260 ;
        RECT 332.200 -210.300 332.975 -210.290 ;
        RECT 330.130 -210.480 332.975 -210.300 ;
        RECT 333.215 -210.375 335.365 -210.225 ;
        RECT 333.215 -210.415 335.310 -210.375 ;
        RECT 336.260 -210.435 336.430 -209.655 ;
        RECT 336.750 -210.195 336.920 -209.655 ;
        RECT 337.240 -210.435 337.410 -209.655 ;
        RECT 337.730 -210.195 337.900 -209.655 ;
        RECT 338.220 -209.710 339.610 -209.360 ;
        RECT 327.725 -211.065 329.150 -210.850 ;
        RECT 326.330 -211.580 326.855 -211.220 ;
        RECT 328.935 -212.095 329.150 -211.065 ;
        RECT 316.495 -212.835 318.745 -212.745 ;
        RECT 314.285 -213.050 318.745 -212.835 ;
        RECT 314.285 -213.140 316.530 -213.050 ;
        RECT 318.440 -214.525 318.745 -213.050 ;
        RECT 322.110 -213.935 322.280 -212.465 ;
        RECT 322.570 -212.545 322.795 -212.195 ;
        RECT 324.530 -212.295 329.150 -212.095 ;
        RECT 324.770 -212.310 329.150 -212.295 ;
        RECT 322.075 -214.525 322.310 -213.935 ;
        RECT 322.600 -214.005 322.770 -212.545 ;
        RECT 323.090 -213.930 323.260 -212.465 ;
        RECT 324.300 -213.880 324.470 -212.465 ;
        RECT 324.770 -212.510 324.990 -212.310 ;
        RECT 323.055 -214.525 323.290 -213.930 ;
        RECT 324.265 -214.525 324.500 -213.880 ;
        RECT 324.790 -214.005 324.960 -212.510 ;
        RECT 318.440 -215.090 325.825 -214.525 ;
        RECT 330.130 -215.460 330.810 -210.480 ;
        RECT 332.200 -210.490 332.975 -210.480 ;
        RECT 332.300 -210.530 332.975 -210.490 ;
        RECT 331.435 -210.780 332.570 -210.770 ;
        RECT 334.625 -210.780 334.995 -210.650 ;
        RECT 331.435 -210.970 334.995 -210.780 ;
        RECT 335.560 -210.865 338.635 -210.435 ;
        RECT 332.565 -210.975 334.995 -210.970 ;
        RECT 332.565 -210.980 332.920 -210.975 ;
        RECT 334.625 -211.005 334.995 -210.975 ;
        RECT 332.725 -212.730 332.895 -211.190 ;
        RECT 333.215 -212.730 333.385 -211.190 ;
        RECT 333.705 -212.730 333.875 -211.190 ;
        RECT 334.195 -212.730 334.365 -211.190 ;
        RECT 334.685 -212.730 334.855 -211.190 ;
        RECT 333.210 -212.990 333.385 -212.730 ;
        RECT 336.780 -212.900 337.085 -210.865 ;
        RECT 339.230 -211.685 339.580 -209.710 ;
        RECT 340.450 -210.980 340.620 -208.060 ;
        RECT 341.485 -208.100 341.695 -207.890 ;
        RECT 340.430 -211.275 340.640 -210.980 ;
        RECT 341.505 -211.010 341.675 -208.100 ;
        RECT 341.995 -211.000 342.165 -208.060 ;
        RECT 342.475 -208.110 342.685 -207.890 ;
        RECT 341.490 -211.275 341.700 -211.010 ;
        RECT 340.430 -211.455 341.700 -211.275 ;
        RECT 341.975 -211.270 342.185 -211.000 ;
        RECT 342.485 -211.100 342.655 -208.110 ;
        RECT 343.545 -211.030 343.715 -208.060 ;
        RECT 341.975 -211.465 342.680 -211.270 ;
        RECT 342.465 -211.525 342.680 -211.465 ;
        RECT 341.255 -211.685 342.030 -211.635 ;
        RECT 339.230 -211.865 342.030 -211.685 ;
        RECT 339.230 -211.875 339.580 -211.865 ;
        RECT 341.255 -211.910 342.030 -211.865 ;
        RECT 342.465 -211.800 343.370 -211.525 ;
        RECT 342.465 -212.150 342.680 -211.800 ;
        RECT 339.905 -212.220 340.680 -212.175 ;
        RECT 339.720 -212.390 340.680 -212.220 ;
        RECT 339.905 -212.450 340.680 -212.390 ;
        RECT 340.910 -212.350 342.680 -212.150 ;
        RECT 343.540 -212.250 343.755 -211.030 ;
        RECT 344.725 -211.375 345.075 -204.690 ;
        RECT 344.670 -211.735 345.195 -211.375 ;
        RECT 347.015 -212.250 348.320 -211.445 ;
        RECT 334.835 -212.990 337.085 -212.900 ;
        RECT 332.625 -213.205 337.085 -212.990 ;
        RECT 332.625 -213.295 334.870 -213.205 ;
        RECT 336.780 -214.680 337.085 -213.205 ;
        RECT 340.450 -214.090 340.620 -212.620 ;
        RECT 340.910 -212.700 341.135 -212.350 ;
        RECT 342.870 -212.450 348.880 -212.250 ;
        RECT 343.110 -212.465 348.880 -212.450 ;
        RECT 340.415 -214.680 340.650 -214.090 ;
        RECT 340.940 -214.160 341.110 -212.700 ;
        RECT 341.430 -214.085 341.600 -212.620 ;
        RECT 342.640 -214.035 342.810 -212.620 ;
        RECT 343.110 -212.665 343.330 -212.465 ;
        RECT 341.395 -214.680 341.630 -214.085 ;
        RECT 342.605 -214.680 342.840 -214.035 ;
        RECT 343.130 -214.160 343.300 -212.665 ;
        RECT 347.015 -212.965 348.320 -212.465 ;
        RECT 336.780 -215.245 344.165 -214.680 ;
        RECT 312.135 -216.140 330.810 -215.460 ;
        RECT 211.545 -223.600 212.745 -223.555 ;
        RECT 309.340 -223.720 311.060 -222.305 ;
        RECT 44.935 -227.385 45.615 -227.375 ;
        RECT 312.135 -227.385 312.815 -216.140 ;
        RECT 355.580 -218.605 356.430 -199.425 ;
        RECT 358.955 -199.485 375.505 -199.425 ;
        RECT 358.955 -200.395 359.335 -199.485 ;
        RECT 358.955 -200.775 359.665 -200.395 ;
        RECT 359.285 -202.720 359.665 -200.775 ;
        RECT 364.330 -200.605 367.655 -200.465 ;
        RECT 364.330 -200.895 369.505 -200.605 ;
        RECT 373.375 -200.890 373.835 -200.465 ;
        RECT 364.330 -201.300 364.760 -200.895 ;
        RECT 365.630 -201.080 365.805 -200.895 ;
        RECT 367.255 -200.910 369.505 -200.895 ;
        RECT 360.070 -201.730 364.760 -201.300 ;
        RECT 359.285 -203.180 359.960 -202.720 ;
        RECT 360.770 -203.010 360.940 -201.730 ;
        RECT 361.260 -203.010 361.430 -201.970 ;
        RECT 361.750 -203.010 361.920 -201.730 ;
        RECT 362.240 -202.840 362.410 -201.970 ;
        RECT 365.145 -202.620 365.315 -201.080 ;
        RECT 365.635 -202.620 365.805 -201.080 ;
        RECT 366.125 -202.620 366.295 -201.080 ;
        RECT 366.615 -202.620 366.785 -201.080 ;
        RECT 367.105 -202.620 367.275 -201.080 ;
        RECT 364.985 -202.835 365.340 -202.830 ;
        RECT 367.045 -202.835 367.415 -202.805 ;
        RECT 364.985 -202.840 367.415 -202.835 ;
        RECT 362.240 -203.010 367.415 -202.840 ;
        RECT 369.200 -202.945 369.505 -200.910 ;
        RECT 362.245 -203.030 367.415 -203.010 ;
        RECT 362.245 -203.040 364.990 -203.030 ;
        RECT 360.180 -203.180 360.545 -203.150 ;
        RECT 367.045 -203.160 367.415 -203.030 ;
        RECT 359.285 -203.265 360.545 -203.180 ;
        RECT 359.310 -203.385 360.545 -203.265 ;
        RECT 364.720 -203.320 365.395 -203.280 ;
        RECT 364.620 -203.330 365.395 -203.320 ;
        RECT 359.310 -203.470 359.960 -203.385 ;
        RECT 360.180 -203.450 360.545 -203.385 ;
        RECT 363.585 -203.510 365.395 -203.330 ;
        RECT 367.980 -203.375 371.905 -202.945 ;
        RECT 364.620 -203.520 365.395 -203.510 ;
        RECT 364.720 -203.550 365.395 -203.520 ;
        RECT 365.635 -203.435 367.730 -203.395 ;
        RECT 365.635 -203.585 367.785 -203.435 ;
        RECT 360.770 -204.660 360.940 -203.620 ;
        RECT 361.750 -204.660 361.920 -203.620 ;
        RECT 362.730 -204.660 362.900 -203.620 ;
        RECT 365.635 -205.305 365.805 -203.585 ;
        RECT 366.615 -205.305 366.785 -203.585 ;
        RECT 367.480 -204.330 367.785 -203.585 ;
        RECT 368.680 -204.155 368.850 -203.375 ;
        RECT 369.170 -204.155 369.340 -203.615 ;
        RECT 369.660 -204.155 369.830 -203.375 ;
        RECT 370.150 -204.155 370.320 -203.615 ;
        RECT 368.090 -204.330 368.455 -204.300 ;
        RECT 367.480 -204.395 368.455 -204.330 ;
        RECT 367.590 -204.535 368.455 -204.395 ;
        RECT 368.090 -204.600 368.455 -204.535 ;
        RECT 370.640 -204.450 372.500 -204.100 ;
        RECT 368.680 -205.310 368.850 -204.770 ;
        RECT 369.660 -205.310 369.830 -204.770 ;
        RECT 370.640 -205.310 370.810 -204.450 ;
        RECT 368.910 -207.650 370.110 -207.480 ;
        RECT 360.640 -209.985 360.810 -208.265 ;
        RECT 361.620 -209.985 361.790 -208.265 ;
        RECT 363.685 -208.800 363.855 -208.260 ;
        RECT 364.665 -208.800 364.835 -208.260 ;
        RECT 363.095 -209.035 363.460 -208.970 ;
        RECT 362.595 -209.175 363.460 -209.035 ;
        RECT 362.485 -209.240 363.460 -209.175 ;
        RECT 362.485 -209.985 362.790 -209.240 ;
        RECT 363.095 -209.270 363.460 -209.240 ;
        RECT 365.645 -209.120 365.815 -208.260 ;
        RECT 359.725 -210.050 360.400 -210.020 ;
        RECT 359.625 -210.060 360.400 -210.050 ;
        RECT 356.985 -210.240 360.400 -210.060 ;
        RECT 360.640 -210.135 362.790 -209.985 ;
        RECT 360.640 -210.175 362.735 -210.135 ;
        RECT 363.685 -210.195 363.855 -209.415 ;
        RECT 364.175 -209.955 364.345 -209.415 ;
        RECT 364.665 -210.195 364.835 -209.415 ;
        RECT 365.155 -209.955 365.325 -209.415 ;
        RECT 365.645 -209.470 367.035 -209.120 ;
        RECT 357.900 -215.375 358.580 -210.240 ;
        RECT 359.625 -210.250 360.400 -210.240 ;
        RECT 359.725 -210.290 360.400 -210.250 ;
        RECT 358.860 -210.540 359.995 -210.530 ;
        RECT 362.050 -210.540 362.420 -210.410 ;
        RECT 358.860 -210.730 362.420 -210.540 ;
        RECT 362.985 -210.625 366.060 -210.195 ;
        RECT 359.990 -210.735 362.420 -210.730 ;
        RECT 359.990 -210.740 360.345 -210.735 ;
        RECT 362.050 -210.765 362.420 -210.735 ;
        RECT 360.150 -212.490 360.320 -210.950 ;
        RECT 360.640 -212.490 360.810 -210.950 ;
        RECT 361.130 -212.490 361.300 -210.950 ;
        RECT 361.620 -212.490 361.790 -210.950 ;
        RECT 362.110 -212.490 362.280 -210.950 ;
        RECT 360.635 -212.750 360.810 -212.490 ;
        RECT 364.205 -212.660 364.510 -210.625 ;
        RECT 366.655 -211.445 367.005 -209.470 ;
        RECT 367.875 -210.740 368.045 -207.820 ;
        RECT 368.910 -207.860 369.120 -207.650 ;
        RECT 367.855 -211.035 368.065 -210.740 ;
        RECT 368.930 -210.770 369.100 -207.860 ;
        RECT 369.420 -210.760 369.590 -207.820 ;
        RECT 369.900 -207.870 370.110 -207.650 ;
        RECT 368.915 -211.035 369.125 -210.770 ;
        RECT 367.855 -211.215 369.125 -211.035 ;
        RECT 369.400 -211.030 369.610 -210.760 ;
        RECT 369.910 -210.860 370.080 -207.870 ;
        RECT 370.970 -210.790 371.140 -207.820 ;
        RECT 369.400 -211.225 370.105 -211.030 ;
        RECT 369.890 -211.285 370.105 -211.225 ;
        RECT 368.680 -211.445 369.455 -211.395 ;
        RECT 366.655 -211.625 369.455 -211.445 ;
        RECT 366.655 -211.635 367.005 -211.625 ;
        RECT 368.680 -211.670 369.455 -211.625 ;
        RECT 369.890 -211.560 370.795 -211.285 ;
        RECT 369.890 -211.910 370.105 -211.560 ;
        RECT 367.330 -211.980 368.105 -211.935 ;
        RECT 367.145 -212.150 368.105 -211.980 ;
        RECT 367.330 -212.210 368.105 -212.150 ;
        RECT 368.335 -212.110 370.105 -211.910 ;
        RECT 370.965 -212.010 371.180 -210.790 ;
        RECT 372.150 -211.135 372.500 -204.450 ;
        RECT 373.490 -210.765 373.705 -200.890 ;
        RECT 375.125 -203.005 375.505 -199.485 ;
        RECT 376.635 -199.265 385.570 -199.075 ;
        RECT 401.960 -198.915 406.365 -198.180 ;
        RECT 432.200 -198.885 432.390 -194.410 ;
        RECT 376.635 -201.155 376.825 -199.265 ;
        RECT 401.960 -199.295 422.325 -198.915 ;
        RECT 401.960 -199.310 406.365 -199.295 ;
        RECT 382.670 -200.760 385.995 -200.620 ;
        RECT 382.670 -201.050 387.845 -200.760 ;
        RECT 376.520 -201.425 376.885 -201.155 ;
        RECT 382.670 -201.455 383.100 -201.050 ;
        RECT 383.970 -201.235 384.145 -201.050 ;
        RECT 385.595 -201.065 387.845 -201.050 ;
        RECT 378.410 -201.885 383.100 -201.455 ;
        RECT 377.650 -203.005 378.300 -202.875 ;
        RECT 375.125 -203.335 378.300 -203.005 ;
        RECT 379.110 -203.165 379.280 -201.885 ;
        RECT 379.600 -203.165 379.770 -202.125 ;
        RECT 380.090 -203.165 380.260 -201.885 ;
        RECT 380.580 -202.995 380.750 -202.125 ;
        RECT 383.485 -202.775 383.655 -201.235 ;
        RECT 383.975 -202.775 384.145 -201.235 ;
        RECT 384.465 -202.775 384.635 -201.235 ;
        RECT 384.955 -202.775 385.125 -201.235 ;
        RECT 385.445 -202.775 385.615 -201.235 ;
        RECT 383.325 -202.990 383.680 -202.985 ;
        RECT 385.385 -202.990 385.755 -202.960 ;
        RECT 383.325 -202.995 385.755 -202.990 ;
        RECT 380.580 -203.165 385.755 -202.995 ;
        RECT 387.540 -203.100 387.845 -201.065 ;
        RECT 380.585 -203.185 385.755 -203.165 ;
        RECT 380.585 -203.195 383.330 -203.185 ;
        RECT 378.520 -203.335 378.885 -203.305 ;
        RECT 385.385 -203.315 385.755 -203.185 ;
        RECT 375.125 -203.385 378.885 -203.335 ;
        RECT 377.650 -203.540 378.885 -203.385 ;
        RECT 383.060 -203.475 383.735 -203.435 ;
        RECT 382.960 -203.485 383.735 -203.475 ;
        RECT 377.650 -203.625 378.300 -203.540 ;
        RECT 378.520 -203.605 378.885 -203.540 ;
        RECT 377.785 -203.875 378.165 -203.625 ;
        RECT 381.925 -203.665 383.735 -203.485 ;
        RECT 386.320 -203.530 390.245 -203.100 ;
        RECT 382.960 -203.675 383.735 -203.665 ;
        RECT 383.060 -203.705 383.735 -203.675 ;
        RECT 383.975 -203.590 386.070 -203.550 ;
        RECT 383.975 -203.740 386.125 -203.590 ;
        RECT 379.110 -204.815 379.280 -203.775 ;
        RECT 380.090 -204.815 380.260 -203.775 ;
        RECT 381.070 -204.815 381.240 -203.775 ;
        RECT 383.975 -205.460 384.145 -203.740 ;
        RECT 384.955 -205.460 385.125 -203.740 ;
        RECT 385.820 -204.485 386.125 -203.740 ;
        RECT 387.020 -204.310 387.190 -203.530 ;
        RECT 387.510 -204.310 387.680 -203.770 ;
        RECT 388.000 -204.310 388.170 -203.530 ;
        RECT 388.490 -204.310 388.660 -203.770 ;
        RECT 386.430 -204.485 386.795 -204.455 ;
        RECT 385.820 -204.550 386.795 -204.485 ;
        RECT 385.930 -204.690 386.795 -204.550 ;
        RECT 386.430 -204.755 386.795 -204.690 ;
        RECT 388.980 -204.605 390.840 -204.255 ;
        RECT 387.020 -205.465 387.190 -204.925 ;
        RECT 388.000 -205.465 388.170 -204.925 ;
        RECT 388.980 -205.465 389.150 -204.605 ;
        RECT 387.250 -207.805 388.450 -207.635 ;
        RECT 378.980 -210.140 379.150 -208.420 ;
        RECT 379.960 -210.140 380.130 -208.420 ;
        RECT 382.025 -208.955 382.195 -208.415 ;
        RECT 383.005 -208.955 383.175 -208.415 ;
        RECT 381.435 -209.190 381.800 -209.125 ;
        RECT 380.935 -209.330 381.800 -209.190 ;
        RECT 380.825 -209.395 381.800 -209.330 ;
        RECT 380.825 -210.140 381.130 -209.395 ;
        RECT 381.435 -209.425 381.800 -209.395 ;
        RECT 383.985 -209.275 384.155 -208.415 ;
        RECT 378.065 -210.205 378.740 -210.175 ;
        RECT 377.965 -210.215 378.740 -210.205 ;
        RECT 375.895 -210.395 378.740 -210.215 ;
        RECT 378.980 -210.290 381.130 -210.140 ;
        RECT 378.980 -210.330 381.075 -210.290 ;
        RECT 382.025 -210.350 382.195 -209.570 ;
        RECT 382.515 -210.110 382.685 -209.570 ;
        RECT 383.005 -210.350 383.175 -209.570 ;
        RECT 383.495 -210.110 383.665 -209.570 ;
        RECT 383.985 -209.625 385.375 -209.275 ;
        RECT 373.490 -210.980 374.915 -210.765 ;
        RECT 372.095 -211.495 372.620 -211.135 ;
        RECT 374.700 -212.010 374.915 -210.980 ;
        RECT 362.260 -212.750 364.510 -212.660 ;
        RECT 360.050 -212.965 364.510 -212.750 ;
        RECT 360.050 -213.055 362.295 -212.965 ;
        RECT 364.205 -214.440 364.510 -212.965 ;
        RECT 367.875 -213.850 368.045 -212.380 ;
        RECT 368.335 -212.460 368.560 -212.110 ;
        RECT 370.295 -212.210 374.915 -212.010 ;
        RECT 370.535 -212.225 374.915 -212.210 ;
        RECT 367.840 -214.440 368.075 -213.850 ;
        RECT 368.365 -213.920 368.535 -212.460 ;
        RECT 368.855 -213.845 369.025 -212.380 ;
        RECT 370.065 -213.795 370.235 -212.380 ;
        RECT 370.535 -212.425 370.755 -212.225 ;
        RECT 368.820 -214.440 369.055 -213.845 ;
        RECT 370.030 -214.440 370.265 -213.795 ;
        RECT 370.555 -213.920 370.725 -212.425 ;
        RECT 364.205 -215.005 371.590 -214.440 ;
        RECT 375.895 -215.375 376.575 -210.395 ;
        RECT 377.965 -210.405 378.740 -210.395 ;
        RECT 378.065 -210.445 378.740 -210.405 ;
        RECT 377.200 -210.695 378.335 -210.685 ;
        RECT 380.390 -210.695 380.760 -210.565 ;
        RECT 377.200 -210.885 380.760 -210.695 ;
        RECT 381.325 -210.780 384.400 -210.350 ;
        RECT 378.330 -210.890 380.760 -210.885 ;
        RECT 378.330 -210.895 378.685 -210.890 ;
        RECT 380.390 -210.920 380.760 -210.890 ;
        RECT 378.490 -212.645 378.660 -211.105 ;
        RECT 378.980 -212.645 379.150 -211.105 ;
        RECT 379.470 -212.645 379.640 -211.105 ;
        RECT 379.960 -212.645 380.130 -211.105 ;
        RECT 380.450 -212.645 380.620 -211.105 ;
        RECT 378.975 -212.905 379.150 -212.645 ;
        RECT 382.545 -212.815 382.850 -210.780 ;
        RECT 384.995 -211.600 385.345 -209.625 ;
        RECT 386.215 -210.895 386.385 -207.975 ;
        RECT 387.250 -208.015 387.460 -207.805 ;
        RECT 386.195 -211.190 386.405 -210.895 ;
        RECT 387.270 -210.925 387.440 -208.015 ;
        RECT 387.760 -210.915 387.930 -207.975 ;
        RECT 388.240 -208.025 388.450 -207.805 ;
        RECT 387.255 -211.190 387.465 -210.925 ;
        RECT 386.195 -211.370 387.465 -211.190 ;
        RECT 387.740 -211.185 387.950 -210.915 ;
        RECT 388.250 -211.015 388.420 -208.025 ;
        RECT 389.310 -210.945 389.480 -207.975 ;
        RECT 387.740 -211.380 388.445 -211.185 ;
        RECT 388.230 -211.440 388.445 -211.380 ;
        RECT 387.020 -211.600 387.795 -211.550 ;
        RECT 384.995 -211.780 387.795 -211.600 ;
        RECT 384.995 -211.790 385.345 -211.780 ;
        RECT 387.020 -211.825 387.795 -211.780 ;
        RECT 388.230 -211.715 389.135 -211.440 ;
        RECT 388.230 -212.065 388.445 -211.715 ;
        RECT 385.670 -212.135 386.445 -212.090 ;
        RECT 385.485 -212.305 386.445 -212.135 ;
        RECT 385.670 -212.365 386.445 -212.305 ;
        RECT 386.675 -212.265 388.445 -212.065 ;
        RECT 389.305 -212.165 389.520 -210.945 ;
        RECT 390.490 -211.290 390.840 -204.605 ;
        RECT 390.435 -211.650 390.960 -211.290 ;
        RECT 393.445 -212.165 393.955 -211.975 ;
        RECT 380.600 -212.905 382.850 -212.815 ;
        RECT 378.390 -213.120 382.850 -212.905 ;
        RECT 378.390 -213.210 380.635 -213.120 ;
        RECT 382.545 -214.595 382.850 -213.120 ;
        RECT 386.215 -214.005 386.385 -212.535 ;
        RECT 386.675 -212.615 386.900 -212.265 ;
        RECT 388.635 -212.365 394.645 -212.165 ;
        RECT 388.875 -212.380 394.645 -212.365 ;
        RECT 386.180 -214.595 386.415 -214.005 ;
        RECT 386.705 -214.075 386.875 -212.615 ;
        RECT 387.195 -214.000 387.365 -212.535 ;
        RECT 388.405 -213.950 388.575 -212.535 ;
        RECT 388.875 -212.580 389.095 -212.380 ;
        RECT 393.445 -212.530 393.955 -212.380 ;
        RECT 387.160 -214.595 387.395 -214.000 ;
        RECT 388.370 -214.595 388.605 -213.950 ;
        RECT 388.895 -214.075 389.065 -212.580 ;
        RECT 382.545 -215.160 389.930 -214.595 ;
        RECT 357.900 -216.055 376.575 -215.375 ;
        RECT 355.385 -219.505 356.615 -218.605 ;
        RECT -121.070 -228.065 312.815 -227.385 ;
        RECT -121.070 -228.090 -111.215 -228.065 ;
        RECT -121.070 -228.880 -120.390 -228.090 ;
        RECT 357.900 -228.880 358.580 -216.055 ;
        RECT 401.960 -222.320 403.090 -199.310 ;
        RECT 405.775 -200.205 406.155 -199.310 ;
        RECT 405.775 -200.585 406.485 -200.205 ;
        RECT 406.105 -202.530 406.485 -200.585 ;
        RECT 411.150 -200.415 414.475 -200.275 ;
        RECT 411.150 -200.705 416.325 -200.415 ;
        RECT 420.195 -200.700 420.655 -200.275 ;
        RECT 411.150 -201.110 411.580 -200.705 ;
        RECT 412.450 -200.890 412.625 -200.705 ;
        RECT 414.075 -200.720 416.325 -200.705 ;
        RECT 406.890 -201.540 411.580 -201.110 ;
        RECT 406.105 -202.990 406.780 -202.530 ;
        RECT 407.590 -202.820 407.760 -201.540 ;
        RECT 408.080 -202.820 408.250 -201.780 ;
        RECT 408.570 -202.820 408.740 -201.540 ;
        RECT 409.060 -202.650 409.230 -201.780 ;
        RECT 411.965 -202.430 412.135 -200.890 ;
        RECT 412.455 -202.430 412.625 -200.890 ;
        RECT 412.945 -202.430 413.115 -200.890 ;
        RECT 413.435 -202.430 413.605 -200.890 ;
        RECT 413.925 -202.430 414.095 -200.890 ;
        RECT 411.805 -202.645 412.160 -202.640 ;
        RECT 413.865 -202.645 414.235 -202.615 ;
        RECT 411.805 -202.650 414.235 -202.645 ;
        RECT 409.060 -202.820 414.235 -202.650 ;
        RECT 416.020 -202.755 416.325 -200.720 ;
        RECT 409.065 -202.840 414.235 -202.820 ;
        RECT 409.065 -202.850 411.810 -202.840 ;
        RECT 407.000 -202.990 407.365 -202.960 ;
        RECT 413.865 -202.970 414.235 -202.840 ;
        RECT 406.105 -203.075 407.365 -202.990 ;
        RECT 406.130 -203.195 407.365 -203.075 ;
        RECT 411.540 -203.130 412.215 -203.090 ;
        RECT 411.440 -203.140 412.215 -203.130 ;
        RECT 406.130 -203.280 406.780 -203.195 ;
        RECT 407.000 -203.260 407.365 -203.195 ;
        RECT 410.405 -203.320 412.215 -203.140 ;
        RECT 414.800 -203.185 418.725 -202.755 ;
        RECT 411.440 -203.330 412.215 -203.320 ;
        RECT 411.540 -203.360 412.215 -203.330 ;
        RECT 412.455 -203.245 414.550 -203.205 ;
        RECT 412.455 -203.395 414.605 -203.245 ;
        RECT 407.590 -204.470 407.760 -203.430 ;
        RECT 408.570 -204.470 408.740 -203.430 ;
        RECT 409.550 -204.470 409.720 -203.430 ;
        RECT 412.455 -205.115 412.625 -203.395 ;
        RECT 413.435 -205.115 413.605 -203.395 ;
        RECT 414.300 -204.140 414.605 -203.395 ;
        RECT 415.500 -203.965 415.670 -203.185 ;
        RECT 415.990 -203.965 416.160 -203.425 ;
        RECT 416.480 -203.965 416.650 -203.185 ;
        RECT 416.970 -203.965 417.140 -203.425 ;
        RECT 414.910 -204.140 415.275 -204.110 ;
        RECT 414.300 -204.205 415.275 -204.140 ;
        RECT 414.410 -204.345 415.275 -204.205 ;
        RECT 414.910 -204.410 415.275 -204.345 ;
        RECT 417.460 -204.260 419.320 -203.910 ;
        RECT 415.500 -205.120 415.670 -204.580 ;
        RECT 416.480 -205.120 416.650 -204.580 ;
        RECT 417.460 -205.120 417.630 -204.260 ;
        RECT 415.730 -207.460 416.930 -207.290 ;
        RECT 407.460 -209.795 407.630 -208.075 ;
        RECT 408.440 -209.795 408.610 -208.075 ;
        RECT 410.505 -208.610 410.675 -208.070 ;
        RECT 411.485 -208.610 411.655 -208.070 ;
        RECT 409.915 -208.845 410.280 -208.780 ;
        RECT 409.415 -208.985 410.280 -208.845 ;
        RECT 409.305 -209.050 410.280 -208.985 ;
        RECT 409.305 -209.795 409.610 -209.050 ;
        RECT 409.915 -209.080 410.280 -209.050 ;
        RECT 412.465 -208.930 412.635 -208.070 ;
        RECT 406.545 -209.860 407.220 -209.830 ;
        RECT 406.445 -209.870 407.220 -209.860 ;
        RECT 403.805 -210.050 407.220 -209.870 ;
        RECT 407.460 -209.945 409.610 -209.795 ;
        RECT 407.460 -209.985 409.555 -209.945 ;
        RECT 410.505 -210.005 410.675 -209.225 ;
        RECT 410.995 -209.765 411.165 -209.225 ;
        RECT 411.485 -210.005 411.655 -209.225 ;
        RECT 411.975 -209.765 412.145 -209.225 ;
        RECT 412.465 -209.280 413.855 -208.930 ;
        RECT 404.720 -215.185 405.400 -210.050 ;
        RECT 406.445 -210.060 407.220 -210.050 ;
        RECT 406.545 -210.100 407.220 -210.060 ;
        RECT 405.680 -210.350 406.815 -210.340 ;
        RECT 408.870 -210.350 409.240 -210.220 ;
        RECT 405.680 -210.540 409.240 -210.350 ;
        RECT 409.805 -210.435 412.880 -210.005 ;
        RECT 406.810 -210.545 409.240 -210.540 ;
        RECT 406.810 -210.550 407.165 -210.545 ;
        RECT 408.870 -210.575 409.240 -210.545 ;
        RECT 406.970 -212.300 407.140 -210.760 ;
        RECT 407.460 -212.300 407.630 -210.760 ;
        RECT 407.950 -212.300 408.120 -210.760 ;
        RECT 408.440 -212.300 408.610 -210.760 ;
        RECT 408.930 -212.300 409.100 -210.760 ;
        RECT 407.455 -212.560 407.630 -212.300 ;
        RECT 411.025 -212.470 411.330 -210.435 ;
        RECT 413.475 -211.255 413.825 -209.280 ;
        RECT 414.695 -210.550 414.865 -207.630 ;
        RECT 415.730 -207.670 415.940 -207.460 ;
        RECT 414.675 -210.845 414.885 -210.550 ;
        RECT 415.750 -210.580 415.920 -207.670 ;
        RECT 416.240 -210.570 416.410 -207.630 ;
        RECT 416.720 -207.680 416.930 -207.460 ;
        RECT 415.735 -210.845 415.945 -210.580 ;
        RECT 414.675 -211.025 415.945 -210.845 ;
        RECT 416.220 -210.840 416.430 -210.570 ;
        RECT 416.730 -210.670 416.900 -207.680 ;
        RECT 417.790 -210.600 417.960 -207.630 ;
        RECT 416.220 -211.035 416.925 -210.840 ;
        RECT 416.710 -211.095 416.925 -211.035 ;
        RECT 415.500 -211.255 416.275 -211.205 ;
        RECT 413.475 -211.435 416.275 -211.255 ;
        RECT 413.475 -211.445 413.825 -211.435 ;
        RECT 415.500 -211.480 416.275 -211.435 ;
        RECT 416.710 -211.370 417.615 -211.095 ;
        RECT 416.710 -211.720 416.925 -211.370 ;
        RECT 414.150 -211.790 414.925 -211.745 ;
        RECT 413.965 -211.960 414.925 -211.790 ;
        RECT 414.150 -212.020 414.925 -211.960 ;
        RECT 415.155 -211.920 416.925 -211.720 ;
        RECT 417.785 -211.820 418.000 -210.600 ;
        RECT 418.970 -210.945 419.320 -204.260 ;
        RECT 420.310 -210.575 420.525 -200.700 ;
        RECT 421.945 -202.815 422.325 -199.295 ;
        RECT 423.455 -199.075 432.390 -198.885 ;
        RECT 423.455 -200.965 423.645 -199.075 ;
        RECT 429.490 -200.570 432.815 -200.430 ;
        RECT 429.490 -200.860 434.665 -200.570 ;
        RECT 423.340 -201.235 423.705 -200.965 ;
        RECT 429.490 -201.265 429.920 -200.860 ;
        RECT 430.790 -201.045 430.965 -200.860 ;
        RECT 432.415 -200.875 434.665 -200.860 ;
        RECT 425.230 -201.695 429.920 -201.265 ;
        RECT 424.470 -202.815 425.120 -202.685 ;
        RECT 421.945 -203.145 425.120 -202.815 ;
        RECT 425.930 -202.975 426.100 -201.695 ;
        RECT 426.420 -202.975 426.590 -201.935 ;
        RECT 426.910 -202.975 427.080 -201.695 ;
        RECT 427.400 -202.805 427.570 -201.935 ;
        RECT 430.305 -202.585 430.475 -201.045 ;
        RECT 430.795 -202.585 430.965 -201.045 ;
        RECT 431.285 -202.585 431.455 -201.045 ;
        RECT 431.775 -202.585 431.945 -201.045 ;
        RECT 432.265 -202.585 432.435 -201.045 ;
        RECT 430.145 -202.800 430.500 -202.795 ;
        RECT 432.205 -202.800 432.575 -202.770 ;
        RECT 430.145 -202.805 432.575 -202.800 ;
        RECT 427.400 -202.975 432.575 -202.805 ;
        RECT 434.360 -202.910 434.665 -200.875 ;
        RECT 427.405 -202.995 432.575 -202.975 ;
        RECT 427.405 -203.005 430.150 -202.995 ;
        RECT 425.340 -203.145 425.705 -203.115 ;
        RECT 432.205 -203.125 432.575 -202.995 ;
        RECT 421.945 -203.195 425.705 -203.145 ;
        RECT 424.470 -203.350 425.705 -203.195 ;
        RECT 429.880 -203.285 430.555 -203.245 ;
        RECT 429.780 -203.295 430.555 -203.285 ;
        RECT 424.470 -203.435 425.120 -203.350 ;
        RECT 425.340 -203.415 425.705 -203.350 ;
        RECT 424.605 -203.685 424.985 -203.435 ;
        RECT 428.745 -203.475 430.555 -203.295 ;
        RECT 433.140 -203.340 437.065 -202.910 ;
        RECT 429.780 -203.485 430.555 -203.475 ;
        RECT 429.880 -203.515 430.555 -203.485 ;
        RECT 430.795 -203.400 432.890 -203.360 ;
        RECT 430.795 -203.550 432.945 -203.400 ;
        RECT 425.930 -204.625 426.100 -203.585 ;
        RECT 426.910 -204.625 427.080 -203.585 ;
        RECT 427.890 -204.625 428.060 -203.585 ;
        RECT 430.795 -205.270 430.965 -203.550 ;
        RECT 431.775 -205.270 431.945 -203.550 ;
        RECT 432.640 -204.295 432.945 -203.550 ;
        RECT 433.840 -204.120 434.010 -203.340 ;
        RECT 434.330 -204.120 434.500 -203.580 ;
        RECT 434.820 -204.120 434.990 -203.340 ;
        RECT 435.310 -204.120 435.480 -203.580 ;
        RECT 433.250 -204.295 433.615 -204.265 ;
        RECT 432.640 -204.360 433.615 -204.295 ;
        RECT 432.750 -204.500 433.615 -204.360 ;
        RECT 433.250 -204.565 433.615 -204.500 ;
        RECT 435.800 -204.415 437.660 -204.065 ;
        RECT 433.840 -205.275 434.010 -204.735 ;
        RECT 434.820 -205.275 434.990 -204.735 ;
        RECT 435.800 -205.275 435.970 -204.415 ;
        RECT 434.070 -207.615 435.270 -207.445 ;
        RECT 425.800 -209.950 425.970 -208.230 ;
        RECT 426.780 -209.950 426.950 -208.230 ;
        RECT 428.845 -208.765 429.015 -208.225 ;
        RECT 429.825 -208.765 429.995 -208.225 ;
        RECT 428.255 -209.000 428.620 -208.935 ;
        RECT 427.755 -209.140 428.620 -209.000 ;
        RECT 427.645 -209.205 428.620 -209.140 ;
        RECT 427.645 -209.950 427.950 -209.205 ;
        RECT 428.255 -209.235 428.620 -209.205 ;
        RECT 430.805 -209.085 430.975 -208.225 ;
        RECT 424.885 -210.015 425.560 -209.985 ;
        RECT 424.785 -210.025 425.560 -210.015 ;
        RECT 422.715 -210.205 425.560 -210.025 ;
        RECT 425.800 -210.100 427.950 -209.950 ;
        RECT 425.800 -210.140 427.895 -210.100 ;
        RECT 428.845 -210.160 429.015 -209.380 ;
        RECT 429.335 -209.920 429.505 -209.380 ;
        RECT 429.825 -210.160 429.995 -209.380 ;
        RECT 430.315 -209.920 430.485 -209.380 ;
        RECT 430.805 -209.435 432.195 -209.085 ;
        RECT 420.310 -210.790 421.735 -210.575 ;
        RECT 418.915 -211.305 419.440 -210.945 ;
        RECT 421.520 -211.820 421.735 -210.790 ;
        RECT 409.080 -212.560 411.330 -212.470 ;
        RECT 406.870 -212.775 411.330 -212.560 ;
        RECT 406.870 -212.865 409.115 -212.775 ;
        RECT 411.025 -214.250 411.330 -212.775 ;
        RECT 414.695 -213.660 414.865 -212.190 ;
        RECT 415.155 -212.270 415.380 -211.920 ;
        RECT 417.115 -212.020 421.735 -211.820 ;
        RECT 417.355 -212.035 421.735 -212.020 ;
        RECT 414.660 -214.250 414.895 -213.660 ;
        RECT 415.185 -213.730 415.355 -212.270 ;
        RECT 415.675 -213.655 415.845 -212.190 ;
        RECT 416.885 -213.605 417.055 -212.190 ;
        RECT 417.355 -212.235 417.575 -212.035 ;
        RECT 415.640 -214.250 415.875 -213.655 ;
        RECT 416.850 -214.250 417.085 -213.605 ;
        RECT 417.375 -213.730 417.545 -212.235 ;
        RECT 411.025 -214.815 418.410 -214.250 ;
        RECT 422.715 -215.185 423.395 -210.205 ;
        RECT 424.785 -210.215 425.560 -210.205 ;
        RECT 424.885 -210.255 425.560 -210.215 ;
        RECT 424.020 -210.505 425.155 -210.495 ;
        RECT 427.210 -210.505 427.580 -210.375 ;
        RECT 424.020 -210.695 427.580 -210.505 ;
        RECT 428.145 -210.590 431.220 -210.160 ;
        RECT 425.150 -210.700 427.580 -210.695 ;
        RECT 425.150 -210.705 425.505 -210.700 ;
        RECT 427.210 -210.730 427.580 -210.700 ;
        RECT 425.310 -212.455 425.480 -210.915 ;
        RECT 425.800 -212.455 425.970 -210.915 ;
        RECT 426.290 -212.455 426.460 -210.915 ;
        RECT 426.780 -212.455 426.950 -210.915 ;
        RECT 427.270 -212.455 427.440 -210.915 ;
        RECT 425.795 -212.715 425.970 -212.455 ;
        RECT 429.365 -212.625 429.670 -210.590 ;
        RECT 431.815 -211.410 432.165 -209.435 ;
        RECT 433.035 -210.705 433.205 -207.785 ;
        RECT 434.070 -207.825 434.280 -207.615 ;
        RECT 433.015 -211.000 433.225 -210.705 ;
        RECT 434.090 -210.735 434.260 -207.825 ;
        RECT 434.580 -210.725 434.750 -207.785 ;
        RECT 435.060 -207.835 435.270 -207.615 ;
        RECT 434.075 -211.000 434.285 -210.735 ;
        RECT 433.015 -211.180 434.285 -211.000 ;
        RECT 434.560 -210.995 434.770 -210.725 ;
        RECT 435.070 -210.825 435.240 -207.835 ;
        RECT 436.130 -210.755 436.300 -207.785 ;
        RECT 434.560 -211.190 435.265 -210.995 ;
        RECT 435.050 -211.250 435.265 -211.190 ;
        RECT 433.840 -211.410 434.615 -211.360 ;
        RECT 431.815 -211.590 434.615 -211.410 ;
        RECT 431.815 -211.600 432.165 -211.590 ;
        RECT 433.840 -211.635 434.615 -211.590 ;
        RECT 435.050 -211.525 435.955 -211.250 ;
        RECT 435.050 -211.875 435.265 -211.525 ;
        RECT 432.490 -211.945 433.265 -211.900 ;
        RECT 432.305 -212.115 433.265 -211.945 ;
        RECT 432.490 -212.175 433.265 -212.115 ;
        RECT 433.495 -212.075 435.265 -211.875 ;
        RECT 436.125 -211.975 436.340 -210.755 ;
        RECT 437.310 -211.100 437.660 -204.415 ;
        RECT 437.255 -211.460 437.780 -211.100 ;
        RECT 440.400 -211.975 442.195 -211.225 ;
        RECT 427.420 -212.715 429.670 -212.625 ;
        RECT 425.210 -212.930 429.670 -212.715 ;
        RECT 425.210 -213.020 427.455 -212.930 ;
        RECT 429.365 -214.405 429.670 -212.930 ;
        RECT 433.035 -213.815 433.205 -212.345 ;
        RECT 433.495 -212.425 433.720 -212.075 ;
        RECT 435.455 -212.175 442.195 -211.975 ;
        RECT 435.695 -212.190 442.195 -212.175 ;
        RECT 433.000 -214.405 433.235 -213.815 ;
        RECT 433.525 -213.885 433.695 -212.425 ;
        RECT 434.015 -213.810 434.185 -212.345 ;
        RECT 435.225 -213.760 435.395 -212.345 ;
        RECT 435.695 -212.390 435.915 -212.190 ;
        RECT 433.980 -214.405 434.215 -213.810 ;
        RECT 435.190 -214.405 435.425 -213.760 ;
        RECT 435.715 -213.885 435.885 -212.390 ;
        RECT 440.400 -212.940 442.195 -212.190 ;
        RECT 429.365 -214.970 436.750 -214.405 ;
        RECT 404.720 -215.865 423.395 -215.185 ;
        RECT 401.515 -223.700 403.450 -222.320 ;
        RECT -121.070 -229.560 358.580 -228.880 ;
        RECT -121.070 -230.730 -120.390 -229.560 ;
        RECT 404.840 -230.730 405.520 -215.865 ;
        RECT -121.070 -231.410 405.520 -230.730 ;
        RECT -36.545 -233.930 88.175 -233.250 ;
        RECT -120.295 -235.115 55.545 -234.440 ;
        RECT -147.240 -274.555 -145.890 -273.805 ;
        RECT -144.245 -274.555 -143.645 -261.155 ;
        RECT -141.180 -261.310 -140.720 -261.180 ;
        RECT -143.220 -261.480 -140.720 -261.310 ;
        RECT -141.180 -261.900 -140.720 -261.480 ;
        RECT -143.220 -262.070 -140.720 -261.900 ;
        RECT -141.180 -262.490 -140.720 -262.070 ;
        RECT -143.220 -262.660 -140.720 -262.490 ;
        RECT -141.180 -263.080 -140.720 -262.660 ;
        RECT -143.220 -263.250 -140.720 -263.080 ;
        RECT -141.180 -263.670 -140.720 -263.250 ;
        RECT -143.220 -263.840 -140.720 -263.670 ;
        RECT -141.180 -264.260 -140.720 -263.840 ;
        RECT -143.220 -264.430 -140.720 -264.260 ;
        RECT -141.180 -264.850 -140.720 -264.430 ;
        RECT -143.220 -265.020 -140.720 -264.850 ;
        RECT -141.180 -265.440 -140.720 -265.020 ;
        RECT 44.720 -261.565 101.060 -259.900 ;
        RECT -143.220 -265.610 -140.720 -265.440 ;
        RECT -60.965 -265.380 -57.825 -265.210 ;
        RECT -68.200 -265.495 -68.030 -265.475 ;
        RECT -141.180 -266.030 -140.720 -265.610 ;
        RECT -143.220 -266.200 -140.720 -266.030 ;
        RECT -141.180 -266.620 -140.720 -266.200 ;
        RECT -143.220 -266.790 -140.720 -266.620 ;
        RECT -141.180 -267.210 -140.720 -266.790 ;
        RECT -68.230 -266.760 -68.000 -265.495 ;
        RECT -67.220 -266.435 -67.050 -265.475 ;
        RECT -66.240 -266.435 -66.070 -265.475 ;
        RECT -64.015 -265.495 -63.845 -265.475 ;
        RECT -65.120 -265.905 -64.835 -265.585 ;
        RECT -65.835 -266.150 -64.835 -265.905 ;
        RECT -67.250 -266.760 -67.020 -266.435 ;
        RECT -66.270 -266.760 -66.040 -266.435 ;
        RECT -68.230 -266.800 -66.040 -266.760 ;
        RECT -65.835 -266.800 -65.605 -266.150 ;
        RECT -65.120 -266.405 -64.835 -266.150 ;
        RECT -69.250 -266.985 -68.410 -266.835 ;
        RECT -143.220 -267.380 -140.720 -267.210 ;
        RECT -141.180 -267.800 -140.720 -267.380 ;
        RECT -143.220 -267.970 -140.720 -267.800 ;
        RECT -141.180 -268.390 -140.720 -267.970 ;
        RECT -143.220 -268.560 -140.720 -268.390 ;
        RECT -141.180 -268.980 -140.720 -268.560 ;
        RECT -143.220 -269.150 -140.720 -268.980 ;
        RECT -69.285 -267.205 -68.410 -266.985 ;
        RECT -68.230 -266.990 -65.605 -266.800 ;
        RECT -64.045 -266.760 -63.815 -265.495 ;
        RECT -63.035 -266.435 -62.865 -265.475 ;
        RECT -62.055 -266.435 -61.885 -265.475 ;
        RECT -60.965 -265.605 -60.785 -265.380 ;
        RECT -63.065 -266.760 -62.835 -266.435 ;
        RECT -62.085 -266.760 -61.855 -266.435 ;
        RECT -64.045 -266.800 -61.855 -266.760 ;
        RECT -61.580 -266.680 -61.210 -265.840 ;
        RECT -60.960 -265.975 -60.790 -265.605 ;
        RECT -61.580 -266.800 -61.215 -266.680 ;
        RECT -65.065 -266.890 -64.225 -266.835 ;
        RECT -65.240 -266.895 -64.225 -266.890 ;
        RECT -69.285 -269.065 -69.045 -267.205 ;
        RECT -68.690 -268.170 -68.520 -267.375 ;
        RECT -68.230 -267.455 -68.000 -266.990 ;
        RECT -68.200 -267.915 -68.030 -267.455 ;
        RECT -67.710 -268.170 -67.540 -267.375 ;
        RECT -67.250 -267.455 -67.020 -266.990 ;
        RECT -66.270 -267.150 -65.605 -266.990 ;
        RECT -67.220 -267.915 -67.050 -267.455 ;
        RECT -66.730 -268.170 -66.560 -267.375 ;
        RECT -66.270 -267.455 -66.040 -267.150 ;
        RECT -65.425 -267.205 -64.225 -266.895 ;
        RECT -64.045 -266.990 -61.215 -266.800 ;
        RECT -66.240 -267.915 -66.070 -267.455 ;
        RECT -65.425 -267.925 -65.125 -267.205 ;
        RECT -64.505 -268.170 -64.335 -267.375 ;
        RECT -64.045 -267.455 -63.815 -266.990 ;
        RECT -64.015 -267.915 -63.845 -267.455 ;
        RECT -63.525 -268.170 -63.355 -267.375 ;
        RECT -63.065 -267.455 -62.835 -266.990 ;
        RECT -62.085 -267.150 -61.215 -266.990 ;
        RECT -60.990 -266.710 -60.755 -265.975 ;
        RECT -60.470 -266.010 -60.300 -265.550 ;
        RECT -59.985 -265.655 -59.775 -265.380 ;
        RECT -60.475 -266.270 -60.295 -266.010 ;
        RECT -59.980 -266.090 -59.810 -265.655 ;
        RECT -59.490 -266.000 -59.320 -265.550 ;
        RECT -59.015 -265.660 -58.805 -265.380 ;
        RECT -59.490 -266.090 -59.305 -266.000 ;
        RECT -59.000 -266.090 -58.830 -265.660 ;
        RECT -58.510 -266.000 -58.340 -265.550 ;
        RECT -58.035 -265.635 -57.825 -265.380 ;
        RECT -47.465 -265.380 -44.325 -265.210 ;
        RECT -54.700 -265.495 -54.530 -265.475 ;
        RECT -59.485 -266.270 -59.305 -266.090 ;
        RECT -58.515 -266.270 -58.335 -266.000 ;
        RECT -58.020 -266.090 -57.850 -265.635 ;
        RECT -57.530 -266.050 -57.360 -265.550 ;
        RECT -57.545 -266.270 -57.335 -266.050 ;
        RECT -60.475 -266.440 -57.335 -266.270 ;
        RECT -60.990 -267.080 -60.130 -266.710 ;
        RECT -58.210 -266.975 -57.335 -266.440 ;
        RECT -54.730 -266.760 -54.500 -265.495 ;
        RECT -53.720 -266.435 -53.550 -265.475 ;
        RECT -52.740 -266.435 -52.570 -265.475 ;
        RECT -50.515 -265.495 -50.345 -265.475 ;
        RECT -51.620 -265.845 -51.335 -265.585 ;
        RECT -52.360 -266.155 -51.335 -265.845 ;
        RECT -53.750 -266.760 -53.520 -266.435 ;
        RECT -52.770 -266.760 -52.540 -266.435 ;
        RECT -54.730 -266.800 -52.540 -266.760 ;
        RECT -52.360 -266.800 -52.050 -266.155 ;
        RECT -51.620 -266.405 -51.335 -266.155 ;
        RECT -55.750 -266.870 -54.910 -266.835 ;
        RECT -63.035 -267.915 -62.865 -267.455 ;
        RECT -62.545 -268.170 -62.375 -267.375 ;
        RECT -62.085 -267.455 -61.855 -267.150 ;
        RECT -62.055 -267.915 -61.885 -267.455 ;
        RECT -60.990 -267.755 -60.755 -267.080 ;
        RECT -58.210 -267.275 -56.880 -266.975 ;
        RECT -55.860 -267.170 -54.910 -266.870 ;
        RECT -55.750 -267.205 -54.910 -267.170 ;
        RECT -54.730 -266.990 -52.050 -266.800 ;
        RECT -50.545 -266.760 -50.315 -265.495 ;
        RECT -49.535 -266.435 -49.365 -265.475 ;
        RECT -48.555 -266.435 -48.385 -265.475 ;
        RECT -47.465 -265.605 -47.285 -265.380 ;
        RECT -49.565 -266.760 -49.335 -266.435 ;
        RECT -48.585 -266.760 -48.355 -266.435 ;
        RECT -50.545 -266.800 -48.355 -266.760 ;
        RECT -48.080 -266.680 -47.710 -265.840 ;
        RECT -47.460 -265.975 -47.290 -265.605 ;
        RECT -48.080 -266.800 -47.715 -266.680 ;
        RECT -51.565 -266.890 -50.725 -266.835 ;
        RECT -60.490 -267.445 -57.335 -267.275 ;
        RECT -60.490 -267.650 -60.285 -267.445 ;
        RECT -60.960 -268.105 -60.790 -267.755 ;
        RECT -68.735 -268.510 -61.880 -268.170 ;
        RECT -60.985 -268.395 -60.765 -268.105 ;
        RECT -60.470 -268.165 -60.300 -267.650 ;
        RECT -59.980 -268.050 -59.810 -267.625 ;
        RECT -59.500 -267.690 -59.295 -267.445 ;
        RECT -60.005 -268.395 -59.785 -268.050 ;
        RECT -59.490 -268.165 -59.320 -267.690 ;
        RECT -59.000 -268.050 -58.830 -267.625 ;
        RECT -58.530 -267.690 -58.325 -267.445 ;
        RECT -57.545 -267.480 -57.335 -267.445 ;
        RECT -59.025 -268.395 -58.805 -268.050 ;
        RECT -58.510 -268.165 -58.340 -267.690 ;
        RECT -58.020 -268.105 -57.850 -267.625 ;
        RECT -57.545 -267.695 -57.340 -267.480 ;
        RECT -58.040 -268.395 -57.820 -268.105 ;
        RECT -57.530 -268.165 -57.360 -267.695 ;
        RECT -55.190 -268.170 -55.020 -267.375 ;
        RECT -54.730 -267.455 -54.500 -266.990 ;
        RECT -54.700 -267.915 -54.530 -267.455 ;
        RECT -54.210 -268.170 -54.040 -267.375 ;
        RECT -53.750 -267.455 -53.520 -266.990 ;
        RECT -52.770 -267.150 -52.050 -266.990 ;
        RECT -53.720 -267.915 -53.550 -267.455 ;
        RECT -53.230 -268.170 -53.060 -267.375 ;
        RECT -52.770 -267.455 -52.540 -267.150 ;
        RECT -51.865 -267.205 -50.725 -266.890 ;
        RECT -50.545 -266.990 -47.715 -266.800 ;
        RECT -52.740 -267.915 -52.570 -267.455 ;
        RECT -51.865 -268.000 -51.565 -267.205 ;
        RECT -51.005 -268.170 -50.835 -267.375 ;
        RECT -50.545 -267.455 -50.315 -266.990 ;
        RECT -50.515 -267.915 -50.345 -267.455 ;
        RECT -50.025 -268.170 -49.855 -267.375 ;
        RECT -49.565 -267.455 -49.335 -266.990 ;
        RECT -48.585 -267.150 -47.715 -266.990 ;
        RECT -47.490 -266.710 -47.255 -265.975 ;
        RECT -46.970 -266.010 -46.800 -265.550 ;
        RECT -46.485 -265.655 -46.275 -265.380 ;
        RECT -46.975 -266.270 -46.795 -266.010 ;
        RECT -46.480 -266.090 -46.310 -265.655 ;
        RECT -45.990 -266.000 -45.820 -265.550 ;
        RECT -45.515 -265.660 -45.305 -265.380 ;
        RECT -45.990 -266.090 -45.805 -266.000 ;
        RECT -45.500 -266.090 -45.330 -265.660 ;
        RECT -45.010 -266.000 -44.840 -265.550 ;
        RECT -44.535 -265.635 -44.325 -265.380 ;
        RECT -36.340 -265.355 -35.140 -265.185 ;
        RECT -45.985 -266.270 -45.805 -266.090 ;
        RECT -45.015 -266.270 -44.835 -266.000 ;
        RECT -44.520 -266.090 -44.350 -265.635 ;
        RECT -44.030 -266.050 -43.860 -265.550 ;
        RECT -44.045 -266.270 -43.835 -266.050 ;
        RECT -46.975 -266.440 -43.835 -266.270 ;
        RECT -47.490 -267.080 -46.630 -266.710 ;
        RECT -44.710 -266.985 -43.835 -266.440 ;
        RECT -49.535 -267.915 -49.365 -267.455 ;
        RECT -49.045 -268.170 -48.875 -267.375 ;
        RECT -48.585 -267.455 -48.355 -267.150 ;
        RECT -48.555 -267.915 -48.385 -267.455 ;
        RECT -47.490 -267.755 -47.255 -267.080 ;
        RECT -44.710 -267.275 -43.460 -266.985 ;
        RECT -46.990 -267.285 -43.460 -267.275 ;
        RECT -46.990 -267.445 -43.835 -267.285 ;
        RECT -46.990 -267.650 -46.785 -267.445 ;
        RECT -47.460 -268.105 -47.290 -267.755 ;
        RECT -67.495 -268.710 -66.940 -268.510 ;
        RECT -67.550 -268.750 -66.865 -268.710 ;
        RECT -63.440 -268.750 -62.885 -268.510 ;
        RECT -60.985 -268.565 -57.820 -268.395 ;
        RECT -55.235 -268.180 -52.565 -268.170 ;
        RECT -51.050 -268.180 -48.380 -268.170 ;
        RECT -55.235 -268.510 -48.380 -268.180 ;
        RECT -47.485 -268.395 -47.265 -268.105 ;
        RECT -46.970 -268.165 -46.800 -267.650 ;
        RECT -46.480 -268.050 -46.310 -267.625 ;
        RECT -46.000 -267.690 -45.795 -267.445 ;
        RECT -46.505 -268.395 -46.285 -268.050 ;
        RECT -45.990 -268.165 -45.820 -267.690 ;
        RECT -45.500 -268.050 -45.330 -267.625 ;
        RECT -45.030 -267.690 -44.825 -267.445 ;
        RECT -44.045 -267.480 -43.835 -267.445 ;
        RECT -45.525 -268.395 -45.305 -268.050 ;
        RECT -45.010 -268.165 -44.840 -267.690 ;
        RECT -44.520 -268.105 -44.350 -267.625 ;
        RECT -44.045 -267.695 -43.840 -267.480 ;
        RECT -44.540 -268.395 -44.320 -268.105 ;
        RECT -44.030 -268.165 -43.860 -267.695 ;
        RECT -54.450 -268.740 -53.895 -268.510 ;
        RECT -53.535 -268.520 -50.935 -268.510 ;
        RECT -54.565 -268.750 -53.880 -268.740 ;
        RECT -50.060 -268.750 -49.505 -268.510 ;
        RECT -47.485 -268.565 -44.320 -268.395 ;
        RECT -37.370 -268.495 -37.200 -265.525 ;
        RECT -36.340 -265.575 -36.130 -265.355 ;
        RECT -41.375 -268.750 -40.715 -268.740 ;
        RECT -67.635 -268.945 -40.710 -268.750 ;
        RECT -67.550 -269.010 -66.865 -268.945 ;
        RECT -54.565 -269.040 -53.880 -268.945 ;
        RECT -41.375 -269.040 -40.715 -268.945 ;
        RECT -141.180 -269.570 -140.720 -269.150 ;
        RECT -143.220 -269.740 -140.720 -269.570 ;
        RECT -141.180 -270.160 -140.720 -269.740 ;
        RECT -143.220 -270.330 -140.720 -270.160 ;
        RECT -141.180 -270.750 -140.720 -270.330 ;
        RECT -143.220 -270.920 -140.720 -270.750 ;
        RECT -106.195 -270.630 -106.025 -269.410 ;
        RECT -105.215 -270.630 -105.045 -269.410 ;
        RECT -104.235 -270.630 -104.065 -269.410 ;
        RECT -106.195 -270.815 -103.420 -270.630 ;
        RECT -141.180 -271.340 -140.720 -270.920 ;
        RECT -143.220 -271.510 -140.720 -271.340 ;
        RECT -141.180 -271.930 -140.720 -271.510 ;
        RECT -143.220 -272.100 -140.720 -271.930 ;
        RECT -103.605 -271.505 -103.420 -270.815 ;
        RECT -101.395 -271.505 -100.720 -271.455 ;
        RECT -103.605 -271.690 -100.720 -271.505 ;
        RECT -103.605 -271.960 -103.420 -271.690 ;
        RECT -101.395 -271.725 -100.720 -271.690 ;
        RECT -141.180 -272.520 -140.720 -272.100 ;
        RECT -143.220 -272.690 -140.720 -272.520 ;
        RECT -141.180 -273.110 -140.720 -272.690 ;
        RECT -143.220 -273.280 -140.720 -273.110 ;
        RECT -141.180 -273.700 -140.720 -273.280 ;
        RECT -143.220 -273.870 -140.720 -273.700 ;
        RECT -141.180 -274.290 -140.720 -273.870 ;
        RECT -106.685 -272.130 -104.470 -271.960 ;
        RECT -103.605 -272.130 -102.440 -271.960 ;
        RECT -106.685 -273.985 -106.515 -272.130 ;
        RECT -105.705 -272.135 -104.470 -272.130 ;
        RECT -143.220 -274.460 -140.720 -274.290 ;
        RECT -147.240 -275.945 -143.645 -274.555 ;
        RECT -141.180 -274.880 -140.720 -274.460 ;
        RECT -143.220 -275.050 -140.720 -274.880 ;
        RECT -106.195 -274.930 -106.025 -272.445 ;
        RECT -105.705 -273.985 -105.535 -272.135 ;
        RECT -104.645 -272.450 -104.470 -272.135 ;
        RECT -105.135 -273.945 -104.965 -272.450 ;
        RECT -105.135 -274.465 -104.960 -273.945 ;
        RECT -104.645 -273.990 -104.475 -272.450 ;
        RECT -104.155 -273.935 -103.985 -272.450 ;
        RECT -104.155 -274.465 -103.980 -273.935 ;
        RECT -103.590 -273.990 -103.420 -272.130 ;
        RECT -105.135 -274.480 -103.980 -274.465 ;
        RECT -103.100 -274.480 -102.930 -272.450 ;
        RECT -102.610 -273.990 -102.440 -272.130 ;
        RECT -105.135 -274.650 -102.930 -274.480 ;
        RECT -101.035 -274.485 -100.865 -272.950 ;
        RECT -100.545 -273.990 -100.375 -269.410 ;
        RECT -98.265 -271.815 -97.580 -271.730 ;
        RECT -96.200 -271.740 -96.030 -270.020 ;
        RECT -95.220 -271.740 -95.050 -270.020 ;
        RECT -93.155 -270.555 -92.985 -270.015 ;
        RECT -92.175 -270.555 -92.005 -270.015 ;
        RECT -93.745 -270.790 -93.380 -270.725 ;
        RECT -94.245 -270.930 -93.380 -270.790 ;
        RECT -94.355 -270.995 -93.380 -270.930 ;
        RECT -94.355 -271.740 -94.050 -270.995 ;
        RECT -93.745 -271.025 -93.380 -270.995 ;
        RECT -91.195 -270.875 -91.025 -270.015 ;
        RECT -84.455 -270.195 -77.070 -269.630 ;
        RECT -69.290 -269.750 -68.990 -269.065 ;
        RECT -56.740 -269.210 -56.055 -269.155 ;
        RECT -52.010 -269.210 -51.350 -269.160 ;
        RECT -67.635 -269.405 -38.985 -269.210 ;
        RECT -56.740 -269.455 -56.055 -269.405 ;
        RECT -52.010 -269.460 -51.350 -269.405 ;
        RECT -65.605 -269.640 -64.945 -269.600 ;
        RECT -42.990 -269.640 -42.330 -269.590 ;
        RECT -91.195 -270.880 -89.175 -270.875 ;
        RECT -91.195 -271.170 -88.855 -270.880 ;
        RECT -97.115 -271.805 -96.440 -271.775 ;
        RECT -97.215 -271.815 -96.440 -271.805 ;
        RECT -98.265 -271.995 -96.440 -271.815 ;
        RECT -96.200 -271.890 -94.050 -271.740 ;
        RECT -96.200 -271.930 -94.105 -271.890 ;
        RECT -93.155 -271.950 -92.985 -271.170 ;
        RECT -92.665 -271.710 -92.495 -271.170 ;
        RECT -92.175 -271.950 -92.005 -271.170 ;
        RECT -91.685 -271.710 -91.515 -271.170 ;
        RECT -91.195 -271.225 -89.175 -271.170 ;
        RECT -88.610 -271.670 -86.365 -271.580 ;
        RECT -84.455 -271.670 -84.150 -270.195 ;
        RECT -80.820 -270.785 -80.585 -270.195 ;
        RECT -90.990 -271.950 -84.150 -271.670 ;
        RECT -98.265 -272.020 -97.580 -271.995 ;
        RECT -97.215 -272.005 -96.440 -271.995 ;
        RECT -97.115 -272.045 -96.440 -272.005 ;
        RECT -93.855 -271.975 -84.150 -271.950 ;
        RECT -93.855 -272.380 -90.685 -271.975 ;
        RECT -88.025 -272.145 -87.850 -271.975 ;
        RECT -96.690 -274.245 -96.520 -272.705 ;
        RECT -96.200 -274.245 -96.030 -272.705 ;
        RECT -95.710 -274.245 -95.540 -272.705 ;
        RECT -95.220 -274.245 -95.050 -272.705 ;
        RECT -94.730 -274.245 -94.560 -272.705 ;
        RECT -96.205 -274.485 -96.030 -274.245 ;
        RECT -92.635 -274.415 -92.330 -272.380 ;
        RECT -90.990 -272.390 -90.685 -272.380 ;
        RECT -88.510 -273.685 -88.340 -272.145 ;
        RECT -88.020 -273.685 -87.850 -272.145 ;
        RECT -87.530 -273.685 -87.360 -272.145 ;
        RECT -87.040 -273.685 -86.870 -272.145 ;
        RECT -86.550 -273.685 -86.380 -272.145 ;
        RECT -88.670 -273.900 -88.315 -273.895 ;
        RECT -86.610 -273.900 -86.240 -273.870 ;
        RECT -88.670 -273.905 -86.240 -273.900 ;
        RECT -89.800 -274.095 -86.240 -273.905 ;
        RECT -84.455 -274.010 -84.150 -271.975 ;
        RECT -80.785 -272.255 -80.615 -270.785 ;
        RECT -80.295 -272.175 -80.125 -270.715 ;
        RECT -79.840 -270.790 -79.605 -270.195 ;
        RECT -81.330 -272.485 -80.555 -272.425 ;
        RECT -81.515 -272.655 -80.555 -272.485 ;
        RECT -81.330 -272.700 -80.555 -272.655 ;
        RECT -80.325 -272.525 -80.100 -272.175 ;
        RECT -79.805 -272.255 -79.635 -270.790 ;
        RECT -78.630 -270.840 -78.395 -270.195 ;
        RECT -78.595 -272.255 -78.425 -270.840 ;
        RECT -78.105 -272.210 -77.935 -270.715 ;
        RECT -69.285 -271.540 -69.045 -269.750 ;
        RECT -67.635 -269.835 -42.330 -269.640 ;
        RECT -39.180 -269.715 -38.985 -269.405 ;
        RECT -37.410 -269.715 -37.195 -268.495 ;
        RECT -36.310 -268.565 -36.140 -265.575 ;
        RECT -35.820 -268.465 -35.650 -265.525 ;
        RECT -35.350 -265.565 -35.140 -265.355 ;
        RECT -35.840 -268.735 -35.630 -268.465 ;
        RECT -35.330 -268.475 -35.160 -265.565 ;
        RECT -34.275 -268.445 -34.105 -265.525 ;
        RECT -30.220 -265.985 -26.580 -265.815 ;
        RECT -30.220 -267.545 -30.050 -265.985 ;
        RECT -29.730 -267.725 -29.560 -266.505 ;
        RECT -29.240 -267.545 -29.070 -265.985 ;
        RECT -28.640 -266.330 -26.930 -266.160 ;
        RECT -28.640 -267.545 -28.470 -266.330 ;
        RECT -28.150 -267.725 -27.980 -266.505 ;
        RECT -27.660 -267.545 -27.490 -266.330 ;
        RECT -30.775 -267.895 -27.405 -267.725 ;
        RECT -36.335 -268.930 -35.630 -268.735 ;
        RECT -35.355 -268.740 -35.145 -268.475 ;
        RECT -34.295 -268.740 -34.085 -268.445 ;
        RECT -35.355 -268.920 -34.085 -268.740 ;
        RECT -36.335 -268.990 -36.120 -268.930 ;
        RECT -37.025 -269.265 -36.120 -268.990 ;
        RECT -36.335 -269.615 -36.120 -269.265 ;
        RECT -35.685 -269.150 -34.910 -269.100 ;
        RECT -32.985 -269.150 -32.325 -268.795 ;
        RECT -35.685 -269.330 -32.325 -269.150 ;
        RECT -35.685 -269.375 -34.910 -269.330 ;
        RECT -65.605 -269.900 -64.945 -269.835 ;
        RECT -42.990 -269.890 -42.330 -269.835 ;
        RECT -39.200 -269.915 -36.525 -269.715 ;
        RECT -36.335 -269.815 -34.565 -269.615 ;
        RECT -39.200 -269.930 -36.765 -269.915 ;
        RECT -68.695 -270.410 -66.025 -270.070 ;
        RECT -64.040 -270.185 -60.875 -270.015 ;
        RECT -68.690 -271.125 -68.520 -270.665 ;
        RECT -68.720 -271.430 -68.490 -271.125 ;
        RECT -68.200 -271.205 -68.030 -270.410 ;
        RECT -67.710 -271.125 -67.540 -270.665 ;
        RECT -68.870 -271.540 -68.490 -271.430 ;
        RECT -69.285 -271.590 -68.490 -271.540 ;
        RECT -67.740 -271.590 -67.510 -271.125 ;
        RECT -67.220 -271.205 -67.050 -270.410 ;
        RECT -66.730 -271.125 -66.560 -270.665 ;
        RECT -66.760 -271.590 -66.530 -271.125 ;
        RECT -66.240 -271.205 -66.070 -270.410 ;
        RECT -64.500 -270.885 -64.330 -270.415 ;
        RECT -64.040 -270.475 -63.820 -270.185 ;
        RECT -64.520 -271.100 -64.315 -270.885 ;
        RECT -64.010 -270.955 -63.840 -270.475 ;
        RECT -63.520 -270.890 -63.350 -270.415 ;
        RECT -63.055 -270.530 -62.835 -270.185 ;
        RECT -64.525 -271.135 -64.315 -271.100 ;
        RECT -63.535 -271.135 -63.330 -270.890 ;
        RECT -63.030 -270.955 -62.860 -270.530 ;
        RECT -62.540 -270.890 -62.370 -270.415 ;
        RECT -62.075 -270.530 -61.855 -270.185 ;
        RECT -62.565 -271.135 -62.360 -270.890 ;
        RECT -62.050 -270.955 -61.880 -270.530 ;
        RECT -61.560 -270.930 -61.390 -270.415 ;
        RECT -61.095 -270.475 -60.875 -270.185 ;
        RECT -59.980 -270.410 -52.525 -270.070 ;
        RECT -50.540 -270.185 -47.375 -270.015 ;
        RECT -61.070 -270.825 -60.900 -270.475 ;
        RECT -61.575 -271.135 -61.370 -270.930 ;
        RECT -64.525 -271.305 -61.370 -271.135 ;
        RECT -69.285 -271.725 -66.530 -271.590 ;
        RECT -69.280 -271.735 -66.530 -271.725 ;
        RECT -68.870 -271.780 -66.530 -271.735 ;
        RECT -66.350 -271.450 -65.510 -271.375 ;
        RECT -64.525 -271.450 -63.650 -271.305 ;
        RECT -66.350 -271.715 -63.650 -271.450 ;
        RECT -61.105 -271.500 -60.870 -270.825 ;
        RECT -59.975 -271.125 -59.805 -270.665 ;
        RECT -60.005 -271.430 -59.775 -271.125 ;
        RECT -59.485 -271.205 -59.315 -270.410 ;
        RECT -58.995 -271.125 -58.825 -270.665 ;
        RECT -66.350 -271.745 -65.510 -271.715 ;
        RECT -68.720 -271.820 -66.530 -271.780 ;
        RECT -68.720 -272.145 -68.490 -271.820 ;
        RECT -67.740 -272.145 -67.510 -271.820 ;
        RECT -78.125 -272.410 -77.905 -272.210 ;
        RECT -78.125 -272.425 -72.425 -272.410 ;
        RECT -80.325 -272.725 -78.555 -272.525 ;
        RECT -78.365 -272.625 -72.425 -272.425 ;
        RECT -82.005 -273.010 -81.655 -273.000 ;
        RECT -79.980 -273.010 -79.205 -272.965 ;
        RECT -82.005 -273.190 -79.205 -273.010 ;
        RECT -89.800 -274.105 -88.665 -274.095 ;
        RECT -86.610 -274.225 -86.240 -274.095 ;
        RECT -94.580 -274.485 -92.330 -274.415 ;
        RECT -85.675 -274.440 -82.600 -274.010 ;
        RECT -101.960 -274.930 -92.180 -274.485 ;
        RECT -141.180 -275.470 -140.720 -275.050 ;
        RECT -143.220 -275.640 -140.720 -275.470 ;
        RECT -147.240 -280.465 -145.890 -275.945 ;
        RECT -144.245 -279.010 -143.645 -275.945 ;
        RECT -141.180 -276.060 -140.720 -275.640 ;
        RECT -143.220 -276.230 -140.720 -276.060 ;
        RECT -141.180 -276.650 -140.720 -276.230 ;
        RECT -109.855 -276.050 -109.550 -275.160 ;
        RECT -106.685 -275.245 -92.180 -274.930 ;
        RECT -88.020 -274.500 -85.925 -274.460 ;
        RECT -88.020 -274.650 -85.870 -274.500 ;
        RECT -106.685 -275.255 -100.315 -275.245 ;
        RECT -98.415 -276.050 -98.150 -275.570 ;
        RECT -109.855 -276.230 -98.150 -276.050 ;
        RECT -109.855 -276.240 -109.550 -276.230 ;
        RECT -88.020 -276.370 -87.850 -274.650 ;
        RECT -87.040 -276.370 -86.870 -274.650 ;
        RECT -86.175 -275.395 -85.870 -274.650 ;
        RECT -84.975 -275.220 -84.805 -274.440 ;
        RECT -84.485 -275.220 -84.315 -274.680 ;
        RECT -83.995 -275.220 -83.825 -274.440 ;
        RECT -83.505 -275.220 -83.335 -274.680 ;
        RECT -82.005 -275.165 -81.655 -273.190 ;
        RECT -79.980 -273.240 -79.205 -273.190 ;
        RECT -78.770 -273.075 -78.555 -272.725 ;
        RECT -78.770 -273.350 -77.865 -273.075 ;
        RECT -78.770 -273.410 -78.555 -273.350 ;
        RECT -80.805 -273.600 -79.535 -273.420 ;
        RECT -80.805 -273.895 -80.595 -273.600 ;
        RECT -79.745 -273.865 -79.535 -273.600 ;
        RECT -79.260 -273.605 -78.555 -273.410 ;
        RECT -85.565 -275.395 -85.200 -275.365 ;
        RECT -86.175 -275.460 -85.200 -275.395 ;
        RECT -86.065 -275.600 -85.200 -275.460 ;
        RECT -85.565 -275.665 -85.200 -275.600 ;
        RECT -83.015 -275.515 -81.625 -275.165 ;
        RECT -84.975 -276.375 -84.805 -275.835 ;
        RECT -83.995 -276.375 -83.825 -275.835 ;
        RECT -83.015 -276.375 -82.845 -275.515 ;
        RECT -143.220 -276.820 -140.720 -276.650 ;
        RECT -80.785 -276.815 -80.615 -273.895 ;
        RECT -79.730 -276.775 -79.560 -273.865 ;
        RECT -79.260 -273.875 -79.050 -273.605 ;
        RECT -141.180 -277.240 -140.720 -276.820 ;
        RECT -79.750 -276.985 -79.540 -276.775 ;
        RECT -79.240 -276.815 -79.070 -273.875 ;
        RECT -78.750 -276.765 -78.580 -273.775 ;
        RECT -77.695 -273.845 -77.480 -272.625 ;
        RECT -76.565 -273.500 -76.040 -273.140 ;
        RECT -78.760 -276.985 -78.550 -276.765 ;
        RECT -77.690 -276.815 -77.520 -273.845 ;
        RECT -79.750 -277.155 -78.550 -276.985 ;
        RECT -143.220 -277.410 -140.720 -277.240 ;
        RECT -141.180 -277.830 -140.720 -277.410 ;
        RECT -143.220 -278.000 -140.720 -277.830 ;
        RECT -141.180 -278.420 -140.720 -278.000 ;
        RECT -143.220 -278.590 -140.720 -278.420 ;
        RECT -141.180 -279.010 -140.860 -278.590 ;
        RECT -144.245 -279.180 -140.860 -279.010 ;
        RECT -144.245 -280.190 -143.645 -279.180 ;
        RECT -141.180 -279.330 -140.860 -279.180 ;
        RECT -140.690 -279.570 -139.910 -279.210 ;
        RECT -144.245 -280.360 -141.180 -280.190 ;
        RECT -144.245 -280.465 -143.645 -280.360 ;
        RECT -147.240 -281.370 -143.645 -280.465 ;
        RECT -140.350 -280.940 -140.180 -279.570 ;
        RECT -140.350 -281.110 -137.140 -280.940 ;
        RECT -108.560 -281.360 -108.260 -280.365 ;
        RECT -105.910 -281.285 -105.740 -279.565 ;
        RECT -104.930 -281.285 -104.760 -279.565 ;
        RECT -102.865 -280.100 -102.695 -279.560 ;
        RECT -101.885 -280.100 -101.715 -279.560 ;
        RECT -103.455 -280.335 -103.090 -280.270 ;
        RECT -103.955 -280.475 -103.090 -280.335 ;
        RECT -104.065 -280.540 -103.090 -280.475 ;
        RECT -104.065 -281.285 -103.760 -280.540 ;
        RECT -103.455 -280.570 -103.090 -280.540 ;
        RECT -100.905 -280.420 -100.735 -279.560 ;
        RECT -97.045 -280.310 -96.875 -279.090 ;
        RECT -96.065 -280.310 -95.895 -279.090 ;
        RECT -95.085 -280.310 -94.915 -279.090 ;
        RECT -97.920 -280.365 -97.245 -280.325 ;
        RECT -99.720 -280.420 -97.245 -280.365 ;
        RECT -100.905 -280.540 -97.245 -280.420 ;
        RECT -97.045 -280.495 -94.270 -280.310 ;
        RECT -106.825 -281.350 -106.150 -281.320 ;
        RECT -106.925 -281.360 -106.150 -281.350 ;
        RECT -147.240 -281.540 -141.180 -281.370 ;
        RECT -108.560 -281.540 -106.150 -281.360 ;
        RECT -105.910 -281.435 -103.760 -281.285 ;
        RECT -105.910 -281.475 -103.815 -281.435 ;
        RECT -102.865 -281.495 -102.695 -280.715 ;
        RECT -102.375 -281.255 -102.205 -280.715 ;
        RECT -101.885 -281.495 -101.715 -280.715 ;
        RECT -101.395 -281.255 -101.225 -280.715 ;
        RECT -100.905 -280.770 -99.515 -280.540 ;
        RECT -98.015 -280.550 -97.245 -280.540 ;
        RECT -97.920 -280.595 -97.245 -280.550 ;
        RECT -98.495 -280.780 -98.205 -280.740 ;
        RECT -96.240 -280.780 -95.565 -280.735 ;
        RECT -98.625 -280.970 -95.565 -280.780 ;
        RECT -147.240 -281.855 -143.645 -281.540 ;
        RECT -108.560 -281.550 -108.260 -281.540 ;
        RECT -106.925 -281.550 -106.150 -281.540 ;
        RECT -106.825 -281.590 -106.150 -281.550 ;
        RECT -147.240 -285.840 -145.890 -281.855 ;
        RECT -144.245 -282.550 -143.645 -281.855 ;
        RECT -109.190 -281.840 -106.555 -281.830 ;
        RECT -104.500 -281.840 -104.130 -281.710 ;
        RECT -109.190 -282.030 -104.130 -281.840 ;
        RECT -103.565 -281.925 -100.490 -281.495 ;
        RECT -139.180 -282.290 -137.140 -282.120 ;
        RECT -144.245 -282.720 -141.180 -282.550 ;
        RECT -109.190 -282.555 -108.990 -282.030 ;
        RECT -106.560 -282.035 -104.130 -282.030 ;
        RECT -106.560 -282.040 -106.205 -282.035 ;
        RECT -104.500 -282.065 -104.130 -282.035 ;
        RECT -144.245 -283.730 -143.645 -282.720 ;
        RECT -139.180 -283.470 -137.140 -283.300 ;
        RECT -144.245 -283.900 -141.180 -283.730 ;
        RECT -109.275 -283.740 -108.975 -282.555 ;
        RECT -106.400 -283.790 -106.230 -282.250 ;
        RECT -105.910 -283.790 -105.740 -282.250 ;
        RECT -105.420 -283.790 -105.250 -282.250 ;
        RECT -104.930 -283.790 -104.760 -282.250 ;
        RECT -104.440 -283.790 -104.270 -282.250 ;
        RECT -144.245 -284.910 -143.645 -283.900 ;
        RECT -105.915 -284.050 -105.740 -283.790 ;
        RECT -102.345 -283.960 -102.040 -281.925 ;
        RECT -100.050 -282.565 -99.760 -281.880 ;
        RECT -98.980 -281.895 -98.690 -281.395 ;
        RECT -98.495 -281.425 -98.205 -280.970 ;
        RECT -96.240 -281.005 -95.565 -280.970 ;
        RECT -95.300 -281.190 -94.625 -281.125 ;
        RECT -98.005 -281.360 -94.625 -281.190 ;
        RECT -98.005 -281.895 -97.835 -281.360 ;
        RECT -95.300 -281.395 -94.625 -281.360 ;
        RECT -94.455 -281.185 -94.270 -280.495 ;
        RECT -92.245 -281.185 -91.570 -281.135 ;
        RECT -94.455 -281.370 -91.570 -281.185 ;
        RECT -94.455 -281.640 -94.270 -281.370 ;
        RECT -92.245 -281.405 -91.570 -281.370 ;
        RECT -91.395 -281.495 -91.225 -279.090 ;
        RECT -87.890 -281.015 -87.720 -279.975 ;
        RECT -86.910 -281.015 -86.740 -279.975 ;
        RECT -85.930 -281.015 -85.760 -279.975 ;
        RECT -83.025 -281.050 -82.855 -279.330 ;
        RECT -82.045 -281.050 -81.875 -279.330 ;
        RECT -79.980 -279.865 -79.810 -279.325 ;
        RECT -79.000 -279.865 -78.830 -279.325 ;
        RECT -80.570 -280.100 -80.205 -280.035 ;
        RECT -81.070 -280.240 -80.205 -280.100 ;
        RECT -81.180 -280.305 -80.205 -280.240 ;
        RECT -81.180 -281.050 -80.875 -280.305 ;
        RECT -80.570 -280.335 -80.205 -280.305 ;
        RECT -78.020 -280.185 -77.850 -279.325 ;
        RECT -76.510 -280.185 -76.160 -273.500 ;
        RECT -83.940 -281.115 -83.265 -281.085 ;
        RECT -84.040 -281.125 -83.265 -281.115 ;
        RECT -89.350 -281.250 -88.700 -281.165 ;
        RECT -88.480 -281.250 -88.115 -281.185 ;
        RECT -89.350 -281.455 -88.115 -281.250 ;
        RECT -85.075 -281.305 -83.265 -281.125 ;
        RECT -83.025 -281.200 -80.875 -281.050 ;
        RECT -83.025 -281.240 -80.930 -281.200 ;
        RECT -79.980 -281.260 -79.810 -280.480 ;
        RECT -79.490 -281.020 -79.320 -280.480 ;
        RECT -79.000 -281.260 -78.830 -280.480 ;
        RECT -78.510 -281.020 -78.340 -280.480 ;
        RECT -78.020 -280.535 -76.160 -280.185 ;
        RECT -84.040 -281.315 -83.265 -281.305 ;
        RECT -83.940 -281.355 -83.265 -281.315 ;
        RECT -89.350 -281.495 -88.700 -281.455 ;
        RECT -88.480 -281.485 -88.115 -281.455 ;
        RECT -98.980 -282.065 -97.835 -281.895 ;
        RECT -97.535 -281.810 -95.320 -281.640 ;
        RECT -94.455 -281.810 -93.290 -281.640 ;
        RECT -98.980 -282.080 -98.690 -282.065 ;
        RECT -97.535 -283.665 -97.365 -281.810 ;
        RECT -96.555 -281.815 -95.320 -281.810 ;
        RECT -104.290 -284.050 -98.445 -283.960 ;
        RECT -106.500 -284.355 -98.445 -284.050 ;
        RECT -139.180 -284.650 -137.140 -284.480 ;
        RECT -104.295 -284.535 -98.445 -284.355 ;
        RECT -99.020 -284.625 -98.445 -284.535 ;
        RECT -97.045 -284.610 -96.875 -282.125 ;
        RECT -96.555 -283.665 -96.385 -281.815 ;
        RECT -95.495 -282.130 -95.320 -281.815 ;
        RECT -95.985 -283.625 -95.815 -282.130 ;
        RECT -95.985 -284.145 -95.810 -283.625 ;
        RECT -95.495 -283.670 -95.325 -282.130 ;
        RECT -95.005 -283.615 -94.835 -282.130 ;
        RECT -95.005 -284.145 -94.830 -283.615 ;
        RECT -94.440 -283.670 -94.270 -281.810 ;
        RECT -95.985 -284.160 -94.830 -284.145 ;
        RECT -93.950 -284.160 -93.780 -282.130 ;
        RECT -93.460 -283.670 -93.290 -281.810 ;
        RECT -91.395 -281.665 -88.700 -281.495 ;
        RECT -86.415 -281.605 -83.670 -281.595 ;
        RECT -81.615 -281.605 -81.245 -281.475 ;
        RECT -86.415 -281.625 -81.245 -281.605 ;
        RECT -95.985 -284.330 -93.780 -284.160 ;
        RECT -91.885 -284.475 -91.715 -282.630 ;
        RECT -91.395 -283.670 -91.225 -281.665 ;
        RECT -89.350 -281.915 -88.700 -281.665 ;
        RECT -87.890 -282.905 -87.720 -281.625 ;
        RECT -87.400 -282.665 -87.230 -281.625 ;
        RECT -86.910 -282.905 -86.740 -281.625 ;
        RECT -86.420 -281.795 -81.245 -281.625 ;
        RECT -80.680 -281.690 -76.755 -281.260 ;
        RECT -86.420 -282.665 -86.250 -281.795 ;
        RECT -83.675 -281.800 -81.245 -281.795 ;
        RECT -83.675 -281.805 -83.320 -281.800 ;
        RECT -81.615 -281.830 -81.245 -281.800 ;
        RECT -88.590 -283.335 -83.900 -282.905 ;
        RECT -84.330 -283.740 -83.900 -283.335 ;
        RECT -83.515 -283.555 -83.345 -282.015 ;
        RECT -83.025 -283.555 -82.855 -282.015 ;
        RECT -82.535 -283.555 -82.365 -282.015 ;
        RECT -82.045 -283.555 -81.875 -282.015 ;
        RECT -81.555 -283.555 -81.385 -282.015 ;
        RECT -83.030 -283.740 -82.855 -283.555 ;
        RECT -79.460 -283.725 -79.155 -281.690 ;
        RECT -81.405 -283.740 -79.155 -283.725 ;
        RECT -84.330 -284.030 -79.155 -283.740 ;
        RECT -84.330 -284.170 -81.005 -284.030 ;
        RECT -84.150 -284.475 -83.100 -284.170 ;
        RECT -92.890 -284.610 -83.100 -284.475 ;
        RECT -97.535 -284.625 -83.100 -284.610 ;
        RECT -144.245 -285.080 -141.180 -284.910 ;
        RECT -144.245 -285.840 -143.645 -285.080 ;
        RECT -99.020 -285.250 -83.100 -284.625 ;
        RECT -78.490 -284.420 -77.150 -284.170 ;
        RECT -73.340 -284.420 -72.425 -272.625 ;
        RECT -68.690 -273.105 -68.520 -272.145 ;
        RECT -67.710 -273.105 -67.540 -272.145 ;
        RECT -66.760 -273.085 -66.530 -271.820 ;
        RECT -64.525 -272.140 -63.650 -271.715 ;
        RECT -61.730 -271.870 -60.870 -271.500 ;
        RECT -64.525 -272.310 -61.385 -272.140 ;
        RECT -64.525 -272.530 -64.315 -272.310 ;
        RECT -64.500 -273.030 -64.330 -272.530 ;
        RECT -64.010 -272.945 -63.840 -272.490 ;
        RECT -63.525 -272.580 -63.345 -272.310 ;
        RECT -62.555 -272.490 -62.375 -272.310 ;
        RECT -66.730 -273.105 -66.560 -273.085 ;
        RECT -64.035 -273.200 -63.825 -272.945 ;
        RECT -63.520 -273.030 -63.350 -272.580 ;
        RECT -63.030 -272.920 -62.860 -272.490 ;
        RECT -62.555 -272.580 -62.370 -272.490 ;
        RECT -63.055 -273.200 -62.845 -272.920 ;
        RECT -62.540 -273.030 -62.370 -272.580 ;
        RECT -62.050 -272.925 -61.880 -272.490 ;
        RECT -61.565 -272.570 -61.385 -272.310 ;
        RECT -62.085 -273.200 -61.875 -272.925 ;
        RECT -61.560 -273.030 -61.390 -272.570 ;
        RECT -61.105 -272.605 -60.870 -271.870 ;
        RECT -60.645 -271.590 -59.775 -271.430 ;
        RECT -59.025 -271.590 -58.795 -271.125 ;
        RECT -58.505 -271.205 -58.335 -270.410 ;
        RECT -58.015 -271.125 -57.845 -270.665 ;
        RECT -58.045 -271.590 -57.815 -271.125 ;
        RECT -57.525 -271.205 -57.355 -270.410 ;
        RECT -60.645 -271.780 -57.815 -271.590 ;
        RECT -57.635 -271.400 -56.795 -271.375 ;
        RECT -56.495 -271.400 -56.195 -271.035 ;
        RECT -57.635 -271.690 -56.195 -271.400 ;
        RECT -55.920 -271.485 -55.620 -270.910 ;
        RECT -55.190 -271.125 -55.020 -270.665 ;
        RECT -55.220 -271.430 -54.990 -271.125 ;
        RECT -54.700 -271.205 -54.530 -270.410 ;
        RECT -54.210 -271.125 -54.040 -270.665 ;
        RECT -55.370 -271.485 -54.990 -271.430 ;
        RECT -57.635 -271.745 -56.795 -271.690 ;
        RECT -56.495 -271.695 -56.195 -271.690 ;
        RECT -55.945 -271.590 -54.990 -271.485 ;
        RECT -54.240 -271.590 -54.010 -271.125 ;
        RECT -53.720 -271.205 -53.550 -270.410 ;
        RECT -53.230 -271.125 -53.060 -270.665 ;
        RECT -53.260 -271.590 -53.030 -271.125 ;
        RECT -52.740 -271.205 -52.570 -270.410 ;
        RECT -51.015 -270.885 -50.785 -270.275 ;
        RECT -50.540 -270.475 -50.320 -270.185 ;
        RECT -51.020 -270.935 -50.785 -270.885 ;
        RECT -51.020 -271.100 -50.815 -270.935 ;
        RECT -50.510 -270.955 -50.340 -270.475 ;
        RECT -50.020 -270.890 -49.850 -270.415 ;
        RECT -49.555 -270.530 -49.335 -270.185 ;
        RECT -51.025 -271.135 -50.815 -271.100 ;
        RECT -50.035 -271.135 -49.830 -270.890 ;
        RECT -49.530 -270.955 -49.360 -270.530 ;
        RECT -49.040 -270.890 -48.870 -270.415 ;
        RECT -48.575 -270.530 -48.355 -270.185 ;
        RECT -49.065 -271.135 -48.860 -270.890 ;
        RECT -48.550 -270.955 -48.380 -270.530 ;
        RECT -48.060 -270.930 -47.890 -270.415 ;
        RECT -47.595 -270.475 -47.375 -270.185 ;
        RECT -46.480 -270.410 -39.400 -270.070 ;
        RECT -47.570 -270.825 -47.400 -270.475 ;
        RECT -48.075 -271.135 -47.870 -270.930 ;
        RECT -51.025 -271.305 -47.870 -271.135 ;
        RECT -55.945 -271.710 -53.030 -271.590 ;
        RECT -60.645 -271.900 -60.280 -271.780 ;
        RECT -61.070 -272.975 -60.900 -272.605 ;
        RECT -60.650 -272.740 -60.280 -271.900 ;
        RECT -60.005 -271.820 -57.815 -271.780 ;
        RECT -60.005 -272.145 -59.775 -271.820 ;
        RECT -59.025 -272.145 -58.795 -271.820 ;
        RECT -61.075 -273.200 -60.895 -272.975 ;
        RECT -59.975 -273.105 -59.805 -272.145 ;
        RECT -58.995 -273.105 -58.825 -272.145 ;
        RECT -58.045 -273.085 -57.815 -271.820 ;
        RECT -57.025 -272.380 -56.740 -272.175 ;
        RECT -55.945 -272.380 -55.720 -271.710 ;
        RECT -55.370 -271.780 -53.030 -271.710 ;
        RECT -52.850 -271.415 -52.010 -271.375 ;
        RECT -51.025 -271.415 -50.150 -271.305 ;
        RECT -52.850 -271.700 -50.150 -271.415 ;
        RECT -47.605 -271.500 -47.370 -270.825 ;
        RECT -46.475 -271.125 -46.305 -270.665 ;
        RECT -46.505 -271.430 -46.275 -271.125 ;
        RECT -45.985 -271.205 -45.815 -270.410 ;
        RECT -45.495 -271.125 -45.325 -270.665 ;
        RECT -52.850 -271.745 -52.010 -271.700 ;
        RECT -55.220 -271.820 -53.030 -271.780 ;
        RECT -55.220 -272.145 -54.990 -271.820 ;
        RECT -54.240 -272.145 -54.010 -271.820 ;
        RECT -57.025 -272.605 -55.720 -272.380 ;
        RECT -57.025 -272.995 -56.740 -272.605 ;
        RECT -58.015 -273.105 -57.845 -273.085 ;
        RECT -55.190 -273.105 -55.020 -272.145 ;
        RECT -54.210 -273.105 -54.040 -272.145 ;
        RECT -53.260 -273.085 -53.030 -271.820 ;
        RECT -51.025 -272.140 -50.150 -271.700 ;
        RECT -48.230 -271.870 -47.370 -271.500 ;
        RECT -51.025 -272.310 -47.885 -272.140 ;
        RECT -51.025 -272.530 -50.815 -272.310 ;
        RECT -51.000 -273.030 -50.830 -272.530 ;
        RECT -50.510 -272.945 -50.340 -272.490 ;
        RECT -50.025 -272.580 -49.845 -272.310 ;
        RECT -49.055 -272.490 -48.875 -272.310 ;
        RECT -53.230 -273.105 -53.060 -273.085 ;
        RECT -64.035 -273.370 -60.895 -273.200 ;
        RECT -50.535 -273.200 -50.325 -272.945 ;
        RECT -50.020 -273.030 -49.850 -272.580 ;
        RECT -49.530 -272.920 -49.360 -272.490 ;
        RECT -49.055 -272.580 -48.870 -272.490 ;
        RECT -49.555 -273.200 -49.345 -272.920 ;
        RECT -49.040 -273.030 -48.870 -272.580 ;
        RECT -48.550 -272.925 -48.380 -272.490 ;
        RECT -48.065 -272.570 -47.885 -272.310 ;
        RECT -48.585 -273.200 -48.375 -272.925 ;
        RECT -48.060 -273.030 -47.890 -272.570 ;
        RECT -47.605 -272.605 -47.370 -271.870 ;
        RECT -47.145 -271.590 -46.275 -271.430 ;
        RECT -45.525 -271.590 -45.295 -271.125 ;
        RECT -45.005 -271.205 -44.835 -270.410 ;
        RECT -44.515 -271.125 -44.345 -270.665 ;
        RECT -44.545 -271.590 -44.315 -271.125 ;
        RECT -44.025 -271.205 -43.855 -270.410 ;
        RECT -47.145 -271.780 -44.315 -271.590 ;
        RECT -44.135 -271.400 -43.295 -271.375 ;
        RECT -44.135 -271.460 -43.120 -271.400 ;
        RECT -42.835 -271.460 -42.535 -271.030 ;
        RECT -42.065 -271.125 -41.895 -270.665 ;
        RECT -42.095 -271.430 -41.865 -271.125 ;
        RECT -41.575 -271.205 -41.405 -270.410 ;
        RECT -41.085 -271.125 -40.915 -270.665 ;
        RECT -42.245 -271.460 -41.865 -271.430 ;
        RECT -44.135 -271.590 -41.865 -271.460 ;
        RECT -41.115 -271.590 -40.885 -271.125 ;
        RECT -40.595 -271.205 -40.425 -270.410 ;
        RECT -40.105 -271.125 -39.935 -270.665 ;
        RECT -40.135 -271.590 -39.905 -271.125 ;
        RECT -39.615 -271.205 -39.445 -270.410 ;
        RECT -39.180 -271.375 -38.985 -269.930 ;
        RECT -36.985 -270.130 -36.765 -269.930 ;
        RECT -44.135 -271.670 -39.905 -271.590 ;
        RECT -44.135 -271.690 -43.120 -271.670 ;
        RECT -42.835 -271.690 -42.535 -271.670 ;
        RECT -44.135 -271.745 -43.295 -271.690 ;
        RECT -42.245 -271.780 -39.905 -271.670 ;
        RECT -39.725 -271.745 -38.885 -271.375 ;
        RECT -36.955 -271.625 -36.785 -270.130 ;
        RECT -36.465 -271.500 -36.295 -270.085 ;
        RECT -47.145 -271.900 -46.780 -271.780 ;
        RECT -47.570 -272.975 -47.400 -272.605 ;
        RECT -47.150 -272.740 -46.780 -271.900 ;
        RECT -46.505 -271.820 -44.315 -271.780 ;
        RECT -46.505 -272.145 -46.275 -271.820 ;
        RECT -45.525 -272.145 -45.295 -271.820 ;
        RECT -47.575 -273.200 -47.395 -272.975 ;
        RECT -46.475 -273.105 -46.305 -272.145 ;
        RECT -45.495 -273.105 -45.325 -272.145 ;
        RECT -44.545 -273.085 -44.315 -271.820 ;
        RECT -42.095 -271.820 -39.905 -271.780 ;
        RECT -42.095 -272.145 -41.865 -271.820 ;
        RECT -41.115 -272.145 -40.885 -271.820 ;
        RECT -43.525 -272.995 -43.240 -272.175 ;
        RECT -44.515 -273.105 -44.345 -273.085 ;
        RECT -42.065 -273.105 -41.895 -272.145 ;
        RECT -41.085 -273.105 -40.915 -272.145 ;
        RECT -40.135 -273.085 -39.905 -271.820 ;
        RECT -38.615 -272.150 -37.225 -272.145 ;
        RECT -36.495 -272.150 -36.260 -271.500 ;
        RECT -35.255 -271.550 -35.085 -270.085 ;
        RECT -34.790 -270.165 -34.565 -269.815 ;
        RECT -34.335 -269.685 -33.560 -269.640 ;
        RECT -34.335 -269.855 -31.525 -269.685 ;
        RECT -34.335 -269.915 -33.560 -269.855 ;
        RECT -35.285 -272.150 -35.050 -271.550 ;
        RECT -34.765 -271.625 -34.595 -270.165 ;
        RECT -34.275 -271.555 -34.105 -270.085 ;
        RECT -34.305 -272.150 -34.070 -271.555 ;
        RECT -38.615 -272.560 -33.660 -272.150 ;
        RECT -40.105 -273.105 -39.935 -273.085 ;
        RECT -50.535 -273.370 -47.395 -273.200 ;
        RECT -59.510 -275.075 -52.125 -274.510 ;
        RECT -63.665 -276.550 -61.420 -276.460 ;
        RECT -59.510 -276.550 -59.205 -275.075 ;
        RECT -55.875 -275.665 -55.640 -275.075 ;
        RECT -63.665 -276.765 -59.205 -276.550 ;
        RECT -63.080 -277.025 -62.905 -276.765 ;
        RECT -61.455 -276.855 -59.205 -276.765 ;
        RECT -63.565 -278.565 -63.395 -277.025 ;
        RECT -63.075 -278.565 -62.905 -277.025 ;
        RECT -62.585 -278.565 -62.415 -277.025 ;
        RECT -62.095 -278.565 -61.925 -277.025 ;
        RECT -61.605 -278.565 -61.435 -277.025 ;
        RECT -59.510 -278.890 -59.205 -276.855 ;
        RECT -55.840 -277.135 -55.670 -275.665 ;
        RECT -55.350 -277.055 -55.180 -275.595 ;
        RECT -54.895 -275.670 -54.660 -275.075 ;
        RECT -56.385 -277.365 -55.610 -277.305 ;
        RECT -56.570 -277.535 -55.610 -277.365 ;
        RECT -56.385 -277.580 -55.610 -277.535 ;
        RECT -55.380 -277.405 -55.155 -277.055 ;
        RECT -54.860 -277.135 -54.690 -275.670 ;
        RECT -53.685 -275.720 -53.450 -275.075 ;
        RECT -53.650 -277.135 -53.480 -275.720 ;
        RECT -53.160 -277.090 -52.990 -275.595 ;
        RECT -53.180 -277.290 -52.960 -277.090 ;
        RECT -53.180 -277.305 -37.780 -277.290 ;
        RECT -55.380 -277.605 -53.610 -277.405 ;
        RECT -53.420 -277.505 -37.780 -277.305 ;
        RECT -57.060 -277.890 -56.710 -277.880 ;
        RECT -55.035 -277.890 -54.260 -277.845 ;
        RECT -57.060 -278.070 -54.260 -277.890 ;
        RECT -66.290 -279.275 -65.360 -278.990 ;
        RECT -63.990 -279.265 -63.315 -279.225 ;
        RECT -64.090 -279.275 -63.315 -279.265 ;
        RECT -66.290 -279.455 -63.315 -279.275 ;
        RECT -60.730 -279.320 -57.655 -278.890 ;
        RECT -66.290 -279.760 -65.360 -279.455 ;
        RECT -64.090 -279.465 -63.315 -279.455 ;
        RECT -63.990 -279.495 -63.315 -279.465 ;
        RECT -63.075 -279.380 -60.980 -279.340 ;
        RECT -63.075 -279.530 -60.925 -279.380 ;
        RECT -63.075 -281.250 -62.905 -279.530 ;
        RECT -62.095 -281.250 -61.925 -279.530 ;
        RECT -61.230 -280.275 -60.925 -279.530 ;
        RECT -60.030 -280.100 -59.860 -279.320 ;
        RECT -59.540 -280.100 -59.370 -279.560 ;
        RECT -59.050 -280.100 -58.880 -279.320 ;
        RECT -58.560 -280.100 -58.390 -279.560 ;
        RECT -57.060 -280.045 -56.710 -278.070 ;
        RECT -55.035 -278.120 -54.260 -278.070 ;
        RECT -53.825 -277.955 -53.610 -277.605 ;
        RECT -53.825 -278.230 -52.920 -277.955 ;
        RECT -53.825 -278.290 -53.610 -278.230 ;
        RECT -55.860 -278.480 -54.590 -278.300 ;
        RECT -55.860 -278.775 -55.650 -278.480 ;
        RECT -54.800 -278.745 -54.590 -278.480 ;
        RECT -54.315 -278.485 -53.610 -278.290 ;
        RECT -60.620 -280.275 -60.255 -280.245 ;
        RECT -61.230 -280.340 -60.255 -280.275 ;
        RECT -61.120 -280.480 -60.255 -280.340 ;
        RECT -60.620 -280.545 -60.255 -280.480 ;
        RECT -58.070 -280.395 -56.680 -280.045 ;
        RECT -60.030 -281.255 -59.860 -280.715 ;
        RECT -59.050 -281.255 -58.880 -280.715 ;
        RECT -58.070 -281.255 -57.900 -280.395 ;
        RECT -55.840 -281.695 -55.670 -278.775 ;
        RECT -54.785 -281.655 -54.615 -278.745 ;
        RECT -54.315 -278.755 -54.105 -278.485 ;
        RECT -54.805 -281.865 -54.595 -281.655 ;
        RECT -54.295 -281.695 -54.125 -278.755 ;
        RECT -53.805 -281.645 -53.635 -278.655 ;
        RECT -52.750 -278.725 -52.535 -277.505 ;
        RECT -38.660 -277.900 -37.780 -277.505 ;
        RECT -51.620 -278.380 -51.095 -278.020 ;
        RECT -53.815 -281.865 -53.605 -281.645 ;
        RECT -52.745 -281.695 -52.575 -278.725 ;
        RECT -54.805 -282.035 -53.605 -281.865 ;
        RECT -99.020 -285.280 -98.445 -285.250 ;
        RECT -139.180 -285.830 -137.140 -285.660 ;
        RECT -147.240 -286.090 -143.645 -285.840 ;
        RECT -132.635 -285.855 -98.445 -285.280 ;
        RECT -78.490 -285.335 -72.425 -284.420 ;
        RECT -78.490 -285.495 -77.150 -285.335 ;
        RECT -147.240 -286.260 -141.180 -286.090 ;
        RECT -147.240 -287.230 -143.645 -286.260 ;
        RECT -139.180 -287.010 -137.140 -286.840 ;
        RECT -147.240 -291.645 -145.890 -287.230 ;
        RECT -144.245 -287.270 -143.645 -287.230 ;
        RECT -144.245 -287.440 -141.180 -287.270 ;
        RECT -144.245 -288.450 -143.645 -287.440 ;
        RECT -139.180 -288.190 -137.140 -288.020 ;
        RECT -144.245 -288.620 -141.180 -288.450 ;
        RECT -144.245 -289.630 -143.645 -288.620 ;
        RECT -140.520 -289.010 -139.740 -288.650 ;
        RECT -143.220 -289.210 -141.180 -289.040 ;
        RECT -144.245 -289.800 -141.180 -289.630 ;
        RECT -144.245 -290.810 -143.645 -289.800 ;
        RECT -143.220 -290.390 -141.180 -290.220 ;
        RECT -144.245 -290.980 -141.180 -290.810 ;
        RECT -144.245 -291.645 -143.645 -290.980 ;
        RECT -140.280 -291.030 -140.110 -289.010 ;
        RECT -139.180 -289.370 -137.140 -289.200 ;
        RECT -140.280 -291.200 -137.140 -291.030 ;
        RECT -143.220 -291.570 -141.180 -291.400 ;
        RECT -147.240 -291.990 -143.645 -291.645 ;
        RECT -147.240 -292.160 -141.180 -291.990 ;
        RECT -147.240 -293.035 -143.645 -292.160 ;
        RECT -139.180 -292.380 -137.140 -292.210 ;
        RECT -143.220 -292.750 -141.180 -292.580 ;
        RECT -147.240 -295.815 -145.890 -293.035 ;
        RECT -144.245 -293.170 -143.645 -293.035 ;
        RECT -144.245 -293.340 -141.180 -293.170 ;
        RECT -144.245 -294.350 -143.645 -293.340 ;
        RECT -143.220 -293.930 -141.180 -293.760 ;
        RECT -140.585 -293.815 -139.885 -293.305 ;
        RECT -139.180 -293.560 -137.140 -293.390 ;
        RECT -144.245 -294.520 -141.180 -294.350 ;
        RECT -144.245 -295.530 -143.645 -294.520 ;
        RECT -143.220 -295.110 -141.180 -294.940 ;
        RECT -140.295 -295.530 -140.125 -293.815 ;
        RECT -139.180 -294.740 -137.140 -294.570 ;
        RECT -144.245 -295.700 -141.180 -295.530 ;
        RECT -140.295 -295.700 -139.510 -295.530 ;
        RECT -144.245 -296.710 -143.645 -295.700 ;
        RECT -143.220 -296.290 -141.180 -296.120 ;
        RECT -140.860 -296.695 -139.975 -296.315 ;
        RECT -139.680 -296.400 -139.510 -295.700 ;
        RECT -139.680 -296.570 -137.140 -296.400 ;
        RECT -144.245 -296.880 -141.180 -296.710 ;
        RECT -144.245 -297.090 -143.645 -296.880 ;
        RECT -140.580 -299.075 -140.275 -296.695 ;
        RECT -139.180 -297.750 -137.140 -297.580 ;
        RECT -140.735 -311.555 -140.050 -299.075 ;
        RECT -136.180 -303.680 -134.480 -302.835 ;
        RECT -132.635 -303.680 -132.060 -285.855 ;
        RECT -62.945 -285.895 -62.775 -284.855 ;
        RECT -61.965 -285.895 -61.795 -284.855 ;
        RECT -60.985 -285.895 -60.815 -284.855 ;
        RECT -58.080 -285.930 -57.910 -284.210 ;
        RECT -57.100 -285.930 -56.930 -284.210 ;
        RECT -55.035 -284.745 -54.865 -284.205 ;
        RECT -54.055 -284.745 -53.885 -284.205 ;
        RECT -55.625 -284.980 -55.260 -284.915 ;
        RECT -56.125 -285.120 -55.260 -284.980 ;
        RECT -56.235 -285.185 -55.260 -285.120 ;
        RECT -56.235 -285.930 -55.930 -285.185 ;
        RECT -55.625 -285.215 -55.260 -285.185 ;
        RECT -53.075 -285.065 -52.905 -284.205 ;
        RECT -51.565 -285.065 -51.215 -278.380 ;
        RECT -31.695 -281.150 -31.525 -269.855 ;
        RECT -30.775 -275.595 -30.605 -267.895 ;
        RECT -30.225 -268.565 -29.530 -268.295 ;
        RECT -27.575 -268.470 -27.405 -267.895 ;
        RECT -27.100 -268.090 -26.930 -266.330 ;
        RECT -26.750 -267.720 -26.580 -265.985 ;
        RECT -17.720 -265.985 -14.080 -265.815 ;
        RECT -25.850 -267.720 -25.680 -266.505 ;
        RECT -26.750 -267.890 -25.680 -267.720 ;
        RECT -24.870 -268.090 -24.700 -266.505 ;
        RECT -23.320 -267.470 -23.150 -266.505 ;
        RECT -21.775 -267.460 -21.605 -266.505 ;
        RECT -27.100 -268.260 -24.700 -268.090 ;
        RECT -24.435 -268.345 -23.740 -268.075 ;
        RECT -27.575 -268.640 -26.845 -268.470 ;
        RECT -30.230 -269.155 -28.575 -268.970 ;
        RECT -28.315 -269.085 -27.620 -268.815 ;
        RECT -27.015 -268.950 -26.845 -268.640 ;
        RECT -26.480 -268.715 -25.785 -268.445 ;
        RECT -27.015 -269.120 -24.210 -268.950 ;
        RECT -30.230 -269.570 -30.045 -269.155 ;
        RECT -28.760 -269.275 -28.575 -269.155 ;
        RECT -28.760 -269.460 -27.980 -269.275 ;
        RECT -30.220 -270.515 -30.050 -269.570 ;
        RECT -30.240 -271.130 -30.045 -270.515 ;
        RECT -29.730 -270.760 -29.560 -269.535 ;
        RECT -28.165 -269.565 -27.980 -269.460 ;
        RECT -28.150 -270.575 -27.980 -269.565 ;
        RECT -27.670 -269.580 -26.170 -269.385 ;
        RECT -27.660 -270.575 -27.490 -269.580 ;
        RECT -26.340 -270.575 -26.170 -269.580 ;
        RECT -25.850 -270.575 -25.680 -269.120 ;
        RECT -24.870 -270.490 -24.700 -269.535 ;
        RECT -24.870 -270.760 -24.690 -270.490 ;
        RECT -24.380 -270.575 -24.210 -269.120 ;
        RECT -23.345 -269.165 -23.130 -267.470 ;
        RECT -21.795 -268.445 -21.580 -267.460 ;
        RECT -17.720 -267.545 -17.550 -265.985 ;
        RECT -17.230 -267.725 -17.060 -266.505 ;
        RECT -16.740 -267.545 -16.570 -265.985 ;
        RECT -16.140 -266.330 -14.430 -266.160 ;
        RECT -16.140 -267.545 -15.970 -266.330 ;
        RECT -15.650 -267.725 -15.480 -266.505 ;
        RECT -15.160 -267.545 -14.990 -266.330 ;
        RECT -18.560 -267.895 -14.905 -267.725 ;
        RECT -21.360 -268.375 -20.665 -268.105 ;
        RECT -22.295 -268.675 -21.580 -268.445 ;
        RECT -22.925 -269.115 -22.230 -268.845 ;
        RECT -23.825 -269.395 -23.130 -269.165 ;
        RECT -23.345 -269.620 -23.130 -269.395 ;
        RECT -23.320 -270.575 -23.150 -269.620 ;
        RECT -22.830 -270.540 -22.660 -269.535 ;
        RECT -21.795 -269.630 -21.580 -268.675 ;
        RECT -29.730 -270.940 -24.690 -270.760 ;
        RECT -22.855 -270.960 -22.640 -270.540 ;
        RECT -21.775 -270.575 -21.605 -269.630 ;
        RECT -21.285 -270.530 -21.115 -269.535 ;
        RECT -18.560 -269.710 -18.390 -267.895 ;
        RECT -17.725 -268.565 -17.030 -268.295 ;
        RECT -15.075 -268.470 -14.905 -267.895 ;
        RECT -14.600 -268.090 -14.430 -266.330 ;
        RECT -14.250 -267.720 -14.080 -265.985 ;
        RECT -5.220 -265.985 -1.580 -265.815 ;
        RECT -13.350 -267.720 -13.180 -266.505 ;
        RECT -14.250 -267.890 -13.180 -267.720 ;
        RECT -12.370 -268.090 -12.200 -266.505 ;
        RECT -10.820 -267.470 -10.650 -266.505 ;
        RECT -9.275 -267.460 -9.105 -266.505 ;
        RECT -14.600 -268.260 -12.200 -268.090 ;
        RECT -11.935 -268.345 -11.240 -268.075 ;
        RECT -15.075 -268.640 -14.345 -268.470 ;
        RECT -17.730 -269.155 -16.075 -268.970 ;
        RECT -15.815 -269.085 -15.120 -268.815 ;
        RECT -14.515 -268.950 -14.345 -268.640 ;
        RECT -13.980 -268.715 -13.285 -268.445 ;
        RECT -14.515 -269.120 -11.710 -268.950 ;
        RECT -17.730 -269.570 -17.545 -269.155 ;
        RECT -16.260 -269.275 -16.075 -269.155 ;
        RECT -16.260 -269.460 -15.480 -269.275 ;
        RECT -18.590 -270.390 -18.360 -269.710 ;
        RECT -17.720 -270.515 -17.550 -269.570 ;
        RECT -21.310 -270.955 -21.095 -270.530 ;
        RECT -17.740 -270.955 -17.545 -270.515 ;
        RECT -17.230 -270.760 -17.060 -269.535 ;
        RECT -15.665 -269.565 -15.480 -269.460 ;
        RECT -15.650 -270.575 -15.480 -269.565 ;
        RECT -15.170 -269.580 -13.670 -269.385 ;
        RECT -15.160 -270.575 -14.990 -269.580 ;
        RECT -13.840 -270.575 -13.670 -269.580 ;
        RECT -13.350 -270.575 -13.180 -269.120 ;
        RECT -12.370 -270.490 -12.200 -269.535 ;
        RECT -12.370 -270.760 -12.190 -270.490 ;
        RECT -11.880 -270.575 -11.710 -269.120 ;
        RECT -10.845 -269.165 -10.630 -267.470 ;
        RECT -9.295 -268.445 -9.080 -267.460 ;
        RECT -5.220 -267.545 -5.050 -265.985 ;
        RECT -4.730 -267.725 -4.560 -266.505 ;
        RECT -4.240 -267.545 -4.070 -265.985 ;
        RECT -3.640 -266.330 -1.930 -266.160 ;
        RECT -3.640 -267.545 -3.470 -266.330 ;
        RECT -3.150 -267.725 -2.980 -266.505 ;
        RECT -2.660 -267.545 -2.490 -266.330 ;
        RECT -5.820 -267.895 -2.405 -267.725 ;
        RECT -8.860 -268.375 -8.165 -268.105 ;
        RECT -9.795 -268.675 -9.080 -268.445 ;
        RECT -10.425 -269.115 -9.730 -268.845 ;
        RECT -11.325 -269.395 -10.630 -269.165 ;
        RECT -10.845 -269.620 -10.630 -269.395 ;
        RECT -10.820 -270.575 -10.650 -269.620 ;
        RECT -10.330 -270.540 -10.160 -269.535 ;
        RECT -9.295 -269.630 -9.080 -268.675 ;
        RECT -17.230 -270.940 -12.190 -270.760 ;
        RECT -21.680 -270.960 -17.545 -270.955 ;
        RECT -10.355 -270.960 -10.140 -270.540 ;
        RECT -9.275 -270.575 -9.105 -269.630 ;
        RECT -8.785 -270.530 -8.615 -269.535 ;
        RECT -5.820 -269.730 -5.650 -267.895 ;
        RECT -5.225 -268.565 -4.530 -268.295 ;
        RECT -2.575 -268.470 -2.405 -267.895 ;
        RECT -2.100 -268.090 -1.930 -266.330 ;
        RECT -1.750 -267.720 -1.580 -265.985 ;
        RECT 7.280 -265.985 10.920 -265.815 ;
        RECT -0.850 -267.720 -0.680 -266.505 ;
        RECT -1.750 -267.890 -0.680 -267.720 ;
        RECT 0.130 -268.090 0.300 -266.505 ;
        RECT 1.680 -267.470 1.850 -266.505 ;
        RECT 3.225 -267.460 3.395 -266.505 ;
        RECT -2.100 -268.260 0.300 -268.090 ;
        RECT 0.565 -268.345 1.260 -268.075 ;
        RECT -2.575 -268.640 -1.845 -268.470 ;
        RECT -5.230 -269.155 -3.575 -268.970 ;
        RECT -3.315 -269.085 -2.620 -268.815 ;
        RECT -2.015 -268.950 -1.845 -268.640 ;
        RECT -1.480 -268.715 -0.785 -268.445 ;
        RECT -2.015 -269.120 0.790 -268.950 ;
        RECT -5.230 -269.570 -5.045 -269.155 ;
        RECT -3.760 -269.275 -3.575 -269.155 ;
        RECT -3.760 -269.460 -2.980 -269.275 ;
        RECT -5.850 -270.410 -5.620 -269.730 ;
        RECT -5.220 -270.515 -5.050 -269.570 ;
        RECT -8.810 -270.960 -8.595 -270.530 ;
        RECT -24.235 -271.130 -17.545 -270.960 ;
        RECT -11.735 -271.130 -8.575 -270.960 ;
        RECT -5.240 -271.130 -5.045 -270.515 ;
        RECT -4.730 -270.760 -4.560 -269.535 ;
        RECT -3.165 -269.565 -2.980 -269.460 ;
        RECT -3.150 -270.575 -2.980 -269.565 ;
        RECT -2.670 -269.580 -1.170 -269.385 ;
        RECT -2.660 -270.575 -2.490 -269.580 ;
        RECT -1.340 -270.575 -1.170 -269.580 ;
        RECT -0.850 -270.575 -0.680 -269.120 ;
        RECT 0.130 -270.490 0.300 -269.535 ;
        RECT 0.130 -270.760 0.310 -270.490 ;
        RECT 0.620 -270.575 0.790 -269.120 ;
        RECT 1.655 -269.165 1.870 -267.470 ;
        RECT 3.205 -268.445 3.420 -267.460 ;
        RECT 7.280 -267.545 7.450 -265.985 ;
        RECT 6.580 -267.725 6.750 -267.720 ;
        RECT 7.770 -267.725 7.940 -266.505 ;
        RECT 8.260 -267.545 8.430 -265.985 ;
        RECT 8.860 -266.330 10.570 -266.160 ;
        RECT 8.860 -267.545 9.030 -266.330 ;
        RECT 9.350 -267.725 9.520 -266.505 ;
        RECT 9.840 -267.545 10.010 -266.330 ;
        RECT 6.580 -267.895 10.095 -267.725 ;
        RECT 3.640 -268.375 4.335 -268.105 ;
        RECT 2.705 -268.675 3.420 -268.445 ;
        RECT 2.075 -269.115 2.770 -268.845 ;
        RECT 1.175 -269.395 1.870 -269.165 ;
        RECT 1.655 -269.620 1.870 -269.395 ;
        RECT 1.680 -270.575 1.850 -269.620 ;
        RECT 2.170 -270.540 2.340 -269.535 ;
        RECT 3.205 -269.630 3.420 -268.675 ;
        RECT -4.730 -270.940 0.310 -270.760 ;
        RECT 2.145 -270.960 2.360 -270.540 ;
        RECT 3.225 -270.575 3.395 -269.630 ;
        RECT 3.715 -270.530 3.885 -269.535 ;
        RECT 6.580 -269.730 6.750 -267.895 ;
        RECT 7.275 -268.565 7.970 -268.295 ;
        RECT 9.925 -268.470 10.095 -267.895 ;
        RECT 10.400 -268.090 10.570 -266.330 ;
        RECT 10.750 -267.720 10.920 -265.985 ;
        RECT 19.780 -265.985 23.420 -265.815 ;
        RECT 11.650 -267.720 11.820 -266.505 ;
        RECT 10.750 -267.890 11.820 -267.720 ;
        RECT 12.630 -268.090 12.800 -266.505 ;
        RECT 14.180 -267.470 14.350 -266.505 ;
        RECT 15.725 -267.460 15.895 -266.505 ;
        RECT 10.400 -268.260 12.800 -268.090 ;
        RECT 13.065 -268.345 13.760 -268.075 ;
        RECT 9.925 -268.640 10.655 -268.470 ;
        RECT 7.270 -269.155 8.925 -268.970 ;
        RECT 9.185 -269.085 9.880 -268.815 ;
        RECT 10.485 -268.950 10.655 -268.640 ;
        RECT 11.020 -268.715 11.715 -268.445 ;
        RECT 10.485 -269.120 13.290 -268.950 ;
        RECT 7.270 -269.570 7.455 -269.155 ;
        RECT 8.740 -269.275 8.925 -269.155 ;
        RECT 8.740 -269.460 9.520 -269.275 ;
        RECT 6.550 -270.410 6.780 -269.730 ;
        RECT 7.280 -270.515 7.450 -269.570 ;
        RECT 3.690 -270.960 3.905 -270.530 ;
        RECT 0.765 -271.130 3.925 -270.960 ;
        RECT 7.260 -271.130 7.455 -270.515 ;
        RECT 7.770 -270.760 7.940 -269.535 ;
        RECT 9.335 -269.565 9.520 -269.460 ;
        RECT 9.350 -270.575 9.520 -269.565 ;
        RECT 9.830 -269.580 11.330 -269.385 ;
        RECT 9.840 -270.575 10.010 -269.580 ;
        RECT 11.160 -270.575 11.330 -269.580 ;
        RECT 11.650 -270.575 11.820 -269.120 ;
        RECT 12.630 -270.490 12.800 -269.535 ;
        RECT 12.630 -270.760 12.810 -270.490 ;
        RECT 13.120 -270.575 13.290 -269.120 ;
        RECT 14.155 -269.165 14.370 -267.470 ;
        RECT 15.705 -268.445 15.920 -267.460 ;
        RECT 19.780 -267.545 19.950 -265.985 ;
        RECT 20.270 -267.725 20.440 -266.505 ;
        RECT 20.760 -267.545 20.930 -265.985 ;
        RECT 21.360 -266.330 23.070 -266.160 ;
        RECT 21.360 -267.545 21.530 -266.330 ;
        RECT 21.850 -267.725 22.020 -266.505 ;
        RECT 22.340 -267.545 22.510 -266.330 ;
        RECT 18.660 -267.895 22.595 -267.725 ;
        RECT 16.140 -268.375 16.835 -268.105 ;
        RECT 15.205 -268.675 15.920 -268.445 ;
        RECT 14.575 -269.115 15.270 -268.845 ;
        RECT 13.675 -269.395 14.370 -269.165 ;
        RECT 14.155 -269.620 14.370 -269.395 ;
        RECT 14.180 -270.575 14.350 -269.620 ;
        RECT 14.670 -270.540 14.840 -269.535 ;
        RECT 15.705 -269.630 15.920 -268.675 ;
        RECT 7.770 -270.940 12.810 -270.760 ;
        RECT 14.645 -270.960 14.860 -270.540 ;
        RECT 15.725 -270.575 15.895 -269.630 ;
        RECT 16.215 -270.530 16.385 -269.535 ;
        RECT 18.660 -269.725 18.830 -267.895 ;
        RECT 19.775 -268.565 20.470 -268.295 ;
        RECT 22.425 -268.470 22.595 -267.895 ;
        RECT 22.900 -268.090 23.070 -266.330 ;
        RECT 23.250 -267.720 23.420 -265.985 ;
        RECT 34.780 -265.985 38.420 -265.815 ;
        RECT 24.150 -267.720 24.320 -266.505 ;
        RECT 23.250 -267.890 24.320 -267.720 ;
        RECT 25.130 -268.090 25.300 -266.505 ;
        RECT 26.680 -267.470 26.850 -266.505 ;
        RECT 28.225 -267.460 28.395 -266.505 ;
        RECT 22.900 -268.260 25.300 -268.090 ;
        RECT 25.565 -268.345 26.260 -268.075 ;
        RECT 22.425 -268.640 23.155 -268.470 ;
        RECT 22.985 -268.950 23.155 -268.640 ;
        RECT 23.520 -268.715 24.215 -268.445 ;
        RECT 19.770 -269.155 21.425 -268.970 ;
        RECT 22.985 -269.120 25.790 -268.950 ;
        RECT 19.770 -269.570 19.955 -269.155 ;
        RECT 21.240 -269.275 21.425 -269.155 ;
        RECT 21.240 -269.460 22.020 -269.275 ;
        RECT 18.660 -269.730 18.835 -269.725 ;
        RECT 18.635 -270.410 18.865 -269.730 ;
        RECT 19.780 -270.515 19.950 -269.570 ;
        RECT 16.190 -270.960 16.405 -270.530 ;
        RECT 13.265 -271.130 16.425 -270.960 ;
        RECT 19.760 -271.130 19.955 -270.515 ;
        RECT 20.270 -270.760 20.440 -269.535 ;
        RECT 21.835 -269.565 22.020 -269.460 ;
        RECT 21.850 -270.575 22.020 -269.565 ;
        RECT 22.330 -269.580 23.830 -269.385 ;
        RECT 22.340 -270.575 22.510 -269.580 ;
        RECT 23.660 -270.575 23.830 -269.580 ;
        RECT 24.150 -270.575 24.320 -269.120 ;
        RECT 25.130 -270.490 25.300 -269.535 ;
        RECT 25.130 -270.760 25.310 -270.490 ;
        RECT 25.620 -270.575 25.790 -269.120 ;
        RECT 26.655 -269.165 26.870 -267.470 ;
        RECT 28.205 -268.445 28.420 -267.460 ;
        RECT 34.780 -267.545 34.950 -265.985 ;
        RECT 35.270 -267.725 35.440 -266.505 ;
        RECT 35.760 -267.545 35.930 -265.985 ;
        RECT 36.360 -266.330 38.070 -266.160 ;
        RECT 36.360 -267.545 36.530 -266.330 ;
        RECT 36.850 -267.725 37.020 -266.505 ;
        RECT 37.340 -267.545 37.510 -266.330 ;
        RECT 33.190 -267.895 37.595 -267.725 ;
        RECT 28.640 -268.375 29.335 -268.105 ;
        RECT 27.705 -268.675 28.420 -268.445 ;
        RECT 26.175 -269.395 26.870 -269.165 ;
        RECT 26.655 -269.620 26.870 -269.395 ;
        RECT 26.680 -270.575 26.850 -269.620 ;
        RECT 27.170 -270.540 27.340 -269.535 ;
        RECT 28.205 -269.630 28.420 -268.675 ;
        RECT 20.270 -270.940 25.310 -270.760 ;
        RECT 27.145 -270.960 27.360 -270.540 ;
        RECT 28.225 -270.575 28.395 -269.630 ;
        RECT 28.715 -270.530 28.885 -269.535 ;
        RECT 33.190 -269.730 33.360 -267.895 ;
        RECT 34.775 -268.565 35.470 -268.295 ;
        RECT 37.425 -268.470 37.595 -267.895 ;
        RECT 37.900 -268.090 38.070 -266.330 ;
        RECT 38.250 -267.720 38.420 -265.985 ;
        RECT 39.150 -267.720 39.320 -266.505 ;
        RECT 38.250 -267.890 39.320 -267.720 ;
        RECT 40.130 -268.090 40.300 -266.505 ;
        RECT 41.680 -267.470 41.850 -266.505 ;
        RECT 43.225 -267.460 43.395 -266.505 ;
        RECT 37.900 -268.260 40.300 -268.090 ;
        RECT 40.565 -268.345 41.260 -268.075 ;
        RECT 37.425 -268.640 38.155 -268.470 ;
        RECT 37.985 -268.950 38.155 -268.640 ;
        RECT 38.520 -268.715 39.215 -268.445 ;
        RECT 34.770 -269.155 36.425 -268.970 ;
        RECT 37.985 -269.120 40.790 -268.950 ;
        RECT 34.770 -269.570 34.955 -269.155 ;
        RECT 36.240 -269.275 36.425 -269.155 ;
        RECT 36.240 -269.460 37.020 -269.275 ;
        RECT 33.160 -270.410 33.390 -269.730 ;
        RECT 34.780 -270.515 34.950 -269.570 ;
        RECT 28.690 -270.960 28.905 -270.530 ;
        RECT 25.765 -271.130 28.925 -270.960 ;
        RECT 34.760 -271.130 34.955 -270.515 ;
        RECT 35.270 -270.760 35.440 -269.535 ;
        RECT 36.835 -269.565 37.020 -269.460 ;
        RECT 36.850 -270.575 37.020 -269.565 ;
        RECT 37.330 -269.580 38.830 -269.385 ;
        RECT 37.340 -270.575 37.510 -269.580 ;
        RECT 38.660 -270.575 38.830 -269.580 ;
        RECT 39.150 -270.575 39.320 -269.120 ;
        RECT 40.130 -270.490 40.300 -269.535 ;
        RECT 40.130 -270.760 40.310 -270.490 ;
        RECT 40.620 -270.575 40.790 -269.120 ;
        RECT 41.655 -269.165 41.870 -267.470 ;
        RECT 43.205 -268.445 43.420 -267.460 ;
        RECT 43.640 -268.375 44.335 -268.105 ;
        RECT 42.705 -268.675 43.420 -268.445 ;
        RECT 41.175 -269.395 41.870 -269.165 ;
        RECT 41.655 -269.620 41.870 -269.395 ;
        RECT 41.680 -270.575 41.850 -269.620 ;
        RECT 42.170 -270.540 42.340 -269.535 ;
        RECT 43.205 -269.630 43.420 -268.675 ;
        RECT 35.270 -270.940 40.310 -270.760 ;
        RECT 42.145 -270.870 42.360 -270.540 ;
        RECT 43.225 -270.575 43.395 -269.630 ;
        RECT 43.715 -270.530 43.885 -269.535 ;
        RECT 43.690 -270.870 43.905 -270.530 ;
        RECT 44.720 -270.870 46.025 -261.565 ;
        RECT 87.795 -263.185 88.780 -262.280 ;
        RECT 86.075 -265.560 87.480 -264.515 ;
        RECT 47.145 -266.575 48.145 -266.405 ;
        RECT 84.275 -266.575 86.085 -266.345 ;
        RECT 47.145 -267.435 86.085 -266.575 ;
        RECT 47.145 -268.260 48.145 -267.435 ;
        RECT 84.275 -267.700 86.085 -267.435 ;
        RECT 40.685 -271.130 46.025 -270.870 ;
        RECT 83.075 -271.065 84.535 -271.060 ;
        RECT -30.240 -271.390 46.025 -271.130 ;
        RECT -30.240 -271.395 -21.075 -271.390 ;
        RECT -17.740 -271.395 46.025 -271.390 ;
        RECT -28.080 -271.495 -25.410 -271.395 ;
        RECT -24.235 -271.440 -21.075 -271.395 ;
        RECT -11.735 -271.440 -8.575 -271.395 ;
        RECT 0.765 -271.440 3.925 -271.395 ;
        RECT 13.265 -271.440 16.425 -271.395 ;
        RECT 25.765 -271.440 28.925 -271.395 ;
        RECT -28.035 -272.290 -27.865 -271.495 ;
        RECT -27.545 -272.210 -27.375 -271.750 ;
        RECT -27.575 -272.675 -27.345 -272.210 ;
        RECT -27.055 -272.290 -26.885 -271.495 ;
        RECT -26.565 -272.210 -26.395 -271.750 ;
        RECT -26.595 -272.675 -26.365 -272.210 ;
        RECT -26.075 -272.290 -25.905 -271.495 ;
        RECT 40.685 -271.505 46.025 -271.395 ;
        RECT -25.585 -272.210 -25.415 -271.750 ;
        RECT -5.025 -271.820 -4.345 -271.590 ;
        RECT 7.460 -271.670 8.140 -271.655 ;
        RECT -4.590 -272.060 -4.345 -271.820 ;
        RECT 7.295 -271.840 18.150 -271.670 ;
        RECT 7.460 -271.885 8.140 -271.840 ;
        RECT -25.615 -272.515 -25.385 -272.210 ;
        RECT -20.500 -272.515 -20.270 -272.185 ;
        RECT -4.590 -272.240 17.670 -272.060 ;
        RECT -25.615 -272.675 -20.270 -272.515 ;
        RECT -27.575 -272.865 -20.270 -272.675 ;
        RECT 17.490 -272.800 17.670 -272.240 ;
        RECT 17.980 -272.460 18.150 -271.840 ;
        RECT 32.900 -271.920 33.580 -271.890 ;
        RECT 18.375 -272.015 19.055 -271.970 ;
        RECT 18.375 -272.185 32.380 -272.015 ;
        RECT 32.900 -272.090 34.260 -271.920 ;
        RECT 32.900 -272.120 33.580 -272.090 ;
        RECT 18.375 -272.200 19.055 -272.185 ;
        RECT 32.210 -272.380 32.380 -272.185 ;
        RECT 17.980 -272.630 25.490 -272.460 ;
        RECT 32.210 -272.550 33.910 -272.380 ;
        RECT -27.575 -272.905 -25.385 -272.865 ;
        RECT -27.575 -274.170 -27.345 -272.905 ;
        RECT -26.595 -273.230 -26.365 -272.905 ;
        RECT -25.615 -273.230 -25.385 -272.905 ;
        RECT 17.490 -272.980 25.095 -272.800 ;
        RECT -27.545 -274.190 -27.375 -274.170 ;
        RECT -26.565 -274.190 -26.395 -273.230 ;
        RECT -25.585 -274.190 -25.415 -273.230 ;
        RECT -18.590 -273.920 -18.360 -273.240 ;
        RECT -18.575 -275.185 -18.375 -273.920 ;
        RECT -18.575 -275.415 -17.895 -275.185 ;
        RECT 16.670 -275.405 17.350 -275.175 ;
        RECT -30.975 -275.825 -30.295 -275.595 ;
        RECT 16.150 -275.825 16.925 -275.595 ;
        RECT -24.665 -277.570 -21.525 -277.400 ;
        RECT -29.320 -278.625 -29.150 -277.665 ;
        RECT -28.340 -278.625 -28.170 -277.665 ;
        RECT -27.360 -277.685 -27.190 -277.665 ;
        RECT -29.350 -278.950 -29.120 -278.625 ;
        RECT -28.370 -278.950 -28.140 -278.625 ;
        RECT -27.390 -278.950 -27.160 -277.685 ;
        RECT -25.130 -278.240 -24.960 -277.740 ;
        RECT -24.665 -277.825 -24.455 -277.570 ;
        RECT -29.350 -278.990 -27.160 -278.950 ;
        RECT -29.500 -279.035 -27.160 -278.990 ;
        RECT -25.155 -278.460 -24.945 -278.240 ;
        RECT -24.640 -278.280 -24.470 -277.825 ;
        RECT -24.150 -278.190 -23.980 -277.740 ;
        RECT -23.685 -277.850 -23.475 -277.570 ;
        RECT -24.155 -278.460 -23.975 -278.190 ;
        RECT -23.660 -278.280 -23.490 -277.850 ;
        RECT -23.170 -278.190 -23.000 -277.740 ;
        RECT -22.715 -277.845 -22.505 -277.570 ;
        RECT -23.185 -278.280 -23.000 -278.190 ;
        RECT -22.680 -278.280 -22.510 -277.845 ;
        RECT -22.190 -278.200 -22.020 -277.740 ;
        RECT -21.705 -277.795 -21.525 -277.570 ;
        RECT -11.165 -277.570 -8.025 -277.400 ;
        RECT -21.700 -278.165 -21.530 -277.795 ;
        RECT -23.185 -278.460 -23.005 -278.280 ;
        RECT -22.195 -278.460 -22.015 -278.200 ;
        RECT -25.155 -278.630 -22.015 -278.460 ;
        RECT -29.910 -279.045 -27.160 -279.035 ;
        RECT -29.915 -279.180 -27.160 -279.045 ;
        RECT -29.915 -279.230 -29.120 -279.180 ;
        RECT -29.915 -281.020 -29.675 -279.230 ;
        RECT -29.500 -279.340 -29.120 -279.230 ;
        RECT -29.350 -279.645 -29.120 -279.340 ;
        RECT -29.320 -280.105 -29.150 -279.645 ;
        RECT -28.830 -280.360 -28.660 -279.565 ;
        RECT -28.370 -279.645 -28.140 -279.180 ;
        RECT -28.340 -280.105 -28.170 -279.645 ;
        RECT -27.850 -280.360 -27.680 -279.565 ;
        RECT -27.390 -279.645 -27.160 -279.180 ;
        RECT -26.980 -279.055 -26.140 -279.025 ;
        RECT -25.155 -279.055 -24.280 -278.630 ;
        RECT -21.735 -278.900 -21.500 -278.165 ;
        RECT -21.280 -278.870 -20.910 -278.030 ;
        RECT -20.605 -278.625 -20.435 -277.665 ;
        RECT -19.625 -278.625 -19.455 -277.665 ;
        RECT -18.645 -277.685 -18.475 -277.665 ;
        RECT -26.980 -279.320 -24.280 -279.055 ;
        RECT -22.360 -279.270 -21.500 -278.900 ;
        RECT -26.980 -279.395 -26.140 -279.320 ;
        RECT -25.155 -279.465 -24.280 -279.320 ;
        RECT -27.360 -280.105 -27.190 -279.645 ;
        RECT -26.870 -280.360 -26.700 -279.565 ;
        RECT -25.155 -279.635 -22.000 -279.465 ;
        RECT -25.155 -279.670 -24.945 -279.635 ;
        RECT -25.150 -279.885 -24.945 -279.670 ;
        RECT -25.130 -280.355 -24.960 -279.885 ;
        RECT -24.640 -280.295 -24.470 -279.815 ;
        RECT -24.165 -279.880 -23.960 -279.635 ;
        RECT -29.325 -280.700 -26.655 -280.360 ;
        RECT -24.670 -280.585 -24.450 -280.295 ;
        RECT -24.150 -280.355 -23.980 -279.880 ;
        RECT -23.660 -280.240 -23.490 -279.815 ;
        RECT -23.195 -279.880 -22.990 -279.635 ;
        RECT -23.685 -280.585 -23.465 -280.240 ;
        RECT -23.170 -280.355 -23.000 -279.880 ;
        RECT -22.680 -280.240 -22.510 -279.815 ;
        RECT -22.205 -279.840 -22.000 -279.635 ;
        RECT -22.705 -280.585 -22.485 -280.240 ;
        RECT -22.190 -280.355 -22.020 -279.840 ;
        RECT -21.735 -279.945 -21.500 -279.270 ;
        RECT -21.275 -278.990 -20.910 -278.870 ;
        RECT -20.635 -278.950 -20.405 -278.625 ;
        RECT -19.655 -278.950 -19.425 -278.625 ;
        RECT -18.675 -278.950 -18.445 -277.685 ;
        RECT -17.655 -278.165 -17.370 -277.775 ;
        RECT -17.655 -278.390 -16.350 -278.165 ;
        RECT -17.655 -278.595 -17.370 -278.390 ;
        RECT -20.635 -278.990 -18.445 -278.950 ;
        RECT -21.275 -279.180 -18.445 -278.990 ;
        RECT -21.275 -279.340 -20.405 -279.180 ;
        RECT -20.635 -279.645 -20.405 -279.340 ;
        RECT -21.700 -280.295 -21.530 -279.945 ;
        RECT -20.605 -280.105 -20.435 -279.645 ;
        RECT -21.725 -280.585 -21.505 -280.295 ;
        RECT -20.115 -280.360 -19.945 -279.565 ;
        RECT -19.655 -279.645 -19.425 -279.180 ;
        RECT -19.625 -280.105 -19.455 -279.645 ;
        RECT -19.135 -280.360 -18.965 -279.565 ;
        RECT -18.675 -279.645 -18.445 -279.180 ;
        RECT -18.265 -279.080 -17.425 -279.025 ;
        RECT -16.575 -279.060 -16.350 -278.390 ;
        RECT -15.820 -278.625 -15.650 -277.665 ;
        RECT -14.840 -278.625 -14.670 -277.665 ;
        RECT -13.860 -277.685 -13.690 -277.665 ;
        RECT -15.850 -278.950 -15.620 -278.625 ;
        RECT -14.870 -278.950 -14.640 -278.625 ;
        RECT -13.890 -278.950 -13.660 -277.685 ;
        RECT -11.630 -278.240 -11.460 -277.740 ;
        RECT -11.165 -277.825 -10.955 -277.570 ;
        RECT -15.850 -278.990 -13.660 -278.950 ;
        RECT -16.000 -279.060 -13.660 -278.990 ;
        RECT -11.655 -278.460 -11.445 -278.240 ;
        RECT -11.140 -278.280 -10.970 -277.825 ;
        RECT -10.650 -278.190 -10.480 -277.740 ;
        RECT -10.185 -277.850 -9.975 -277.570 ;
        RECT -10.655 -278.460 -10.475 -278.190 ;
        RECT -10.160 -278.280 -9.990 -277.850 ;
        RECT -9.670 -278.190 -9.500 -277.740 ;
        RECT -9.215 -277.845 -9.005 -277.570 ;
        RECT -9.685 -278.280 -9.500 -278.190 ;
        RECT -9.180 -278.280 -9.010 -277.845 ;
        RECT -8.690 -278.200 -8.520 -277.740 ;
        RECT -8.205 -277.795 -8.025 -277.570 ;
        RECT -8.200 -278.165 -8.030 -277.795 ;
        RECT -9.685 -278.460 -9.505 -278.280 ;
        RECT -8.695 -278.460 -8.515 -278.200 ;
        RECT -11.655 -278.630 -8.515 -278.460 ;
        RECT -17.125 -279.080 -16.825 -279.075 ;
        RECT -18.265 -279.370 -16.825 -279.080 ;
        RECT -16.575 -279.180 -13.660 -279.060 ;
        RECT -16.575 -279.285 -15.620 -279.180 ;
        RECT -18.265 -279.395 -17.425 -279.370 ;
        RECT -18.645 -280.105 -18.475 -279.645 ;
        RECT -18.155 -280.360 -17.985 -279.565 ;
        RECT -17.125 -279.735 -16.825 -279.370 ;
        RECT -16.550 -279.860 -16.250 -279.285 ;
        RECT -16.000 -279.340 -15.620 -279.285 ;
        RECT -15.850 -279.645 -15.620 -279.340 ;
        RECT -15.820 -280.105 -15.650 -279.645 ;
        RECT -15.330 -280.360 -15.160 -279.565 ;
        RECT -14.870 -279.645 -14.640 -279.180 ;
        RECT -14.840 -280.105 -14.670 -279.645 ;
        RECT -14.350 -280.360 -14.180 -279.565 ;
        RECT -13.890 -279.645 -13.660 -279.180 ;
        RECT -13.480 -279.070 -12.640 -279.025 ;
        RECT -11.655 -279.070 -10.780 -278.630 ;
        RECT -8.235 -278.900 -8.000 -278.165 ;
        RECT -7.780 -278.870 -7.410 -278.030 ;
        RECT -7.105 -278.625 -6.935 -277.665 ;
        RECT -6.125 -278.625 -5.955 -277.665 ;
        RECT -5.145 -277.685 -4.975 -277.665 ;
        RECT -13.480 -279.355 -10.780 -279.070 ;
        RECT -8.860 -279.270 -8.000 -278.900 ;
        RECT -13.480 -279.395 -12.640 -279.355 ;
        RECT -11.655 -279.465 -10.780 -279.355 ;
        RECT -13.860 -280.105 -13.690 -279.645 ;
        RECT -13.370 -280.360 -13.200 -279.565 ;
        RECT -11.655 -279.635 -8.500 -279.465 ;
        RECT -11.655 -279.670 -11.445 -279.635 ;
        RECT -11.650 -279.835 -11.445 -279.670 ;
        RECT -11.650 -279.885 -11.415 -279.835 ;
        RECT -24.670 -280.755 -21.505 -280.585 ;
        RECT -20.610 -280.700 -13.155 -280.360 ;
        RECT -11.645 -280.495 -11.415 -279.885 ;
        RECT -11.140 -280.295 -10.970 -279.815 ;
        RECT -10.665 -279.880 -10.460 -279.635 ;
        RECT -11.170 -280.585 -10.950 -280.295 ;
        RECT -10.650 -280.355 -10.480 -279.880 ;
        RECT -10.160 -280.240 -9.990 -279.815 ;
        RECT -9.695 -279.880 -9.490 -279.635 ;
        RECT -10.185 -280.585 -9.965 -280.240 ;
        RECT -9.670 -280.355 -9.500 -279.880 ;
        RECT -9.180 -280.240 -9.010 -279.815 ;
        RECT -8.705 -279.840 -8.500 -279.635 ;
        RECT -9.205 -280.585 -8.985 -280.240 ;
        RECT -8.690 -280.355 -8.520 -279.840 ;
        RECT -8.235 -279.945 -8.000 -279.270 ;
        RECT -7.775 -278.990 -7.410 -278.870 ;
        RECT -7.135 -278.950 -6.905 -278.625 ;
        RECT -6.155 -278.950 -5.925 -278.625 ;
        RECT -5.175 -278.950 -4.945 -277.685 ;
        RECT -4.155 -278.595 -3.870 -277.775 ;
        RECT -2.695 -278.625 -2.525 -277.665 ;
        RECT -1.715 -278.625 -1.545 -277.665 ;
        RECT -0.735 -277.685 -0.565 -277.665 ;
        RECT -7.135 -278.990 -4.945 -278.950 ;
        RECT -2.725 -278.950 -2.495 -278.625 ;
        RECT -1.745 -278.950 -1.515 -278.625 ;
        RECT -0.765 -278.950 -0.535 -277.685 ;
        RECT -2.725 -278.990 -0.535 -278.950 ;
        RECT -7.775 -279.180 -4.945 -278.990 ;
        RECT -7.775 -279.340 -6.905 -279.180 ;
        RECT -7.135 -279.645 -6.905 -279.340 ;
        RECT -8.200 -280.295 -8.030 -279.945 ;
        RECT -7.105 -280.105 -6.935 -279.645 ;
        RECT -8.225 -280.585 -8.005 -280.295 ;
        RECT -6.615 -280.360 -6.445 -279.565 ;
        RECT -6.155 -279.645 -5.925 -279.180 ;
        RECT -6.125 -280.105 -5.955 -279.645 ;
        RECT -5.635 -280.360 -5.465 -279.565 ;
        RECT -5.175 -279.645 -4.945 -279.180 ;
        RECT -3.465 -279.100 -3.165 -279.080 ;
        RECT -2.875 -279.100 -0.535 -278.990 ;
        RECT -3.465 -279.180 -0.535 -279.100 ;
        RECT -3.465 -279.310 -2.495 -279.180 ;
        RECT -5.145 -280.105 -4.975 -279.645 ;
        RECT -4.655 -280.360 -4.485 -279.565 ;
        RECT -3.465 -279.740 -3.165 -279.310 ;
        RECT -2.875 -279.340 -2.495 -279.310 ;
        RECT -2.725 -279.645 -2.495 -279.340 ;
        RECT -2.695 -280.105 -2.525 -279.645 ;
        RECT -2.205 -280.360 -2.035 -279.565 ;
        RECT -1.745 -279.645 -1.515 -279.180 ;
        RECT -1.715 -280.105 -1.545 -279.645 ;
        RECT -1.225 -280.360 -1.055 -279.565 ;
        RECT -0.765 -279.645 -0.535 -279.180 ;
        RECT -0.735 -280.105 -0.565 -279.645 ;
        RECT -0.245 -280.360 -0.075 -279.565 ;
        RECT 1.955 -279.800 2.125 -277.750 ;
        RECT 5.645 -278.970 5.815 -277.750 ;
        RECT 6.625 -278.970 6.795 -277.750 ;
        RECT 7.605 -278.970 7.775 -277.750 ;
        RECT 5.000 -279.155 7.775 -278.970 ;
        RECT 8.705 -278.985 8.935 -278.565 ;
        RECT 10.620 -278.675 10.790 -277.815 ;
        RECT 11.600 -278.355 11.770 -277.815 ;
        RECT 12.580 -278.355 12.750 -277.815 ;
        RECT 1.200 -280.065 2.125 -279.800 ;
        RECT 2.300 -279.845 2.975 -279.795 ;
        RECT 5.000 -279.845 5.185 -279.155 ;
        RECT 7.975 -279.255 8.935 -278.985 ;
        RECT 9.935 -279.025 10.790 -278.675 ;
        RECT 12.975 -278.590 13.340 -278.525 ;
        RECT 12.975 -278.730 13.840 -278.590 ;
        RECT 12.975 -278.795 13.950 -278.730 ;
        RECT 12.975 -278.825 13.340 -278.795 ;
        RECT 6.295 -279.440 6.970 -279.395 ;
        RECT 9.110 -279.440 9.790 -279.435 ;
        RECT 6.295 -279.630 9.790 -279.440 ;
        RECT 6.295 -279.665 6.970 -279.630 ;
        RECT 9.110 -279.665 9.790 -279.630 ;
        RECT 2.300 -280.030 5.185 -279.845 ;
        RECT 2.300 -280.065 2.975 -280.030 ;
        RECT -11.170 -280.755 -8.005 -280.585 ;
        RECT -7.110 -280.700 -0.030 -280.360 ;
        RECT -31.695 -281.465 -30.775 -281.150 ;
        RECT -31.590 -281.470 -30.775 -281.465 ;
        RECT -29.920 -281.705 -29.620 -281.020 ;
        RECT -17.370 -281.365 -16.685 -281.315 ;
        RECT -12.640 -281.365 -11.980 -281.310 ;
        RECT -2.570 -281.365 -1.910 -281.315 ;
        RECT -28.265 -281.560 -1.910 -281.365 ;
        RECT -17.370 -281.615 -16.685 -281.560 ;
        RECT -12.640 -281.610 -11.980 -281.560 ;
        RECT -2.570 -281.615 -1.910 -281.560 ;
        RECT -29.915 -283.565 -29.675 -281.705 ;
        RECT -28.180 -281.825 -27.495 -281.760 ;
        RECT -15.195 -281.825 -14.510 -281.730 ;
        RECT -1.355 -281.825 -0.695 -281.730 ;
        RECT -28.265 -282.020 -0.690 -281.825 ;
        RECT -28.180 -282.060 -27.495 -282.020 ;
        RECT -28.125 -282.260 -27.570 -282.060 ;
        RECT -24.070 -282.260 -23.515 -282.020 ;
        RECT -15.195 -282.030 -14.510 -282.020 ;
        RECT -29.365 -282.600 -22.510 -282.260 ;
        RECT -21.615 -282.375 -18.450 -282.205 ;
        RECT -15.080 -282.260 -14.525 -282.030 ;
        RECT -14.165 -282.260 -11.565 -282.250 ;
        RECT -10.690 -282.260 -10.135 -282.020 ;
        RECT -29.320 -283.395 -29.150 -282.600 ;
        RECT -28.830 -283.315 -28.660 -282.855 ;
        RECT -29.915 -283.785 -29.040 -283.565 ;
        RECT -29.880 -283.935 -29.040 -283.785 ;
        RECT -28.860 -283.780 -28.630 -283.315 ;
        RECT -28.340 -283.395 -28.170 -282.600 ;
        RECT -27.850 -283.315 -27.680 -282.855 ;
        RECT -27.880 -283.780 -27.650 -283.315 ;
        RECT -27.360 -283.395 -27.190 -282.600 ;
        RECT -26.870 -283.315 -26.700 -282.855 ;
        RECT -26.900 -283.620 -26.670 -283.315 ;
        RECT -25.135 -283.395 -24.965 -282.600 ;
        RECT -24.645 -283.315 -24.475 -282.855 ;
        RECT -26.900 -283.780 -26.235 -283.620 ;
        RECT -58.995 -285.995 -58.320 -285.965 ;
        RECT -59.095 -286.005 -58.320 -285.995 ;
        RECT -90.420 -287.205 -72.730 -286.175 ;
        RECT -60.130 -286.185 -58.320 -286.005 ;
        RECT -58.080 -286.080 -55.930 -285.930 ;
        RECT -58.080 -286.120 -55.985 -286.080 ;
        RECT -55.035 -286.140 -54.865 -285.360 ;
        RECT -54.545 -285.900 -54.375 -285.360 ;
        RECT -54.055 -286.140 -53.885 -285.360 ;
        RECT -53.565 -285.900 -53.395 -285.360 ;
        RECT -53.075 -285.415 -51.215 -285.065 ;
        RECT -28.860 -283.970 -26.235 -283.780 ;
        RECT -28.860 -284.010 -26.670 -283.970 ;
        RECT -28.860 -285.275 -28.630 -284.010 ;
        RECT -27.880 -284.335 -27.650 -284.010 ;
        RECT -26.900 -284.335 -26.670 -284.010 ;
        RECT -28.830 -285.295 -28.660 -285.275 ;
        RECT -27.850 -285.295 -27.680 -284.335 ;
        RECT -26.870 -285.295 -26.700 -284.335 ;
        RECT -26.465 -284.620 -26.235 -283.970 ;
        RECT -24.675 -283.780 -24.445 -283.315 ;
        RECT -24.155 -283.395 -23.985 -282.600 ;
        RECT -23.665 -283.315 -23.495 -282.855 ;
        RECT -23.695 -283.780 -23.465 -283.315 ;
        RECT -23.175 -283.395 -23.005 -282.600 ;
        RECT -21.615 -282.665 -21.395 -282.375 ;
        RECT -22.685 -283.315 -22.515 -282.855 ;
        RECT -21.590 -283.015 -21.420 -282.665 ;
        RECT -22.715 -283.620 -22.485 -283.315 ;
        RECT -22.715 -283.780 -21.845 -283.620 ;
        RECT -24.675 -283.970 -21.845 -283.780 ;
        RECT -24.675 -284.010 -22.485 -283.970 ;
        RECT -25.750 -284.620 -25.465 -284.365 ;
        RECT -26.465 -284.865 -25.465 -284.620 ;
        RECT -25.750 -285.185 -25.465 -284.865 ;
        RECT -24.675 -285.275 -24.445 -284.010 ;
        RECT -23.695 -284.335 -23.465 -284.010 ;
        RECT -22.715 -284.335 -22.485 -284.010 ;
        RECT -22.210 -284.090 -21.845 -283.970 ;
        RECT -21.620 -283.690 -21.385 -283.015 ;
        RECT -21.100 -283.120 -20.930 -282.605 ;
        RECT -20.635 -282.720 -20.415 -282.375 ;
        RECT -21.120 -283.325 -20.915 -283.120 ;
        RECT -20.610 -283.145 -20.440 -282.720 ;
        RECT -20.120 -283.080 -19.950 -282.605 ;
        RECT -19.655 -282.720 -19.435 -282.375 ;
        RECT -20.130 -283.325 -19.925 -283.080 ;
        RECT -19.630 -283.145 -19.460 -282.720 ;
        RECT -19.140 -283.080 -18.970 -282.605 ;
        RECT -18.670 -282.665 -18.450 -282.375 ;
        RECT -15.865 -282.590 -9.010 -282.260 ;
        RECT -15.865 -282.600 -13.195 -282.590 ;
        RECT -11.680 -282.600 -9.010 -282.590 ;
        RECT -8.115 -282.375 -4.950 -282.205 ;
        RECT -19.160 -283.325 -18.955 -283.080 ;
        RECT -18.650 -283.145 -18.480 -282.665 ;
        RECT -18.160 -283.075 -17.990 -282.605 ;
        RECT -18.175 -283.290 -17.970 -283.075 ;
        RECT -18.175 -283.325 -17.965 -283.290 ;
        RECT -21.120 -283.495 -17.965 -283.325 ;
        RECT -15.820 -283.395 -15.650 -282.600 ;
        RECT -15.330 -283.315 -15.160 -282.855 ;
        RECT -21.620 -284.060 -20.760 -283.690 ;
        RECT -18.840 -283.795 -17.510 -283.495 ;
        RECT -16.380 -283.600 -15.540 -283.565 ;
        RECT -24.645 -285.295 -24.475 -285.275 ;
        RECT -23.665 -285.295 -23.495 -284.335 ;
        RECT -22.685 -285.295 -22.515 -284.335 ;
        RECT -22.210 -284.930 -21.840 -284.090 ;
        RECT -21.620 -284.795 -21.385 -284.060 ;
        RECT -18.840 -284.330 -17.965 -283.795 ;
        RECT -16.490 -283.900 -15.540 -283.600 ;
        RECT -16.380 -283.935 -15.540 -283.900 ;
        RECT -15.360 -283.780 -15.130 -283.315 ;
        RECT -14.840 -283.395 -14.670 -282.600 ;
        RECT -14.350 -283.315 -14.180 -282.855 ;
        RECT -14.380 -283.780 -14.150 -283.315 ;
        RECT -13.860 -283.395 -13.690 -282.600 ;
        RECT -13.370 -283.315 -13.200 -282.855 ;
        RECT -13.400 -283.620 -13.170 -283.315 ;
        RECT -12.495 -283.565 -12.195 -282.770 ;
        RECT -11.635 -283.395 -11.465 -282.600 ;
        RECT -11.145 -283.315 -10.975 -282.855 ;
        RECT -13.400 -283.780 -12.680 -283.620 ;
        RECT -21.105 -284.500 -17.965 -284.330 ;
        RECT -21.105 -284.760 -20.925 -284.500 ;
        RECT -20.115 -284.680 -19.935 -284.500 ;
        RECT -21.590 -285.165 -21.420 -284.795 ;
        RECT -21.595 -285.390 -21.415 -285.165 ;
        RECT -21.100 -285.220 -20.930 -284.760 ;
        RECT -20.610 -285.115 -20.440 -284.680 ;
        RECT -20.120 -284.770 -19.935 -284.680 ;
        RECT -20.615 -285.390 -20.405 -285.115 ;
        RECT -20.120 -285.220 -19.950 -284.770 ;
        RECT -19.630 -285.110 -19.460 -284.680 ;
        RECT -19.145 -284.770 -18.965 -284.500 ;
        RECT -19.645 -285.390 -19.435 -285.110 ;
        RECT -19.140 -285.220 -18.970 -284.770 ;
        RECT -18.650 -285.135 -18.480 -284.680 ;
        RECT -18.175 -284.720 -17.965 -284.500 ;
        RECT -15.360 -283.970 -12.680 -283.780 ;
        RECT -12.495 -283.880 -11.355 -283.565 ;
        RECT -12.195 -283.935 -11.355 -283.880 ;
        RECT -11.175 -283.780 -10.945 -283.315 ;
        RECT -10.655 -283.395 -10.485 -282.600 ;
        RECT -10.165 -283.315 -9.995 -282.855 ;
        RECT -10.195 -283.780 -9.965 -283.315 ;
        RECT -9.675 -283.395 -9.505 -282.600 ;
        RECT -8.115 -282.665 -7.895 -282.375 ;
        RECT -9.185 -283.315 -9.015 -282.855 ;
        RECT -8.090 -283.015 -7.920 -282.665 ;
        RECT -9.215 -283.620 -8.985 -283.315 ;
        RECT -9.215 -283.780 -8.345 -283.620 ;
        RECT -15.360 -284.010 -13.170 -283.970 ;
        RECT -18.665 -285.390 -18.455 -285.135 ;
        RECT -18.160 -285.220 -17.990 -284.720 ;
        RECT -15.360 -285.275 -15.130 -284.010 ;
        RECT -14.380 -284.335 -14.150 -284.010 ;
        RECT -13.400 -284.335 -13.170 -284.010 ;
        RECT -15.330 -285.295 -15.160 -285.275 ;
        RECT -14.350 -285.295 -14.180 -284.335 ;
        RECT -13.370 -285.295 -13.200 -284.335 ;
        RECT -12.990 -284.615 -12.680 -283.970 ;
        RECT -11.175 -283.970 -8.345 -283.780 ;
        RECT -11.175 -284.010 -8.985 -283.970 ;
        RECT -12.250 -284.615 -11.965 -284.365 ;
        RECT -12.990 -284.925 -11.965 -284.615 ;
        RECT -12.250 -285.185 -11.965 -284.925 ;
        RECT -11.175 -285.275 -10.945 -284.010 ;
        RECT -10.195 -284.335 -9.965 -284.010 ;
        RECT -9.215 -284.335 -8.985 -284.010 ;
        RECT -8.710 -284.090 -8.345 -283.970 ;
        RECT -8.120 -283.690 -7.885 -283.015 ;
        RECT -7.600 -283.120 -7.430 -282.605 ;
        RECT -7.135 -282.720 -6.915 -282.375 ;
        RECT -7.620 -283.325 -7.415 -283.120 ;
        RECT -7.110 -283.145 -6.940 -282.720 ;
        RECT -6.620 -283.080 -6.450 -282.605 ;
        RECT -6.155 -282.720 -5.935 -282.375 ;
        RECT -6.630 -283.325 -6.425 -283.080 ;
        RECT -6.130 -283.145 -5.960 -282.720 ;
        RECT -5.640 -283.080 -5.470 -282.605 ;
        RECT -5.170 -282.665 -4.950 -282.375 ;
        RECT -5.660 -283.325 -5.455 -283.080 ;
        RECT -5.150 -283.145 -4.980 -282.665 ;
        RECT -4.660 -283.075 -4.490 -282.605 ;
        RECT -4.675 -283.290 -4.470 -283.075 ;
        RECT -4.675 -283.325 -4.465 -283.290 ;
        RECT -7.620 -283.485 -4.465 -283.325 ;
        RECT -7.620 -283.495 -4.090 -283.485 ;
        RECT -8.120 -284.060 -7.260 -283.690 ;
        RECT -5.340 -283.785 -4.090 -283.495 ;
        RECT -11.145 -285.295 -10.975 -285.275 ;
        RECT -10.165 -285.295 -9.995 -284.335 ;
        RECT -9.185 -285.295 -9.015 -284.335 ;
        RECT -8.710 -284.930 -8.340 -284.090 ;
        RECT -8.120 -284.795 -7.885 -284.060 ;
        RECT -5.340 -284.330 -4.465 -283.785 ;
        RECT -7.605 -284.500 -4.465 -284.330 ;
        RECT -7.605 -284.760 -7.425 -284.500 ;
        RECT -6.615 -284.680 -6.435 -284.500 ;
        RECT -8.090 -285.165 -7.920 -284.795 ;
        RECT -21.595 -285.560 -18.455 -285.390 ;
        RECT -8.095 -285.390 -7.915 -285.165 ;
        RECT -7.600 -285.220 -7.430 -284.760 ;
        RECT -7.110 -285.115 -6.940 -284.680 ;
        RECT -6.620 -284.770 -6.435 -284.680 ;
        RECT -7.115 -285.390 -6.905 -285.115 ;
        RECT -6.620 -285.220 -6.450 -284.770 ;
        RECT -6.130 -285.110 -5.960 -284.680 ;
        RECT -5.645 -284.770 -5.465 -284.500 ;
        RECT -6.145 -285.390 -5.935 -285.110 ;
        RECT -5.640 -285.220 -5.470 -284.770 ;
        RECT -5.150 -285.135 -4.980 -284.680 ;
        RECT -4.675 -284.720 -4.465 -284.500 ;
        RECT -5.165 -285.390 -4.955 -285.135 ;
        RECT -4.660 -285.220 -4.490 -284.720 ;
        RECT -3.270 -284.920 -1.780 -282.020 ;
        RECT -1.355 -282.030 -0.695 -282.020 ;
        RECT 1.955 -282.330 2.125 -280.065 ;
        RECT 5.000 -280.300 5.185 -280.030 ;
        RECT 5.355 -279.850 6.030 -279.785 ;
        RECT 9.965 -279.850 10.135 -279.025 ;
        RECT 11.110 -279.510 11.280 -278.970 ;
        RECT 11.600 -279.750 11.770 -278.970 ;
        RECT 12.090 -279.510 12.260 -278.970 ;
        RECT 12.580 -279.750 12.750 -278.970 ;
        RECT 13.645 -279.540 13.950 -278.795 ;
        RECT 14.645 -279.540 14.815 -277.820 ;
        RECT 15.625 -279.540 15.795 -277.820 ;
        RECT 13.645 -279.690 15.795 -279.540 ;
        RECT 16.745 -279.575 16.925 -275.825 ;
        RECT 13.700 -279.730 15.795 -279.690 ;
        RECT 16.035 -279.615 16.925 -279.575 ;
        RECT 5.355 -280.020 10.135 -279.850 ;
        RECT 5.355 -280.055 6.030 -280.020 ;
        RECT 10.375 -280.180 13.450 -279.750 ;
        RECT 16.035 -279.795 16.970 -279.615 ;
        RECT 16.035 -279.815 16.860 -279.795 ;
        RECT 16.035 -279.845 16.710 -279.815 ;
        RECT 14.015 -280.095 14.385 -279.965 ;
        RECT 17.150 -280.085 17.350 -275.405 ;
        RECT 18.645 -278.685 18.815 -277.825 ;
        RECT 19.625 -278.365 19.795 -277.825 ;
        RECT 20.605 -278.365 20.775 -277.825 ;
        RECT 16.440 -280.095 17.350 -280.085 ;
        RECT 4.020 -280.470 5.185 -280.300 ;
        RECT 6.050 -280.470 8.265 -280.300 ;
        RECT 2.445 -283.270 2.615 -281.290 ;
        RECT 4.020 -282.330 4.190 -280.470 ;
        RECT 4.510 -282.820 4.680 -280.790 ;
        RECT 5.000 -282.330 5.170 -280.470 ;
        RECT 6.050 -280.475 7.285 -280.470 ;
        RECT 6.050 -280.790 6.225 -280.475 ;
        RECT 5.565 -282.275 5.735 -280.790 ;
        RECT 5.560 -282.805 5.735 -282.275 ;
        RECT 6.055 -282.330 6.225 -280.790 ;
        RECT 6.545 -282.285 6.715 -280.790 ;
        RECT 6.540 -282.805 6.715 -282.285 ;
        RECT 7.115 -282.325 7.285 -280.475 ;
        RECT 5.560 -282.820 6.715 -282.805 ;
        RECT 4.510 -282.990 6.715 -282.820 ;
        RECT 7.605 -283.270 7.775 -280.785 ;
        RECT 8.095 -282.325 8.265 -280.470 ;
        RECT 11.925 -282.215 12.230 -280.180 ;
        RECT 14.015 -280.285 17.350 -280.095 ;
        RECT 17.825 -279.035 18.815 -278.685 ;
        RECT 21.000 -278.600 21.365 -278.535 ;
        RECT 21.000 -278.740 21.865 -278.600 ;
        RECT 21.000 -278.805 21.975 -278.740 ;
        RECT 21.000 -278.835 21.365 -278.805 ;
        RECT 14.015 -280.290 16.445 -280.285 ;
        RECT 14.015 -280.320 14.385 -280.290 ;
        RECT 16.090 -280.295 16.445 -280.290 ;
        RECT 14.155 -282.045 14.325 -280.505 ;
        RECT 14.645 -282.045 14.815 -280.505 ;
        RECT 15.135 -282.045 15.305 -280.505 ;
        RECT 15.625 -282.045 15.795 -280.505 ;
        RECT 16.115 -282.045 16.285 -280.505 ;
        RECT 11.925 -282.305 14.175 -282.215 ;
        RECT 15.625 -282.305 15.800 -282.045 ;
        RECT 11.925 -282.520 16.385 -282.305 ;
        RECT 1.895 -283.595 8.265 -283.270 ;
        RECT 1.960 -284.920 2.610 -283.595 ;
        RECT 3.490 -284.920 4.140 -283.595 ;
        RECT 5.075 -284.920 5.725 -283.595 ;
        RECT 7.305 -284.920 7.955 -283.595 ;
        RECT 11.925 -284.920 12.680 -282.520 ;
        RECT 13.810 -282.610 16.385 -282.520 ;
        RECT 13.810 -284.920 14.430 -282.610 ;
        RECT 15.460 -284.920 16.080 -282.610 ;
        RECT 17.825 -282.710 18.175 -279.035 ;
        RECT 19.135 -279.520 19.305 -278.980 ;
        RECT 19.625 -279.760 19.795 -278.980 ;
        RECT 20.115 -279.520 20.285 -278.980 ;
        RECT 20.605 -279.760 20.775 -278.980 ;
        RECT 21.670 -279.550 21.975 -278.805 ;
        RECT 22.670 -279.550 22.840 -277.830 ;
        RECT 23.650 -279.550 23.820 -277.830 ;
        RECT 21.670 -279.700 23.820 -279.550 ;
        RECT 21.725 -279.740 23.820 -279.700 ;
        RECT 24.060 -279.615 24.735 -279.585 ;
        RECT 24.915 -279.615 25.095 -272.980 ;
        RECT 18.400 -280.190 21.475 -279.760 ;
        RECT 24.060 -279.805 25.095 -279.615 ;
        RECT 24.060 -279.815 24.995 -279.805 ;
        RECT 24.060 -279.855 24.735 -279.815 ;
        RECT 22.040 -280.105 22.410 -279.975 ;
        RECT 25.290 -280.095 25.490 -272.630 ;
        RECT 24.465 -280.105 25.490 -280.095 ;
        RECT 17.495 -282.940 18.175 -282.710 ;
        RECT 19.950 -282.225 20.255 -280.190 ;
        RECT 22.040 -280.295 25.490 -280.105 ;
        RECT 22.040 -280.300 24.470 -280.295 ;
        RECT 22.040 -280.330 22.410 -280.300 ;
        RECT 24.115 -280.305 24.470 -280.300 ;
        RECT 22.180 -282.055 22.350 -280.515 ;
        RECT 22.670 -282.055 22.840 -280.515 ;
        RECT 23.160 -282.055 23.330 -280.515 ;
        RECT 23.650 -282.055 23.820 -280.515 ;
        RECT 24.140 -282.055 24.310 -280.515 ;
        RECT 26.765 -280.705 26.935 -277.705 ;
        RECT 30.455 -278.925 30.625 -277.705 ;
        RECT 31.435 -278.925 31.605 -277.705 ;
        RECT 32.415 -278.925 32.585 -277.705 ;
        RECT 29.810 -279.110 32.585 -278.925 ;
        RECT 32.785 -278.980 33.460 -278.940 ;
        RECT 27.110 -279.800 27.785 -279.750 ;
        RECT 29.810 -279.800 29.995 -279.110 ;
        RECT 32.780 -279.165 33.555 -278.980 ;
        RECT 32.780 -279.210 33.460 -279.165 ;
        RECT 31.105 -279.395 31.780 -279.350 ;
        RECT 33.740 -279.395 33.910 -272.550 ;
        RECT 31.105 -279.585 33.910 -279.395 ;
        RECT 31.105 -279.620 31.780 -279.585 ;
        RECT 27.110 -279.985 29.995 -279.800 ;
        RECT 27.110 -280.020 27.785 -279.985 ;
        RECT 29.810 -280.255 29.995 -279.985 ;
        RECT 30.165 -279.805 30.840 -279.740 ;
        RECT 34.090 -279.805 34.260 -272.090 ;
        RECT 34.830 -277.240 38.470 -277.070 ;
        RECT 34.830 -278.800 35.000 -277.240 ;
        RECT 35.320 -278.980 35.490 -277.760 ;
        RECT 35.810 -278.800 35.980 -277.240 ;
        RECT 36.410 -277.585 38.120 -277.415 ;
        RECT 36.410 -278.800 36.580 -277.585 ;
        RECT 36.900 -278.980 37.070 -277.760 ;
        RECT 37.390 -278.800 37.560 -277.585 ;
        RECT 34.575 -279.150 37.645 -278.980 ;
        RECT 30.165 -279.975 34.260 -279.805 ;
        RECT 34.825 -279.820 35.520 -279.550 ;
        RECT 37.475 -279.725 37.645 -279.150 ;
        RECT 37.950 -279.345 38.120 -277.585 ;
        RECT 38.300 -278.975 38.470 -277.240 ;
        RECT 39.200 -278.975 39.370 -277.760 ;
        RECT 38.300 -279.145 39.370 -278.975 ;
        RECT 40.180 -279.345 40.350 -277.760 ;
        RECT 41.730 -278.725 41.900 -277.760 ;
        RECT 43.275 -278.715 43.445 -277.760 ;
        RECT 37.950 -279.515 40.350 -279.345 ;
        RECT 40.615 -279.600 41.310 -279.330 ;
        RECT 37.475 -279.895 38.205 -279.725 ;
        RECT 30.165 -280.010 30.840 -279.975 ;
        RECT 38.035 -280.205 38.205 -279.895 ;
        RECT 38.570 -279.970 39.265 -279.700 ;
        RECT 25.685 -280.995 26.935 -280.705 ;
        RECT 19.950 -282.315 22.200 -282.225 ;
        RECT 23.650 -282.315 23.825 -282.055 ;
        RECT 19.950 -282.530 24.410 -282.315 ;
        RECT 19.950 -284.920 20.705 -282.530 ;
        RECT 22.160 -282.620 24.410 -282.530 ;
        RECT 22.160 -284.920 22.915 -282.620 ;
        RECT 23.625 -284.920 24.380 -282.620 ;
        RECT 25.685 -283.270 26.010 -280.995 ;
        RECT 26.765 -282.285 26.935 -280.995 ;
        RECT 28.830 -280.425 29.995 -280.255 ;
        RECT 30.860 -280.425 33.075 -280.255 ;
        RECT 27.255 -283.225 27.425 -281.245 ;
        RECT 28.830 -282.285 29.000 -280.425 ;
        RECT 29.320 -282.775 29.490 -280.745 ;
        RECT 29.810 -282.285 29.980 -280.425 ;
        RECT 30.860 -280.430 32.095 -280.425 ;
        RECT 30.860 -280.745 31.035 -280.430 ;
        RECT 30.375 -282.230 30.545 -280.745 ;
        RECT 30.370 -282.760 30.545 -282.230 ;
        RECT 30.865 -282.285 31.035 -280.745 ;
        RECT 31.355 -282.240 31.525 -280.745 ;
        RECT 31.350 -282.760 31.525 -282.240 ;
        RECT 31.925 -282.280 32.095 -280.430 ;
        RECT 30.370 -282.775 31.525 -282.760 ;
        RECT 29.320 -282.945 31.525 -282.775 ;
        RECT 32.415 -283.225 32.585 -280.740 ;
        RECT 32.905 -282.280 33.075 -280.425 ;
        RECT 34.820 -280.410 36.475 -280.225 ;
        RECT 38.035 -280.375 40.840 -280.205 ;
        RECT 34.820 -280.825 35.005 -280.410 ;
        RECT 36.290 -280.530 36.475 -280.410 ;
        RECT 36.290 -280.715 37.070 -280.530 ;
        RECT 34.830 -281.770 35.000 -280.825 ;
        RECT 34.810 -282.385 35.005 -281.770 ;
        RECT 35.320 -282.015 35.490 -280.790 ;
        RECT 36.885 -280.820 37.070 -280.715 ;
        RECT 36.900 -281.830 37.070 -280.820 ;
        RECT 37.380 -280.835 38.880 -280.640 ;
        RECT 37.390 -281.830 37.560 -280.835 ;
        RECT 38.710 -281.830 38.880 -280.835 ;
        RECT 39.200 -281.830 39.370 -280.375 ;
        RECT 40.180 -281.745 40.350 -280.790 ;
        RECT 40.180 -282.015 40.360 -281.745 ;
        RECT 40.670 -281.830 40.840 -280.375 ;
        RECT 41.705 -280.420 41.920 -278.725 ;
        RECT 43.255 -279.700 43.470 -278.715 ;
        RECT 43.690 -279.630 44.385 -279.360 ;
        RECT 42.755 -279.930 43.470 -279.700 ;
        RECT 41.225 -280.650 41.920 -280.420 ;
        RECT 41.705 -280.875 41.920 -280.650 ;
        RECT 41.730 -281.830 41.900 -280.875 ;
        RECT 42.220 -281.795 42.390 -280.790 ;
        RECT 43.255 -280.885 43.470 -279.930 ;
        RECT 35.320 -282.195 40.360 -282.015 ;
        RECT 42.195 -282.215 42.410 -281.795 ;
        RECT 43.275 -281.830 43.445 -280.885 ;
        RECT 43.765 -281.785 43.935 -280.790 ;
        RECT 43.740 -282.215 43.955 -281.785 ;
        RECT 40.815 -282.385 43.975 -282.215 ;
        RECT 34.810 -282.650 43.975 -282.385 ;
        RECT 25.335 -283.500 26.015 -283.270 ;
        RECT 26.705 -283.550 33.075 -283.225 ;
        RECT 26.825 -284.920 27.555 -283.550 ;
        RECT 29.050 -284.920 29.780 -283.550 ;
        RECT 30.380 -284.920 31.110 -283.550 ;
        RECT 32.180 -284.920 32.910 -283.550 ;
        RECT 35.000 -284.920 35.985 -282.650 ;
        RECT 37.665 -284.920 38.650 -282.650 ;
        RECT 40.230 -282.695 43.975 -282.650 ;
        RECT 40.230 -284.920 41.215 -282.695 ;
        RECT 42.745 -284.920 43.730 -282.695 ;
        RECT 44.720 -284.920 46.025 -271.505 ;
        RECT 48.205 -271.760 84.535 -271.065 ;
        RECT 82.910 -276.160 84.245 -275.980 ;
        RECT 56.185 -277.335 84.245 -276.160 ;
        RECT 82.910 -277.470 84.245 -277.335 ;
        RECT 48.345 -279.130 49.435 -279.090 ;
        RECT 84.225 -279.130 84.990 -278.935 ;
        RECT 48.345 -279.505 84.990 -279.130 ;
        RECT 48.345 -279.535 49.435 -279.505 ;
        RECT 84.225 -279.690 84.990 -279.505 ;
        RECT 53.255 -280.235 53.505 -280.205 ;
        RECT 80.815 -280.235 81.305 -280.165 ;
        RECT 53.210 -280.850 81.305 -280.235 ;
        RECT 53.255 -280.870 53.505 -280.850 ;
        RECT 80.815 -280.985 81.305 -280.850 ;
        RECT 85.400 -282.260 86.040 -267.700 ;
        RECT 86.665 -281.815 87.325 -265.560 ;
        RECT 87.875 -278.935 88.320 -263.185 ;
        RECT 98.335 -269.255 101.060 -261.565 ;
        RECT 95.420 -271.785 425.285 -269.255 ;
        RECT 87.875 -279.690 88.360 -278.935 ;
        RECT 98.335 -279.105 101.060 -271.785 ;
        RECT 147.065 -274.090 148.480 -271.785 ;
        RECT 145.845 -274.230 149.170 -274.090 ;
        RECT 173.905 -274.165 175.690 -273.830 ;
        RECT 179.795 -274.165 181.580 -274.000 ;
        RECT 189.060 -274.145 190.475 -271.785 ;
        RECT 145.845 -274.520 151.020 -274.230 ;
        RECT 145.845 -274.925 146.275 -274.520 ;
        RECT 147.145 -274.705 147.320 -274.520 ;
        RECT 148.770 -274.535 151.020 -274.520 ;
        RECT 141.585 -275.355 146.275 -274.925 ;
        RECT 140.825 -276.805 141.475 -276.345 ;
        RECT 142.285 -276.635 142.455 -275.355 ;
        RECT 142.775 -276.635 142.945 -275.595 ;
        RECT 143.265 -276.635 143.435 -275.355 ;
        RECT 143.755 -276.465 143.925 -275.595 ;
        RECT 146.660 -276.245 146.830 -274.705 ;
        RECT 147.150 -276.245 147.320 -274.705 ;
        RECT 147.640 -276.245 147.810 -274.705 ;
        RECT 148.130 -276.245 148.300 -274.705 ;
        RECT 148.620 -276.245 148.790 -274.705 ;
        RECT 146.500 -276.460 146.855 -276.455 ;
        RECT 148.560 -276.460 148.930 -276.430 ;
        RECT 146.500 -276.465 148.930 -276.460 ;
        RECT 143.755 -276.635 148.930 -276.465 ;
        RECT 150.715 -276.570 151.020 -274.535 ;
        RECT 173.905 -275.110 181.580 -274.165 ;
        RECT 188.045 -274.285 191.370 -274.145 ;
        RECT 188.045 -274.575 193.220 -274.285 ;
        RECT 233.620 -274.340 235.035 -271.785 ;
        RECT 279.715 -274.170 281.130 -271.785 ;
        RECT 306.460 -274.010 308.340 -273.535 ;
        RECT 323.690 -273.840 325.225 -271.785 ;
        RECT 314.465 -274.010 315.715 -273.875 ;
        RECT 188.045 -274.980 188.475 -274.575 ;
        RECT 189.345 -274.760 189.520 -274.575 ;
        RECT 190.970 -274.590 193.220 -274.575 ;
        RECT 173.905 -275.165 175.690 -275.110 ;
        RECT 179.795 -275.335 181.580 -275.110 ;
        RECT 183.785 -275.410 188.475 -274.980 ;
        RECT 143.760 -276.655 148.930 -276.635 ;
        RECT 143.760 -276.665 146.505 -276.655 ;
        RECT 141.695 -276.805 142.060 -276.775 ;
        RECT 148.560 -276.785 148.930 -276.655 ;
        RECT 140.825 -277.010 142.060 -276.805 ;
        RECT 149.495 -277.000 153.420 -276.570 ;
        RECT 183.025 -276.860 183.675 -276.400 ;
        RECT 184.485 -276.690 184.655 -275.410 ;
        RECT 184.975 -276.690 185.145 -275.650 ;
        RECT 185.465 -276.690 185.635 -275.410 ;
        RECT 185.955 -276.520 186.125 -275.650 ;
        RECT 188.860 -276.300 189.030 -274.760 ;
        RECT 189.350 -276.300 189.520 -274.760 ;
        RECT 189.840 -276.300 190.010 -274.760 ;
        RECT 190.330 -276.300 190.500 -274.760 ;
        RECT 190.820 -276.300 190.990 -274.760 ;
        RECT 188.700 -276.515 189.055 -276.510 ;
        RECT 190.760 -276.515 191.130 -276.485 ;
        RECT 188.700 -276.520 191.130 -276.515 ;
        RECT 185.955 -276.690 191.130 -276.520 ;
        RECT 192.915 -276.625 193.220 -274.590 ;
        RECT 216.685 -274.610 218.010 -274.455 ;
        RECT 224.315 -274.610 225.800 -274.445 ;
        RECT 216.685 -275.445 225.800 -274.610 ;
        RECT 232.360 -274.480 235.685 -274.340 ;
        RECT 232.360 -274.770 237.535 -274.480 ;
        RECT 232.360 -275.175 232.790 -274.770 ;
        RECT 233.660 -274.955 233.835 -274.770 ;
        RECT 235.285 -274.785 237.535 -274.770 ;
        RECT 216.685 -275.780 218.010 -275.445 ;
        RECT 224.315 -275.555 225.800 -275.445 ;
        RECT 228.100 -275.605 232.790 -275.175 ;
        RECT 185.960 -276.710 191.130 -276.690 ;
        RECT 185.960 -276.720 188.705 -276.710 ;
        RECT 183.895 -276.860 184.260 -276.830 ;
        RECT 190.760 -276.840 191.130 -276.710 ;
        RECT 140.825 -277.095 141.475 -277.010 ;
        RECT 141.695 -277.075 142.060 -277.010 ;
        RECT 147.150 -277.060 149.245 -277.020 ;
        RECT 147.150 -277.210 149.300 -277.060 ;
        RECT 142.285 -278.285 142.455 -277.245 ;
        RECT 143.265 -278.285 143.435 -277.245 ;
        RECT 144.245 -278.285 144.415 -277.245 ;
        RECT 105.385 -278.915 108.525 -278.745 ;
        RECT 93.845 -279.635 102.695 -279.105 ;
        RECT 104.920 -279.585 105.090 -279.085 ;
        RECT 105.385 -279.170 105.595 -278.915 ;
        RECT 87.875 -281.355 88.320 -279.690 ;
        RECT 94.365 -280.365 94.605 -279.635 ;
        RECT 94.390 -281.220 94.560 -280.365 ;
        RECT 94.880 -281.135 95.050 -280.180 ;
        RECT 95.335 -280.380 95.575 -279.635 ;
        RECT 93.460 -281.355 94.185 -281.320 ;
        RECT 87.875 -281.560 94.185 -281.355 ;
        RECT 93.460 -281.600 94.185 -281.560 ;
        RECT 94.860 -281.390 95.070 -281.135 ;
        RECT 95.370 -281.220 95.540 -280.380 ;
        RECT 95.860 -281.135 96.030 -280.180 ;
        RECT 95.840 -281.390 96.050 -281.135 ;
        RECT 94.860 -281.600 98.790 -281.390 ;
        RECT 98.095 -281.690 98.790 -281.600 ;
        RECT 95.105 -281.815 95.830 -281.795 ;
        RECT 86.665 -282.020 95.830 -281.815 ;
        RECT 95.105 -282.075 95.830 -282.020 ;
        RECT 96.705 -282.235 97.430 -281.955 ;
        RECT 96.705 -282.260 97.005 -282.235 ;
        RECT 85.400 -282.465 97.005 -282.260 ;
        RECT 98.095 -282.600 98.305 -281.690 ;
        RECT 94.370 -282.830 96.615 -282.645 ;
        RECT 94.370 -283.085 94.575 -282.830 ;
        RECT 95.425 -283.050 95.635 -282.830 ;
        RECT -8.095 -285.560 -4.955 -285.390 ;
        RECT -59.095 -286.195 -58.320 -286.185 ;
        RECT -58.995 -286.235 -58.320 -286.195 ;
        RECT -61.470 -286.485 -58.725 -286.475 ;
        RECT -56.670 -286.485 -56.300 -286.355 ;
        RECT -61.470 -286.505 -56.300 -286.485 ;
        RECT -73.770 -287.215 -72.730 -287.205 ;
        RECT -62.945 -287.785 -62.775 -286.505 ;
        RECT -62.455 -287.545 -62.285 -286.505 ;
        RECT -61.965 -287.785 -61.795 -286.505 ;
        RECT -61.475 -286.675 -56.300 -286.505 ;
        RECT -55.735 -286.570 -51.810 -286.140 ;
        RECT -3.270 -286.225 46.025 -284.920 ;
        RECT 94.390 -286.040 94.560 -283.085 ;
        RECT 95.450 -286.040 95.620 -283.050 ;
        RECT 95.940 -286.010 96.110 -283.000 ;
        RECT 96.405 -283.055 96.615 -282.830 ;
        RECT 97.465 -282.810 98.305 -282.600 ;
        RECT -61.475 -287.545 -61.305 -286.675 ;
        RECT -58.730 -286.680 -56.300 -286.675 ;
        RECT -58.730 -286.685 -58.375 -286.680 ;
        RECT -56.670 -286.710 -56.300 -286.680 ;
        RECT -63.645 -288.215 -58.955 -287.785 ;
        RECT -78.465 -288.505 -77.125 -288.270 ;
        RECT -136.180 -304.255 -132.060 -303.680 ;
        RECT -115.480 -289.435 -77.125 -288.505 ;
        RECT -59.385 -288.620 -58.955 -288.215 ;
        RECT -58.570 -288.435 -58.400 -286.895 ;
        RECT -58.080 -288.435 -57.910 -286.895 ;
        RECT -57.590 -288.435 -57.420 -286.895 ;
        RECT -57.100 -288.435 -56.930 -286.895 ;
        RECT -56.610 -288.435 -56.440 -286.895 ;
        RECT -58.085 -288.620 -57.910 -288.435 ;
        RECT -54.515 -288.605 -54.210 -286.570 ;
        RECT -56.460 -288.620 -54.210 -288.605 ;
        RECT -59.385 -288.910 -54.210 -288.620 ;
        RECT -59.385 -289.050 -56.060 -288.910 ;
        RECT -136.180 -304.965 -134.480 -304.255 ;
        RECT -115.480 -311.360 -114.550 -289.435 ;
        RECT -78.465 -289.595 -77.125 -289.435 ;
        RECT -60.965 -290.015 -57.825 -289.845 ;
        RECT -68.200 -290.130 -68.030 -290.110 ;
        RECT -68.230 -291.395 -68.000 -290.130 ;
        RECT -67.220 -291.070 -67.050 -290.110 ;
        RECT -66.240 -291.070 -66.070 -290.110 ;
        RECT -64.015 -290.130 -63.845 -290.110 ;
        RECT -65.120 -290.540 -64.835 -290.220 ;
        RECT -65.835 -290.785 -64.835 -290.540 ;
        RECT -67.250 -291.395 -67.020 -291.070 ;
        RECT -66.270 -291.395 -66.040 -291.070 ;
        RECT -68.230 -291.435 -66.040 -291.395 ;
        RECT -65.835 -291.435 -65.605 -290.785 ;
        RECT -65.120 -291.040 -64.835 -290.785 ;
        RECT -69.250 -291.620 -68.410 -291.470 ;
        RECT -69.285 -291.840 -68.410 -291.620 ;
        RECT -68.230 -291.625 -65.605 -291.435 ;
        RECT -64.045 -291.395 -63.815 -290.130 ;
        RECT -63.035 -291.070 -62.865 -290.110 ;
        RECT -62.055 -291.070 -61.885 -290.110 ;
        RECT -60.965 -290.240 -60.785 -290.015 ;
        RECT -63.065 -291.395 -62.835 -291.070 ;
        RECT -62.085 -291.395 -61.855 -291.070 ;
        RECT -64.045 -291.435 -61.855 -291.395 ;
        RECT -61.580 -291.315 -61.210 -290.475 ;
        RECT -60.960 -290.610 -60.790 -290.240 ;
        RECT -61.580 -291.435 -61.215 -291.315 ;
        RECT -65.065 -291.525 -64.225 -291.470 ;
        RECT -65.240 -291.530 -64.225 -291.525 ;
        RECT -69.285 -293.700 -69.045 -291.840 ;
        RECT -68.690 -292.805 -68.520 -292.010 ;
        RECT -68.230 -292.090 -68.000 -291.625 ;
        RECT -68.200 -292.550 -68.030 -292.090 ;
        RECT -67.710 -292.805 -67.540 -292.010 ;
        RECT -67.250 -292.090 -67.020 -291.625 ;
        RECT -66.270 -291.785 -65.605 -291.625 ;
        RECT -67.220 -292.550 -67.050 -292.090 ;
        RECT -66.730 -292.805 -66.560 -292.010 ;
        RECT -66.270 -292.090 -66.040 -291.785 ;
        RECT -65.425 -291.840 -64.225 -291.530 ;
        RECT -64.045 -291.625 -61.215 -291.435 ;
        RECT -66.240 -292.550 -66.070 -292.090 ;
        RECT -65.425 -292.560 -65.125 -291.840 ;
        RECT -64.505 -292.805 -64.335 -292.010 ;
        RECT -64.045 -292.090 -63.815 -291.625 ;
        RECT -64.015 -292.550 -63.845 -292.090 ;
        RECT -63.525 -292.805 -63.355 -292.010 ;
        RECT -63.065 -292.090 -62.835 -291.625 ;
        RECT -62.085 -291.785 -61.215 -291.625 ;
        RECT -60.990 -291.345 -60.755 -290.610 ;
        RECT -60.470 -290.645 -60.300 -290.185 ;
        RECT -59.985 -290.290 -59.775 -290.015 ;
        RECT -60.475 -290.905 -60.295 -290.645 ;
        RECT -59.980 -290.725 -59.810 -290.290 ;
        RECT -59.490 -290.635 -59.320 -290.185 ;
        RECT -59.015 -290.295 -58.805 -290.015 ;
        RECT -59.490 -290.725 -59.305 -290.635 ;
        RECT -59.000 -290.725 -58.830 -290.295 ;
        RECT -58.510 -290.635 -58.340 -290.185 ;
        RECT -58.035 -290.270 -57.825 -290.015 ;
        RECT -47.465 -290.015 -44.325 -289.845 ;
        RECT -54.700 -290.130 -54.530 -290.110 ;
        RECT -59.485 -290.905 -59.305 -290.725 ;
        RECT -58.515 -290.905 -58.335 -290.635 ;
        RECT -58.020 -290.725 -57.850 -290.270 ;
        RECT -57.530 -290.685 -57.360 -290.185 ;
        RECT -57.545 -290.905 -57.335 -290.685 ;
        RECT -60.475 -291.075 -57.335 -290.905 ;
        RECT -60.990 -291.715 -60.130 -291.345 ;
        RECT -58.210 -291.610 -57.335 -291.075 ;
        RECT -54.730 -291.395 -54.500 -290.130 ;
        RECT -53.720 -291.070 -53.550 -290.110 ;
        RECT -52.740 -291.070 -52.570 -290.110 ;
        RECT -50.515 -290.130 -50.345 -290.110 ;
        RECT -51.620 -290.480 -51.335 -290.220 ;
        RECT -52.360 -290.790 -51.335 -290.480 ;
        RECT -53.750 -291.395 -53.520 -291.070 ;
        RECT -52.770 -291.395 -52.540 -291.070 ;
        RECT -54.730 -291.435 -52.540 -291.395 ;
        RECT -52.360 -291.435 -52.050 -290.790 ;
        RECT -51.620 -291.040 -51.335 -290.790 ;
        RECT -55.750 -291.505 -54.910 -291.470 ;
        RECT -63.035 -292.550 -62.865 -292.090 ;
        RECT -62.545 -292.805 -62.375 -292.010 ;
        RECT -62.085 -292.090 -61.855 -291.785 ;
        RECT -62.055 -292.550 -61.885 -292.090 ;
        RECT -60.990 -292.390 -60.755 -291.715 ;
        RECT -58.210 -291.910 -56.880 -291.610 ;
        RECT -55.860 -291.805 -54.910 -291.505 ;
        RECT -55.750 -291.840 -54.910 -291.805 ;
        RECT -54.730 -291.625 -52.050 -291.435 ;
        RECT -50.545 -291.395 -50.315 -290.130 ;
        RECT -49.535 -291.070 -49.365 -290.110 ;
        RECT -48.555 -291.070 -48.385 -290.110 ;
        RECT -47.465 -290.240 -47.285 -290.015 ;
        RECT -49.565 -291.395 -49.335 -291.070 ;
        RECT -48.585 -291.395 -48.355 -291.070 ;
        RECT -50.545 -291.435 -48.355 -291.395 ;
        RECT -48.080 -291.315 -47.710 -290.475 ;
        RECT -47.460 -290.610 -47.290 -290.240 ;
        RECT -48.080 -291.435 -47.715 -291.315 ;
        RECT -51.565 -291.525 -50.725 -291.470 ;
        RECT -60.490 -292.080 -57.335 -291.910 ;
        RECT -60.490 -292.285 -60.285 -292.080 ;
        RECT -60.960 -292.740 -60.790 -292.390 ;
        RECT -68.735 -293.145 -61.880 -292.805 ;
        RECT -60.985 -293.030 -60.765 -292.740 ;
        RECT -60.470 -292.800 -60.300 -292.285 ;
        RECT -59.980 -292.685 -59.810 -292.260 ;
        RECT -59.500 -292.325 -59.295 -292.080 ;
        RECT -60.005 -293.030 -59.785 -292.685 ;
        RECT -59.490 -292.800 -59.320 -292.325 ;
        RECT -59.000 -292.685 -58.830 -292.260 ;
        RECT -58.530 -292.325 -58.325 -292.080 ;
        RECT -57.545 -292.115 -57.335 -292.080 ;
        RECT -59.025 -293.030 -58.805 -292.685 ;
        RECT -58.510 -292.800 -58.340 -292.325 ;
        RECT -58.020 -292.740 -57.850 -292.260 ;
        RECT -57.545 -292.330 -57.340 -292.115 ;
        RECT -58.040 -293.030 -57.820 -292.740 ;
        RECT -57.530 -292.800 -57.360 -292.330 ;
        RECT -55.190 -292.805 -55.020 -292.010 ;
        RECT -54.730 -292.090 -54.500 -291.625 ;
        RECT -54.700 -292.550 -54.530 -292.090 ;
        RECT -54.210 -292.805 -54.040 -292.010 ;
        RECT -53.750 -292.090 -53.520 -291.625 ;
        RECT -52.770 -291.785 -52.050 -291.625 ;
        RECT -53.720 -292.550 -53.550 -292.090 ;
        RECT -53.230 -292.805 -53.060 -292.010 ;
        RECT -52.770 -292.090 -52.540 -291.785 ;
        RECT -51.865 -291.840 -50.725 -291.525 ;
        RECT -50.545 -291.625 -47.715 -291.435 ;
        RECT -52.740 -292.550 -52.570 -292.090 ;
        RECT -51.865 -292.635 -51.565 -291.840 ;
        RECT -51.005 -292.805 -50.835 -292.010 ;
        RECT -50.545 -292.090 -50.315 -291.625 ;
        RECT -50.515 -292.550 -50.345 -292.090 ;
        RECT -50.025 -292.805 -49.855 -292.010 ;
        RECT -49.565 -292.090 -49.335 -291.625 ;
        RECT -48.585 -291.785 -47.715 -291.625 ;
        RECT -47.490 -291.345 -47.255 -290.610 ;
        RECT -46.970 -290.645 -46.800 -290.185 ;
        RECT -46.485 -290.290 -46.275 -290.015 ;
        RECT -46.975 -290.905 -46.795 -290.645 ;
        RECT -46.480 -290.725 -46.310 -290.290 ;
        RECT -45.990 -290.635 -45.820 -290.185 ;
        RECT -45.515 -290.295 -45.305 -290.015 ;
        RECT -45.990 -290.725 -45.805 -290.635 ;
        RECT -45.500 -290.725 -45.330 -290.295 ;
        RECT -45.010 -290.635 -44.840 -290.185 ;
        RECT -44.535 -290.270 -44.325 -290.015 ;
        RECT -36.205 -290.025 -35.005 -289.855 ;
        RECT -45.985 -290.905 -45.805 -290.725 ;
        RECT -45.015 -290.905 -44.835 -290.635 ;
        RECT -44.520 -290.725 -44.350 -290.270 ;
        RECT -44.030 -290.685 -43.860 -290.185 ;
        RECT -44.045 -290.905 -43.835 -290.685 ;
        RECT -46.975 -291.075 -43.835 -290.905 ;
        RECT -47.490 -291.715 -46.630 -291.345 ;
        RECT -44.710 -291.620 -43.835 -291.075 ;
        RECT -49.535 -292.550 -49.365 -292.090 ;
        RECT -49.045 -292.805 -48.875 -292.010 ;
        RECT -48.585 -292.090 -48.355 -291.785 ;
        RECT -48.555 -292.550 -48.385 -292.090 ;
        RECT -47.490 -292.390 -47.255 -291.715 ;
        RECT -44.710 -291.910 -43.460 -291.620 ;
        RECT -46.990 -291.920 -43.460 -291.910 ;
        RECT -46.990 -292.080 -43.835 -291.920 ;
        RECT -46.990 -292.285 -46.785 -292.080 ;
        RECT -47.460 -292.740 -47.290 -292.390 ;
        RECT -67.495 -293.345 -66.940 -293.145 ;
        RECT -67.550 -293.385 -66.865 -293.345 ;
        RECT -63.440 -293.385 -62.885 -293.145 ;
        RECT -60.985 -293.200 -57.820 -293.030 ;
        RECT -55.235 -292.815 -52.565 -292.805 ;
        RECT -51.050 -292.815 -48.380 -292.805 ;
        RECT -55.235 -293.145 -48.380 -292.815 ;
        RECT -47.485 -293.030 -47.265 -292.740 ;
        RECT -46.970 -292.800 -46.800 -292.285 ;
        RECT -46.480 -292.685 -46.310 -292.260 ;
        RECT -46.000 -292.325 -45.795 -292.080 ;
        RECT -46.505 -293.030 -46.285 -292.685 ;
        RECT -45.990 -292.800 -45.820 -292.325 ;
        RECT -45.500 -292.685 -45.330 -292.260 ;
        RECT -45.030 -292.325 -44.825 -292.080 ;
        RECT -44.045 -292.115 -43.835 -292.080 ;
        RECT -45.525 -293.030 -45.305 -292.685 ;
        RECT -45.010 -292.800 -44.840 -292.325 ;
        RECT -44.520 -292.740 -44.350 -292.260 ;
        RECT -44.045 -292.330 -43.840 -292.115 ;
        RECT -44.540 -293.030 -44.320 -292.740 ;
        RECT -44.030 -292.800 -43.860 -292.330 ;
        RECT -54.450 -293.375 -53.895 -293.145 ;
        RECT -53.535 -293.155 -50.935 -293.145 ;
        RECT -54.565 -293.385 -53.880 -293.375 ;
        RECT -50.060 -293.385 -49.505 -293.145 ;
        RECT -47.485 -293.200 -44.320 -293.030 ;
        RECT -37.235 -293.165 -37.065 -290.195 ;
        RECT -36.205 -290.245 -35.995 -290.025 ;
        RECT -41.375 -293.385 -40.715 -293.375 ;
        RECT -67.635 -293.580 -40.710 -293.385 ;
        RECT -67.550 -293.645 -66.865 -293.580 ;
        RECT -54.565 -293.675 -53.880 -293.580 ;
        RECT -41.375 -293.675 -40.715 -293.580 ;
        RECT -69.290 -294.385 -68.990 -293.700 ;
        RECT -56.740 -293.845 -56.055 -293.790 ;
        RECT -52.010 -293.845 -51.350 -293.795 ;
        RECT -67.635 -294.040 -38.985 -293.845 ;
        RECT -56.740 -294.090 -56.055 -294.040 ;
        RECT -52.010 -294.095 -51.350 -294.040 ;
        RECT -65.605 -294.275 -64.945 -294.235 ;
        RECT -42.990 -294.275 -42.330 -294.225 ;
        RECT -98.535 -295.000 -97.315 -294.810 ;
        RECT -104.085 -295.355 -101.770 -295.185 ;
        RECT -105.585 -298.490 -105.415 -295.535 ;
        RECT -105.605 -298.745 -105.400 -298.490 ;
        RECT -104.525 -298.525 -104.355 -295.535 ;
        RECT -104.085 -295.565 -103.820 -295.355 ;
        RECT -104.550 -298.745 -104.340 -298.525 ;
        RECT -104.035 -298.575 -103.865 -295.565 ;
        RECT -103.545 -298.520 -103.375 -295.535 ;
        RECT -103.040 -295.565 -102.760 -295.355 ;
        RECT -103.570 -298.745 -103.360 -298.520 ;
        RECT -102.980 -298.575 -102.810 -295.565 ;
        RECT -102.490 -298.485 -102.320 -295.535 ;
        RECT -102.050 -295.565 -101.770 -295.355 ;
        RECT -105.605 -298.930 -103.360 -298.745 ;
        RECT -102.510 -298.765 -102.300 -298.485 ;
        RECT -102.000 -298.575 -101.830 -295.565 ;
        RECT -99.555 -297.195 -99.385 -295.180 ;
        RECT -98.535 -295.320 -98.305 -295.000 ;
        RECT -99.560 -297.390 -99.380 -297.195 ;
        RECT -98.500 -297.220 -98.330 -295.320 ;
        RECT -98.010 -297.170 -97.840 -295.180 ;
        RECT -97.545 -295.320 -97.315 -295.000 ;
        RECT -94.010 -295.005 -92.790 -294.815 ;
        RECT -97.520 -296.990 -97.350 -295.320 ;
        RECT -98.045 -297.390 -97.820 -297.170 ;
        RECT -99.560 -297.570 -97.820 -297.390 ;
        RECT -97.535 -298.150 -97.285 -296.990 ;
        RECT -95.030 -297.200 -94.860 -295.185 ;
        RECT -94.010 -295.325 -93.780 -295.005 ;
        RECT -96.365 -297.805 -96.075 -297.330 ;
        RECT -95.035 -297.395 -94.855 -297.200 ;
        RECT -93.975 -297.225 -93.805 -295.325 ;
        RECT -93.485 -297.175 -93.315 -295.185 ;
        RECT -93.020 -295.325 -92.790 -295.005 ;
        RECT -84.455 -295.195 -77.070 -294.630 ;
        RECT -92.995 -296.995 -92.825 -295.325 ;
        RECT -88.610 -296.670 -86.365 -296.580 ;
        RECT -84.455 -296.670 -84.150 -295.195 ;
        RECT -80.820 -295.785 -80.585 -295.195 ;
        RECT -91.170 -296.975 -84.150 -296.670 ;
        RECT -93.520 -297.395 -93.295 -297.175 ;
        RECT -95.035 -297.575 -93.295 -297.395 ;
        RECT -94.385 -297.805 -93.670 -297.770 ;
        RECT -96.365 -297.985 -93.670 -297.805 ;
        RECT -96.365 -298.015 -96.075 -297.985 ;
        RECT -94.385 -298.070 -93.670 -297.985 ;
        RECT -100.570 -298.245 -100.280 -298.180 ;
        RECT -100.025 -298.245 -99.295 -298.165 ;
        RECT -97.535 -298.215 -96.805 -298.150 ;
        RECT -93.010 -298.155 -92.760 -296.995 ;
        RECT -100.570 -298.425 -99.295 -298.245 ;
        RECT -97.815 -298.260 -96.805 -298.215 ;
        RECT -102.510 -298.975 -101.670 -298.765 ;
        RECT -100.570 -298.865 -100.280 -298.425 ;
        RECT -100.025 -298.465 -99.295 -298.425 ;
        RECT -99.090 -298.440 -96.805 -298.260 ;
        RECT -95.980 -298.250 -95.690 -298.190 ;
        RECT -95.500 -298.250 -94.770 -298.170 ;
        RECT -93.010 -298.220 -92.150 -298.155 ;
        RECT -95.980 -298.430 -94.770 -298.250 ;
        RECT -93.290 -298.265 -92.150 -298.220 ;
        RECT -101.880 -299.895 -101.670 -298.975 ;
        RECT -99.555 -299.435 -99.385 -298.640 ;
        RECT -99.090 -298.685 -98.865 -298.440 ;
        RECT -101.925 -299.975 -101.240 -299.895 ;
        RECT -105.115 -300.185 -101.240 -299.975 ;
        RECT -105.585 -301.210 -105.415 -300.355 ;
        RECT -105.115 -300.440 -104.905 -300.185 ;
        RECT -105.610 -301.855 -105.370 -301.210 ;
        RECT -105.095 -301.395 -104.925 -300.440 ;
        RECT -104.605 -301.195 -104.435 -300.355 ;
        RECT -104.135 -300.440 -103.925 -300.185 ;
        RECT -99.575 -300.195 -99.355 -299.435 ;
        RECT -99.065 -299.680 -98.895 -298.685 ;
        RECT -98.575 -299.440 -98.405 -298.640 ;
        RECT -95.980 -298.875 -95.690 -298.430 ;
        RECT -95.500 -298.470 -94.770 -298.430 ;
        RECT -94.565 -298.445 -92.150 -298.265 ;
        RECT -95.030 -299.440 -94.860 -298.645 ;
        RECT -94.565 -298.690 -94.340 -298.445 ;
        RECT -98.605 -300.195 -98.385 -299.440 ;
        RECT -100.220 -300.370 -97.235 -300.195 ;
        RECT -95.050 -300.200 -94.830 -299.440 ;
        RECT -94.540 -299.685 -94.370 -298.690 ;
        RECT -94.050 -299.445 -93.880 -298.645 ;
        RECT -91.170 -298.765 -90.865 -296.975 ;
        RECT -88.025 -297.145 -87.850 -296.975 ;
        RECT -88.510 -298.685 -88.340 -297.145 ;
        RECT -88.020 -298.685 -87.850 -297.145 ;
        RECT -87.530 -298.685 -87.360 -297.145 ;
        RECT -87.040 -298.685 -86.870 -297.145 ;
        RECT -86.550 -298.685 -86.380 -297.145 ;
        RECT -93.105 -299.070 -90.865 -298.765 ;
        RECT -88.670 -298.900 -88.315 -298.895 ;
        RECT -86.610 -298.900 -86.240 -298.870 ;
        RECT -88.670 -298.905 -86.240 -298.900 ;
        RECT -94.080 -300.200 -93.860 -299.445 ;
        RECT -93.105 -300.200 -92.800 -299.070 ;
        RECT -89.800 -299.095 -86.240 -298.905 ;
        RECT -84.455 -299.010 -84.150 -296.975 ;
        RECT -80.785 -297.255 -80.615 -295.785 ;
        RECT -80.295 -297.175 -80.125 -295.715 ;
        RECT -79.840 -295.790 -79.605 -295.195 ;
        RECT -81.330 -297.485 -80.555 -297.425 ;
        RECT -81.515 -297.655 -80.555 -297.485 ;
        RECT -81.330 -297.700 -80.555 -297.655 ;
        RECT -80.325 -297.525 -80.100 -297.175 ;
        RECT -79.805 -297.255 -79.635 -295.790 ;
        RECT -78.630 -295.840 -78.395 -295.195 ;
        RECT -78.595 -297.255 -78.425 -295.840 ;
        RECT -78.105 -297.210 -77.935 -295.715 ;
        RECT -69.285 -296.175 -69.045 -294.385 ;
        RECT -67.635 -294.470 -42.330 -294.275 ;
        RECT -65.605 -294.535 -64.945 -294.470 ;
        RECT -42.990 -294.525 -42.330 -294.470 ;
        RECT -39.180 -294.385 -38.985 -294.040 ;
        RECT -37.275 -294.385 -37.060 -293.165 ;
        RECT -36.175 -293.235 -36.005 -290.245 ;
        RECT -35.685 -293.135 -35.515 -290.195 ;
        RECT -35.215 -290.235 -35.005 -290.025 ;
        RECT -35.705 -293.405 -35.495 -293.135 ;
        RECT -35.195 -293.145 -35.025 -290.235 ;
        RECT -34.140 -293.115 -33.970 -290.195 ;
        RECT -3.270 -290.515 -1.780 -286.225 ;
        RECT 4.775 -290.515 6.080 -286.225 ;
        RECT 8.960 -290.515 10.265 -286.225 ;
        RECT 14.160 -290.515 15.465 -286.225 ;
        RECT 21.450 -290.515 22.755 -286.225 ;
        RECT 27.520 -290.515 28.825 -286.225 ;
        RECT 37.250 -290.515 38.555 -286.225 ;
        RECT 44.720 -290.515 46.025 -286.225 ;
        RECT 95.890 -286.220 96.155 -286.010 ;
        RECT 96.430 -286.040 96.600 -283.055 ;
        RECT 96.995 -286.010 97.165 -283.000 ;
        RECT 97.465 -283.090 97.675 -282.810 ;
        RECT 96.935 -286.220 97.215 -286.010 ;
        RECT 97.485 -286.040 97.655 -283.090 ;
        RECT 97.975 -286.010 98.145 -283.000 ;
        RECT 97.925 -286.220 98.205 -286.010 ;
        RECT 95.890 -286.390 98.205 -286.220 ;
        RECT -21.595 -291.350 -18.455 -291.180 ;
        RECT -28.830 -291.465 -28.660 -291.445 ;
        RECT -28.860 -292.730 -28.630 -291.465 ;
        RECT -27.850 -292.405 -27.680 -291.445 ;
        RECT -26.870 -292.405 -26.700 -291.445 ;
        RECT -24.645 -291.465 -24.475 -291.445 ;
        RECT -25.750 -291.875 -25.465 -291.555 ;
        RECT -26.465 -292.120 -25.465 -291.875 ;
        RECT -27.880 -292.730 -27.650 -292.405 ;
        RECT -26.900 -292.730 -26.670 -292.405 ;
        RECT -28.860 -292.770 -26.670 -292.730 ;
        RECT -26.465 -292.770 -26.235 -292.120 ;
        RECT -25.750 -292.375 -25.465 -292.120 ;
        RECT -29.880 -292.955 -29.040 -292.805 ;
        RECT -36.200 -293.600 -35.495 -293.405 ;
        RECT -35.220 -293.410 -35.010 -293.145 ;
        RECT -34.160 -293.410 -33.950 -293.115 ;
        RECT -35.220 -293.590 -33.950 -293.410 ;
        RECT -29.915 -293.175 -29.040 -292.955 ;
        RECT -28.860 -292.960 -26.235 -292.770 ;
        RECT -24.675 -292.730 -24.445 -291.465 ;
        RECT -23.665 -292.405 -23.495 -291.445 ;
        RECT -22.685 -292.405 -22.515 -291.445 ;
        RECT -21.595 -291.575 -21.415 -291.350 ;
        RECT -23.695 -292.730 -23.465 -292.405 ;
        RECT -22.715 -292.730 -22.485 -292.405 ;
        RECT -24.675 -292.770 -22.485 -292.730 ;
        RECT -22.210 -292.650 -21.840 -291.810 ;
        RECT -21.590 -291.945 -21.420 -291.575 ;
        RECT -22.210 -292.770 -21.845 -292.650 ;
        RECT -25.695 -292.860 -24.855 -292.805 ;
        RECT -25.870 -292.865 -24.855 -292.860 ;
        RECT -36.200 -293.660 -35.985 -293.600 ;
        RECT -36.890 -293.935 -35.985 -293.660 ;
        RECT -36.200 -294.285 -35.985 -293.935 ;
        RECT -35.550 -293.820 -34.775 -293.770 ;
        RECT -32.985 -293.820 -32.325 -293.560 ;
        RECT -35.550 -294.000 -32.325 -293.820 ;
        RECT -35.550 -294.045 -34.775 -294.000 ;
        RECT -39.180 -294.585 -36.390 -294.385 ;
        RECT -36.200 -294.485 -34.430 -294.285 ;
        RECT -39.180 -294.600 -36.630 -294.585 ;
        RECT -68.695 -295.045 -66.025 -294.705 ;
        RECT -64.040 -294.820 -60.875 -294.650 ;
        RECT -68.690 -295.760 -68.520 -295.300 ;
        RECT -68.720 -296.065 -68.490 -295.760 ;
        RECT -68.200 -295.840 -68.030 -295.045 ;
        RECT -67.710 -295.760 -67.540 -295.300 ;
        RECT -68.870 -296.175 -68.490 -296.065 ;
        RECT -69.285 -296.225 -68.490 -296.175 ;
        RECT -67.740 -296.225 -67.510 -295.760 ;
        RECT -67.220 -295.840 -67.050 -295.045 ;
        RECT -66.730 -295.760 -66.560 -295.300 ;
        RECT -66.760 -296.225 -66.530 -295.760 ;
        RECT -66.240 -295.840 -66.070 -295.045 ;
        RECT -64.500 -295.520 -64.330 -295.050 ;
        RECT -64.040 -295.110 -63.820 -294.820 ;
        RECT -64.520 -295.735 -64.315 -295.520 ;
        RECT -64.010 -295.590 -63.840 -295.110 ;
        RECT -63.520 -295.525 -63.350 -295.050 ;
        RECT -63.055 -295.165 -62.835 -294.820 ;
        RECT -64.525 -295.770 -64.315 -295.735 ;
        RECT -63.535 -295.770 -63.330 -295.525 ;
        RECT -63.030 -295.590 -62.860 -295.165 ;
        RECT -62.540 -295.525 -62.370 -295.050 ;
        RECT -62.075 -295.165 -61.855 -294.820 ;
        RECT -62.565 -295.770 -62.360 -295.525 ;
        RECT -62.050 -295.590 -61.880 -295.165 ;
        RECT -61.560 -295.565 -61.390 -295.050 ;
        RECT -61.095 -295.110 -60.875 -294.820 ;
        RECT -59.980 -295.045 -52.525 -294.705 ;
        RECT -50.540 -294.820 -47.375 -294.650 ;
        RECT -61.070 -295.460 -60.900 -295.110 ;
        RECT -61.575 -295.770 -61.370 -295.565 ;
        RECT -64.525 -295.940 -61.370 -295.770 ;
        RECT -69.285 -296.360 -66.530 -296.225 ;
        RECT -69.280 -296.370 -66.530 -296.360 ;
        RECT -68.870 -296.415 -66.530 -296.370 ;
        RECT -66.350 -296.085 -65.510 -296.010 ;
        RECT -64.525 -296.085 -63.650 -295.940 ;
        RECT -66.350 -296.350 -63.650 -296.085 ;
        RECT -61.105 -296.135 -60.870 -295.460 ;
        RECT -59.975 -295.760 -59.805 -295.300 ;
        RECT -60.005 -296.065 -59.775 -295.760 ;
        RECT -59.485 -295.840 -59.315 -295.045 ;
        RECT -58.995 -295.760 -58.825 -295.300 ;
        RECT -66.350 -296.380 -65.510 -296.350 ;
        RECT -68.720 -296.455 -66.530 -296.415 ;
        RECT -68.720 -296.780 -68.490 -296.455 ;
        RECT -67.740 -296.780 -67.510 -296.455 ;
        RECT -78.125 -297.410 -77.905 -297.210 ;
        RECT -73.665 -297.410 -72.980 -297.060 ;
        RECT -78.125 -297.425 -72.980 -297.410 ;
        RECT -80.325 -297.725 -78.555 -297.525 ;
        RECT -78.365 -297.625 -72.980 -297.425 ;
        RECT -82.005 -298.010 -81.655 -298.000 ;
        RECT -79.980 -298.010 -79.205 -297.965 ;
        RECT -82.005 -298.190 -79.205 -298.010 ;
        RECT -89.800 -299.105 -88.665 -299.095 ;
        RECT -86.610 -299.225 -86.240 -299.095 ;
        RECT -91.530 -299.395 -90.945 -299.320 ;
        RECT -88.935 -299.385 -88.260 -299.345 ;
        RECT -89.035 -299.395 -88.260 -299.385 ;
        RECT -91.530 -299.575 -88.260 -299.395 ;
        RECT -85.675 -299.440 -82.600 -299.010 ;
        RECT -91.530 -299.935 -90.945 -299.575 ;
        RECT -89.035 -299.585 -88.260 -299.575 ;
        RECT -88.935 -299.615 -88.260 -299.585 ;
        RECT -88.020 -299.500 -85.925 -299.460 ;
        RECT -88.020 -299.650 -85.870 -299.500 ;
        RECT -95.695 -300.370 -92.710 -300.200 ;
        RECT -104.640 -301.855 -104.400 -301.195 ;
        RECT -104.115 -301.395 -103.945 -300.440 ;
        RECT -102.995 -300.645 -92.710 -300.370 ;
        RECT -102.995 -300.950 -93.790 -300.645 ;
        RECT -102.995 -301.855 -102.415 -300.950 ;
        RECT -88.020 -301.370 -87.850 -299.650 ;
        RECT -87.040 -301.370 -86.870 -299.650 ;
        RECT -86.175 -300.395 -85.870 -299.650 ;
        RECT -84.975 -300.220 -84.805 -299.440 ;
        RECT -84.485 -300.220 -84.315 -299.680 ;
        RECT -83.995 -300.220 -83.825 -299.440 ;
        RECT -83.505 -300.220 -83.335 -299.680 ;
        RECT -82.005 -300.165 -81.655 -298.190 ;
        RECT -79.980 -298.240 -79.205 -298.190 ;
        RECT -78.770 -298.075 -78.555 -297.725 ;
        RECT -78.770 -298.350 -77.865 -298.075 ;
        RECT -78.770 -298.410 -78.555 -298.350 ;
        RECT -80.805 -298.600 -79.535 -298.420 ;
        RECT -80.805 -298.895 -80.595 -298.600 ;
        RECT -79.745 -298.865 -79.535 -298.600 ;
        RECT -79.260 -298.605 -78.555 -298.410 ;
        RECT -85.565 -300.395 -85.200 -300.365 ;
        RECT -86.175 -300.460 -85.200 -300.395 ;
        RECT -86.065 -300.600 -85.200 -300.460 ;
        RECT -85.565 -300.665 -85.200 -300.600 ;
        RECT -83.015 -300.515 -81.625 -300.165 ;
        RECT -84.975 -301.375 -84.805 -300.835 ;
        RECT -83.995 -301.375 -83.825 -300.835 ;
        RECT -83.015 -301.375 -82.845 -300.515 ;
        RECT -80.785 -301.815 -80.615 -298.895 ;
        RECT -79.730 -301.775 -79.560 -298.865 ;
        RECT -79.260 -298.875 -79.050 -298.605 ;
        RECT -106.285 -301.940 -102.265 -301.855 ;
        RECT -106.285 -302.470 -101.845 -301.940 ;
        RECT -79.750 -301.985 -79.540 -301.775 ;
        RECT -79.240 -301.815 -79.070 -298.875 ;
        RECT -78.750 -301.765 -78.580 -298.775 ;
        RECT -77.695 -298.845 -77.480 -297.625 ;
        RECT -73.665 -297.890 -72.980 -297.625 ;
        RECT -68.690 -297.740 -68.520 -296.780 ;
        RECT -67.710 -297.740 -67.540 -296.780 ;
        RECT -66.760 -297.720 -66.530 -296.455 ;
        RECT -64.525 -296.775 -63.650 -296.350 ;
        RECT -61.730 -296.505 -60.870 -296.135 ;
        RECT -64.525 -296.945 -61.385 -296.775 ;
        RECT -64.525 -297.165 -64.315 -296.945 ;
        RECT -64.500 -297.665 -64.330 -297.165 ;
        RECT -64.010 -297.580 -63.840 -297.125 ;
        RECT -63.525 -297.215 -63.345 -296.945 ;
        RECT -62.555 -297.125 -62.375 -296.945 ;
        RECT -66.730 -297.740 -66.560 -297.720 ;
        RECT -64.035 -297.835 -63.825 -297.580 ;
        RECT -63.520 -297.665 -63.350 -297.215 ;
        RECT -63.030 -297.555 -62.860 -297.125 ;
        RECT -62.555 -297.215 -62.370 -297.125 ;
        RECT -63.055 -297.835 -62.845 -297.555 ;
        RECT -62.540 -297.665 -62.370 -297.215 ;
        RECT -62.050 -297.560 -61.880 -297.125 ;
        RECT -61.565 -297.205 -61.385 -296.945 ;
        RECT -62.085 -297.835 -61.875 -297.560 ;
        RECT -61.560 -297.665 -61.390 -297.205 ;
        RECT -61.105 -297.240 -60.870 -296.505 ;
        RECT -60.645 -296.225 -59.775 -296.065 ;
        RECT -59.025 -296.225 -58.795 -295.760 ;
        RECT -58.505 -295.840 -58.335 -295.045 ;
        RECT -58.015 -295.760 -57.845 -295.300 ;
        RECT -58.045 -296.225 -57.815 -295.760 ;
        RECT -57.525 -295.840 -57.355 -295.045 ;
        RECT -60.645 -296.415 -57.815 -296.225 ;
        RECT -57.635 -296.035 -56.795 -296.010 ;
        RECT -56.495 -296.035 -56.195 -295.670 ;
        RECT -57.635 -296.325 -56.195 -296.035 ;
        RECT -55.920 -296.120 -55.620 -295.545 ;
        RECT -55.190 -295.760 -55.020 -295.300 ;
        RECT -55.220 -296.065 -54.990 -295.760 ;
        RECT -54.700 -295.840 -54.530 -295.045 ;
        RECT -54.210 -295.760 -54.040 -295.300 ;
        RECT -55.370 -296.120 -54.990 -296.065 ;
        RECT -57.635 -296.380 -56.795 -296.325 ;
        RECT -56.495 -296.330 -56.195 -296.325 ;
        RECT -55.945 -296.225 -54.990 -296.120 ;
        RECT -54.240 -296.225 -54.010 -295.760 ;
        RECT -53.720 -295.840 -53.550 -295.045 ;
        RECT -53.230 -295.760 -53.060 -295.300 ;
        RECT -53.260 -296.225 -53.030 -295.760 ;
        RECT -52.740 -295.840 -52.570 -295.045 ;
        RECT -51.015 -295.520 -50.785 -294.910 ;
        RECT -50.540 -295.110 -50.320 -294.820 ;
        RECT -51.020 -295.570 -50.785 -295.520 ;
        RECT -51.020 -295.735 -50.815 -295.570 ;
        RECT -50.510 -295.590 -50.340 -295.110 ;
        RECT -50.020 -295.525 -49.850 -295.050 ;
        RECT -49.555 -295.165 -49.335 -294.820 ;
        RECT -51.025 -295.770 -50.815 -295.735 ;
        RECT -50.035 -295.770 -49.830 -295.525 ;
        RECT -49.530 -295.590 -49.360 -295.165 ;
        RECT -49.040 -295.525 -48.870 -295.050 ;
        RECT -48.575 -295.165 -48.355 -294.820 ;
        RECT -49.065 -295.770 -48.860 -295.525 ;
        RECT -48.550 -295.590 -48.380 -295.165 ;
        RECT -48.060 -295.565 -47.890 -295.050 ;
        RECT -47.595 -295.110 -47.375 -294.820 ;
        RECT -46.480 -295.045 -39.400 -294.705 ;
        RECT -47.570 -295.460 -47.400 -295.110 ;
        RECT -48.075 -295.770 -47.870 -295.565 ;
        RECT -51.025 -295.940 -47.870 -295.770 ;
        RECT -55.945 -296.345 -53.030 -296.225 ;
        RECT -60.645 -296.535 -60.280 -296.415 ;
        RECT -61.070 -297.610 -60.900 -297.240 ;
        RECT -60.650 -297.375 -60.280 -296.535 ;
        RECT -60.005 -296.455 -57.815 -296.415 ;
        RECT -60.005 -296.780 -59.775 -296.455 ;
        RECT -59.025 -296.780 -58.795 -296.455 ;
        RECT -61.075 -297.835 -60.895 -297.610 ;
        RECT -59.975 -297.740 -59.805 -296.780 ;
        RECT -58.995 -297.740 -58.825 -296.780 ;
        RECT -58.045 -297.720 -57.815 -296.455 ;
        RECT -57.025 -297.015 -56.740 -296.810 ;
        RECT -55.945 -297.015 -55.720 -296.345 ;
        RECT -55.370 -296.415 -53.030 -296.345 ;
        RECT -52.850 -296.050 -52.010 -296.010 ;
        RECT -51.025 -296.050 -50.150 -295.940 ;
        RECT -52.850 -296.335 -50.150 -296.050 ;
        RECT -47.605 -296.135 -47.370 -295.460 ;
        RECT -46.475 -295.760 -46.305 -295.300 ;
        RECT -46.505 -296.065 -46.275 -295.760 ;
        RECT -45.985 -295.840 -45.815 -295.045 ;
        RECT -45.495 -295.760 -45.325 -295.300 ;
        RECT -52.850 -296.380 -52.010 -296.335 ;
        RECT -55.220 -296.455 -53.030 -296.415 ;
        RECT -55.220 -296.780 -54.990 -296.455 ;
        RECT -54.240 -296.780 -54.010 -296.455 ;
        RECT -57.025 -297.240 -55.720 -297.015 ;
        RECT -57.025 -297.630 -56.740 -297.240 ;
        RECT -58.015 -297.740 -57.845 -297.720 ;
        RECT -55.190 -297.740 -55.020 -296.780 ;
        RECT -54.210 -297.740 -54.040 -296.780 ;
        RECT -53.260 -297.720 -53.030 -296.455 ;
        RECT -51.025 -296.775 -50.150 -296.335 ;
        RECT -48.230 -296.505 -47.370 -296.135 ;
        RECT -51.025 -296.945 -47.885 -296.775 ;
        RECT -51.025 -297.165 -50.815 -296.945 ;
        RECT -51.000 -297.665 -50.830 -297.165 ;
        RECT -50.510 -297.580 -50.340 -297.125 ;
        RECT -50.025 -297.215 -49.845 -296.945 ;
        RECT -49.055 -297.125 -48.875 -296.945 ;
        RECT -53.230 -297.740 -53.060 -297.720 ;
        RECT -64.035 -298.005 -60.895 -297.835 ;
        RECT -50.535 -297.835 -50.325 -297.580 ;
        RECT -50.020 -297.665 -49.850 -297.215 ;
        RECT -49.530 -297.555 -49.360 -297.125 ;
        RECT -49.055 -297.215 -48.870 -297.125 ;
        RECT -49.555 -297.835 -49.345 -297.555 ;
        RECT -49.040 -297.665 -48.870 -297.215 ;
        RECT -48.550 -297.560 -48.380 -297.125 ;
        RECT -48.065 -297.205 -47.885 -296.945 ;
        RECT -48.585 -297.835 -48.375 -297.560 ;
        RECT -48.060 -297.665 -47.890 -297.205 ;
        RECT -47.605 -297.240 -47.370 -296.505 ;
        RECT -47.145 -296.225 -46.275 -296.065 ;
        RECT -45.525 -296.225 -45.295 -295.760 ;
        RECT -45.005 -295.840 -44.835 -295.045 ;
        RECT -44.515 -295.760 -44.345 -295.300 ;
        RECT -44.545 -296.225 -44.315 -295.760 ;
        RECT -44.025 -295.840 -43.855 -295.045 ;
        RECT -47.145 -296.415 -44.315 -296.225 ;
        RECT -44.135 -296.035 -43.295 -296.010 ;
        RECT -44.135 -296.095 -43.120 -296.035 ;
        RECT -42.835 -296.095 -42.535 -295.665 ;
        RECT -42.065 -295.760 -41.895 -295.300 ;
        RECT -42.095 -296.065 -41.865 -295.760 ;
        RECT -41.575 -295.840 -41.405 -295.045 ;
        RECT -41.085 -295.760 -40.915 -295.300 ;
        RECT -42.245 -296.095 -41.865 -296.065 ;
        RECT -44.135 -296.225 -41.865 -296.095 ;
        RECT -41.115 -296.225 -40.885 -295.760 ;
        RECT -40.595 -295.840 -40.425 -295.045 ;
        RECT -40.105 -295.760 -39.935 -295.300 ;
        RECT -40.135 -296.225 -39.905 -295.760 ;
        RECT -39.615 -295.840 -39.445 -295.045 ;
        RECT -39.180 -296.010 -38.985 -294.600 ;
        RECT -36.850 -294.800 -36.630 -294.600 ;
        RECT -44.135 -296.305 -39.905 -296.225 ;
        RECT -44.135 -296.325 -43.120 -296.305 ;
        RECT -42.835 -296.325 -42.535 -296.305 ;
        RECT -44.135 -296.380 -43.295 -296.325 ;
        RECT -42.245 -296.415 -39.905 -296.305 ;
        RECT -39.725 -296.380 -38.885 -296.010 ;
        RECT -36.820 -296.295 -36.650 -294.800 ;
        RECT -36.330 -296.170 -36.160 -294.755 ;
        RECT -47.145 -296.535 -46.780 -296.415 ;
        RECT -47.570 -297.610 -47.400 -297.240 ;
        RECT -47.150 -297.375 -46.780 -296.535 ;
        RECT -46.505 -296.455 -44.315 -296.415 ;
        RECT -46.505 -296.780 -46.275 -296.455 ;
        RECT -45.525 -296.780 -45.295 -296.455 ;
        RECT -47.575 -297.835 -47.395 -297.610 ;
        RECT -46.475 -297.740 -46.305 -296.780 ;
        RECT -45.495 -297.740 -45.325 -296.780 ;
        RECT -44.545 -297.720 -44.315 -296.455 ;
        RECT -42.095 -296.455 -39.905 -296.415 ;
        RECT -42.095 -296.780 -41.865 -296.455 ;
        RECT -41.115 -296.780 -40.885 -296.455 ;
        RECT -43.525 -297.630 -43.240 -296.810 ;
        RECT -44.515 -297.740 -44.345 -297.720 ;
        RECT -42.065 -297.740 -41.895 -296.780 ;
        RECT -41.085 -297.740 -40.915 -296.780 ;
        RECT -40.135 -297.720 -39.905 -296.455 ;
        RECT -36.360 -296.820 -36.125 -296.170 ;
        RECT -35.120 -296.220 -34.950 -294.755 ;
        RECT -34.655 -294.835 -34.430 -294.485 ;
        RECT -34.200 -294.355 -33.425 -294.310 ;
        RECT -31.610 -294.355 -30.900 -294.270 ;
        RECT -34.200 -294.525 -30.900 -294.355 ;
        RECT -34.200 -294.585 -33.425 -294.525 ;
        RECT -31.610 -294.590 -30.900 -294.525 ;
        RECT -35.150 -296.820 -34.915 -296.220 ;
        RECT -34.630 -296.295 -34.460 -294.835 ;
        RECT -34.140 -296.225 -33.970 -294.755 ;
        RECT -29.915 -295.035 -29.675 -293.175 ;
        RECT -29.320 -294.140 -29.150 -293.345 ;
        RECT -28.860 -293.425 -28.630 -292.960 ;
        RECT -28.830 -293.885 -28.660 -293.425 ;
        RECT -28.340 -294.140 -28.170 -293.345 ;
        RECT -27.880 -293.425 -27.650 -292.960 ;
        RECT -26.900 -293.120 -26.235 -292.960 ;
        RECT -27.850 -293.885 -27.680 -293.425 ;
        RECT -27.360 -294.140 -27.190 -293.345 ;
        RECT -26.900 -293.425 -26.670 -293.120 ;
        RECT -26.055 -293.175 -24.855 -292.865 ;
        RECT -24.675 -292.960 -21.845 -292.770 ;
        RECT -26.870 -293.885 -26.700 -293.425 ;
        RECT -26.055 -293.895 -25.755 -293.175 ;
        RECT -25.135 -294.140 -24.965 -293.345 ;
        RECT -24.675 -293.425 -24.445 -292.960 ;
        RECT -24.645 -293.885 -24.475 -293.425 ;
        RECT -24.155 -294.140 -23.985 -293.345 ;
        RECT -23.695 -293.425 -23.465 -292.960 ;
        RECT -22.715 -293.120 -21.845 -292.960 ;
        RECT -21.620 -292.680 -21.385 -291.945 ;
        RECT -21.100 -291.980 -20.930 -291.520 ;
        RECT -20.615 -291.625 -20.405 -291.350 ;
        RECT -21.105 -292.240 -20.925 -291.980 ;
        RECT -20.610 -292.060 -20.440 -291.625 ;
        RECT -20.120 -291.970 -19.950 -291.520 ;
        RECT -19.645 -291.630 -19.435 -291.350 ;
        RECT -20.120 -292.060 -19.935 -291.970 ;
        RECT -19.630 -292.060 -19.460 -291.630 ;
        RECT -19.140 -291.970 -18.970 -291.520 ;
        RECT -18.665 -291.605 -18.455 -291.350 ;
        RECT -8.095 -291.350 -4.955 -291.180 ;
        RECT -15.330 -291.465 -15.160 -291.445 ;
        RECT -20.115 -292.240 -19.935 -292.060 ;
        RECT -19.145 -292.240 -18.965 -291.970 ;
        RECT -18.650 -292.060 -18.480 -291.605 ;
        RECT -18.160 -292.020 -17.990 -291.520 ;
        RECT -18.175 -292.240 -17.965 -292.020 ;
        RECT -21.105 -292.410 -17.965 -292.240 ;
        RECT -21.620 -293.050 -20.760 -292.680 ;
        RECT -18.840 -292.945 -17.965 -292.410 ;
        RECT -15.360 -292.730 -15.130 -291.465 ;
        RECT -14.350 -292.405 -14.180 -291.445 ;
        RECT -13.370 -292.405 -13.200 -291.445 ;
        RECT -11.145 -291.465 -10.975 -291.445 ;
        RECT -12.250 -291.815 -11.965 -291.555 ;
        RECT -12.990 -292.125 -11.965 -291.815 ;
        RECT -14.380 -292.730 -14.150 -292.405 ;
        RECT -13.400 -292.730 -13.170 -292.405 ;
        RECT -15.360 -292.770 -13.170 -292.730 ;
        RECT -12.990 -292.770 -12.680 -292.125 ;
        RECT -12.250 -292.375 -11.965 -292.125 ;
        RECT -16.380 -292.840 -15.540 -292.805 ;
        RECT -23.665 -293.885 -23.495 -293.425 ;
        RECT -23.175 -294.140 -23.005 -293.345 ;
        RECT -22.715 -293.425 -22.485 -293.120 ;
        RECT -22.685 -293.885 -22.515 -293.425 ;
        RECT -21.620 -293.725 -21.385 -293.050 ;
        RECT -18.840 -293.245 -17.510 -292.945 ;
        RECT -16.490 -293.140 -15.540 -292.840 ;
        RECT -16.380 -293.175 -15.540 -293.140 ;
        RECT -15.360 -292.960 -12.680 -292.770 ;
        RECT -21.120 -293.415 -17.965 -293.245 ;
        RECT -21.120 -293.620 -20.915 -293.415 ;
        RECT -21.590 -294.075 -21.420 -293.725 ;
        RECT -29.365 -294.480 -22.510 -294.140 ;
        RECT -21.615 -294.365 -21.395 -294.075 ;
        RECT -21.100 -294.135 -20.930 -293.620 ;
        RECT -20.610 -294.020 -20.440 -293.595 ;
        RECT -20.130 -293.660 -19.925 -293.415 ;
        RECT -20.635 -294.365 -20.415 -294.020 ;
        RECT -20.120 -294.135 -19.950 -293.660 ;
        RECT -19.630 -294.020 -19.460 -293.595 ;
        RECT -19.160 -293.660 -18.955 -293.415 ;
        RECT -18.175 -293.450 -17.965 -293.415 ;
        RECT -19.655 -294.365 -19.435 -294.020 ;
        RECT -19.140 -294.135 -18.970 -293.660 ;
        RECT -18.650 -294.075 -18.480 -293.595 ;
        RECT -18.175 -293.665 -17.970 -293.450 ;
        RECT -18.670 -294.365 -18.450 -294.075 ;
        RECT -18.160 -294.135 -17.990 -293.665 ;
        RECT -15.820 -294.140 -15.650 -293.345 ;
        RECT -15.360 -293.425 -15.130 -292.960 ;
        RECT -15.330 -293.885 -15.160 -293.425 ;
        RECT -14.840 -294.140 -14.670 -293.345 ;
        RECT -14.380 -293.425 -14.150 -292.960 ;
        RECT -13.400 -293.120 -12.680 -292.960 ;
        RECT -11.175 -292.730 -10.945 -291.465 ;
        RECT -10.165 -292.405 -9.995 -291.445 ;
        RECT -9.185 -292.405 -9.015 -291.445 ;
        RECT -8.095 -291.575 -7.915 -291.350 ;
        RECT -10.195 -292.730 -9.965 -292.405 ;
        RECT -9.215 -292.730 -8.985 -292.405 ;
        RECT -11.175 -292.770 -8.985 -292.730 ;
        RECT -8.710 -292.650 -8.340 -291.810 ;
        RECT -8.090 -291.945 -7.920 -291.575 ;
        RECT -8.710 -292.770 -8.345 -292.650 ;
        RECT -11.175 -292.960 -8.345 -292.770 ;
        RECT -14.350 -293.885 -14.180 -293.425 ;
        RECT -13.860 -294.140 -13.690 -293.345 ;
        RECT -13.400 -293.425 -13.170 -293.120 ;
        RECT -13.370 -293.885 -13.200 -293.425 ;
        RECT -11.635 -294.140 -11.465 -293.345 ;
        RECT -11.175 -293.425 -10.945 -292.960 ;
        RECT -11.145 -293.885 -10.975 -293.425 ;
        RECT -10.655 -294.140 -10.485 -293.345 ;
        RECT -10.195 -293.425 -9.965 -292.960 ;
        RECT -9.215 -293.120 -8.345 -292.960 ;
        RECT -8.120 -292.680 -7.885 -291.945 ;
        RECT -7.600 -291.980 -7.430 -291.520 ;
        RECT -7.115 -291.625 -6.905 -291.350 ;
        RECT -7.605 -292.240 -7.425 -291.980 ;
        RECT -7.110 -292.060 -6.940 -291.625 ;
        RECT -6.620 -291.970 -6.450 -291.520 ;
        RECT -6.145 -291.630 -5.935 -291.350 ;
        RECT -6.620 -292.060 -6.435 -291.970 ;
        RECT -6.130 -292.060 -5.960 -291.630 ;
        RECT -5.640 -291.970 -5.470 -291.520 ;
        RECT -5.165 -291.605 -4.955 -291.350 ;
        RECT -6.615 -292.240 -6.435 -292.060 ;
        RECT -5.645 -292.240 -5.465 -291.970 ;
        RECT -5.150 -292.060 -4.980 -291.605 ;
        RECT -4.660 -292.020 -4.490 -291.520 ;
        RECT -3.270 -291.820 46.025 -290.515 ;
        RECT 74.755 -289.880 77.325 -289.065 ;
        RECT 83.555 -289.880 84.660 -289.740 ;
        RECT 74.755 -290.530 84.660 -289.880 ;
        RECT 74.755 -291.190 77.325 -290.530 ;
        RECT -4.675 -292.240 -4.465 -292.020 ;
        RECT -7.605 -292.410 -4.465 -292.240 ;
        RECT -8.120 -293.050 -7.260 -292.680 ;
        RECT -5.340 -292.955 -4.465 -292.410 ;
        RECT -10.165 -293.885 -9.995 -293.425 ;
        RECT -9.675 -294.140 -9.505 -293.345 ;
        RECT -9.215 -293.425 -8.985 -293.120 ;
        RECT -9.185 -293.885 -9.015 -293.425 ;
        RECT -8.120 -293.725 -7.885 -293.050 ;
        RECT -5.340 -293.245 -4.090 -292.955 ;
        RECT -7.620 -293.255 -4.090 -293.245 ;
        RECT -7.620 -293.415 -4.465 -293.255 ;
        RECT -7.620 -293.620 -7.415 -293.415 ;
        RECT -8.090 -294.075 -7.920 -293.725 ;
        RECT -28.125 -294.680 -27.570 -294.480 ;
        RECT -28.180 -294.720 -27.495 -294.680 ;
        RECT -24.070 -294.720 -23.515 -294.480 ;
        RECT -21.615 -294.535 -18.450 -294.365 ;
        RECT -15.865 -294.150 -13.195 -294.140 ;
        RECT -11.680 -294.150 -9.010 -294.140 ;
        RECT -15.865 -294.480 -9.010 -294.150 ;
        RECT -8.115 -294.365 -7.895 -294.075 ;
        RECT -7.600 -294.135 -7.430 -293.620 ;
        RECT -7.110 -294.020 -6.940 -293.595 ;
        RECT -6.630 -293.660 -6.425 -293.415 ;
        RECT -7.135 -294.365 -6.915 -294.020 ;
        RECT -6.620 -294.135 -6.450 -293.660 ;
        RECT -6.130 -294.020 -5.960 -293.595 ;
        RECT -5.660 -293.660 -5.455 -293.415 ;
        RECT -4.675 -293.450 -4.465 -293.415 ;
        RECT -6.155 -294.365 -5.935 -294.020 ;
        RECT -5.640 -294.135 -5.470 -293.660 ;
        RECT -5.150 -294.075 -4.980 -293.595 ;
        RECT -4.675 -293.665 -4.470 -293.450 ;
        RECT -5.170 -294.365 -4.950 -294.075 ;
        RECT -4.660 -294.135 -4.490 -293.665 ;
        RECT -15.080 -294.710 -14.525 -294.480 ;
        RECT -14.165 -294.490 -11.565 -294.480 ;
        RECT -15.195 -294.720 -14.510 -294.710 ;
        RECT -10.690 -294.720 -10.135 -294.480 ;
        RECT -8.115 -294.535 -4.950 -294.365 ;
        RECT -3.270 -294.710 -1.780 -291.820 ;
        RECT 1.960 -293.145 2.610 -291.820 ;
        RECT 3.490 -293.145 4.140 -291.820 ;
        RECT 5.075 -293.145 5.725 -291.820 ;
        RECT 7.305 -293.145 7.955 -291.820 ;
        RECT 1.895 -293.470 8.265 -293.145 ;
        RECT -3.270 -294.720 -1.345 -294.710 ;
        RECT -28.265 -294.915 -1.340 -294.720 ;
        RECT -28.180 -294.980 -27.495 -294.915 ;
        RECT -15.195 -295.010 -14.510 -294.915 ;
        RECT -2.005 -295.010 -1.345 -294.915 ;
        RECT -29.920 -295.720 -29.620 -295.035 ;
        RECT -26.235 -295.610 -25.575 -295.570 ;
        RECT -3.620 -295.610 -2.960 -295.560 ;
        RECT -34.170 -296.820 -33.935 -296.225 ;
        RECT -31.615 -296.820 -31.090 -296.790 ;
        RECT -37.260 -297.230 -31.090 -296.820 ;
        RECT -31.615 -297.265 -31.090 -297.230 ;
        RECT -29.915 -297.510 -29.675 -295.720 ;
        RECT -28.265 -295.805 -2.960 -295.610 ;
        RECT -26.235 -295.870 -25.575 -295.805 ;
        RECT -3.620 -295.860 -2.960 -295.805 ;
        RECT -29.325 -296.380 -26.655 -296.040 ;
        RECT -24.670 -296.155 -21.505 -295.985 ;
        RECT -29.320 -297.095 -29.150 -296.635 ;
        RECT -29.350 -297.400 -29.120 -297.095 ;
        RECT -28.830 -297.175 -28.660 -296.380 ;
        RECT -28.340 -297.095 -28.170 -296.635 ;
        RECT -29.500 -297.510 -29.120 -297.400 ;
        RECT -29.915 -297.560 -29.120 -297.510 ;
        RECT -28.370 -297.560 -28.140 -297.095 ;
        RECT -27.850 -297.175 -27.680 -296.380 ;
        RECT -27.360 -297.095 -27.190 -296.635 ;
        RECT -27.390 -297.560 -27.160 -297.095 ;
        RECT -26.870 -297.175 -26.700 -296.380 ;
        RECT -25.130 -296.855 -24.960 -296.385 ;
        RECT -24.670 -296.445 -24.450 -296.155 ;
        RECT -25.150 -297.070 -24.945 -296.855 ;
        RECT -24.640 -296.925 -24.470 -296.445 ;
        RECT -24.150 -296.860 -23.980 -296.385 ;
        RECT -23.685 -296.500 -23.465 -296.155 ;
        RECT -25.155 -297.105 -24.945 -297.070 ;
        RECT -24.165 -297.105 -23.960 -296.860 ;
        RECT -23.660 -296.925 -23.490 -296.500 ;
        RECT -23.170 -296.860 -23.000 -296.385 ;
        RECT -22.705 -296.500 -22.485 -296.155 ;
        RECT -23.195 -297.105 -22.990 -296.860 ;
        RECT -22.680 -296.925 -22.510 -296.500 ;
        RECT -22.190 -296.900 -22.020 -296.385 ;
        RECT -21.725 -296.445 -21.505 -296.155 ;
        RECT -20.610 -296.380 -13.155 -296.040 ;
        RECT -11.170 -296.155 -8.005 -295.985 ;
        RECT -21.700 -296.795 -21.530 -296.445 ;
        RECT -22.205 -297.105 -22.000 -296.900 ;
        RECT -25.155 -297.275 -22.000 -297.105 ;
        RECT -29.915 -297.695 -27.160 -297.560 ;
        RECT -29.910 -297.705 -27.160 -297.695 ;
        RECT -40.105 -297.740 -39.935 -297.720 ;
        RECT -29.500 -297.750 -27.160 -297.705 ;
        RECT -26.980 -297.420 -26.140 -297.345 ;
        RECT -25.155 -297.420 -24.280 -297.275 ;
        RECT -26.980 -297.685 -24.280 -297.420 ;
        RECT -21.735 -297.470 -21.500 -296.795 ;
        RECT -20.605 -297.095 -20.435 -296.635 ;
        RECT -20.635 -297.400 -20.405 -297.095 ;
        RECT -20.115 -297.175 -19.945 -296.380 ;
        RECT -19.625 -297.095 -19.455 -296.635 ;
        RECT -26.980 -297.715 -26.140 -297.685 ;
        RECT -50.535 -298.005 -47.395 -297.835 ;
        RECT -29.350 -297.790 -27.160 -297.750 ;
        RECT -29.350 -298.115 -29.120 -297.790 ;
        RECT -28.370 -298.115 -28.140 -297.790 ;
        RECT -76.565 -298.500 -76.040 -298.140 ;
        RECT -78.760 -301.985 -78.550 -301.765 ;
        RECT -77.690 -301.815 -77.520 -298.845 ;
        RECT -79.750 -302.155 -78.550 -301.985 ;
        RECT -106.285 -302.605 -102.265 -302.470 ;
        RECT -109.855 -303.430 -109.565 -303.415 ;
        RECT -100.580 -303.430 -100.290 -302.950 ;
        RECT -109.855 -303.635 -100.290 -303.430 ;
        RECT -109.855 -304.100 -109.565 -303.635 ;
        RECT -109.285 -303.825 -108.995 -303.820 ;
        RECT -96.475 -303.825 -96.185 -303.345 ;
        RECT -109.285 -304.030 -96.185 -303.825 ;
        RECT -109.285 -304.505 -108.995 -304.030 ;
        RECT -96.010 -304.210 -95.720 -303.730 ;
        RECT -108.560 -304.415 -95.720 -304.210 ;
        RECT -108.560 -304.895 -108.270 -304.415 ;
        RECT -107.350 -304.820 -102.435 -304.665 ;
        RECT -107.350 -305.145 -100.960 -304.820 ;
        RECT -107.350 -305.240 -102.435 -305.145 ;
        RECT -107.270 -310.665 -107.100 -306.085 ;
        RECT -106.780 -307.125 -106.610 -305.240 ;
        RECT -104.715 -305.595 -102.510 -305.425 ;
        RECT -105.205 -307.945 -105.035 -306.085 ;
        RECT -104.715 -307.625 -104.545 -305.595 ;
        RECT -103.665 -305.610 -102.510 -305.595 ;
        RECT -104.225 -307.945 -104.055 -306.085 ;
        RECT -103.665 -306.140 -103.490 -305.610 ;
        RECT -103.660 -307.625 -103.490 -306.140 ;
        RECT -103.170 -307.625 -103.000 -306.085 ;
        RECT -102.685 -306.130 -102.510 -305.610 ;
        RECT -102.680 -307.625 -102.510 -306.130 ;
        RECT -103.175 -307.940 -103.000 -307.625 ;
        RECT -102.110 -307.940 -101.940 -306.090 ;
        RECT -101.620 -307.630 -101.450 -305.145 ;
        RECT -87.890 -306.015 -87.720 -304.975 ;
        RECT -86.910 -306.015 -86.740 -304.975 ;
        RECT -85.930 -306.015 -85.760 -304.975 ;
        RECT -83.025 -306.050 -82.855 -304.330 ;
        RECT -82.045 -306.050 -81.875 -304.330 ;
        RECT -79.980 -304.865 -79.810 -304.325 ;
        RECT -79.000 -304.865 -78.830 -304.325 ;
        RECT -80.570 -305.100 -80.205 -305.035 ;
        RECT -81.070 -305.240 -80.205 -305.100 ;
        RECT -81.180 -305.305 -80.205 -305.240 ;
        RECT -81.180 -306.050 -80.875 -305.305 ;
        RECT -80.570 -305.335 -80.205 -305.305 ;
        RECT -78.020 -305.185 -77.850 -304.325 ;
        RECT -76.510 -305.185 -76.160 -298.500 ;
        RECT -29.320 -299.075 -29.150 -298.115 ;
        RECT -28.340 -299.075 -28.170 -298.115 ;
        RECT -27.390 -299.055 -27.160 -297.790 ;
        RECT -25.155 -298.110 -24.280 -297.685 ;
        RECT -22.360 -297.840 -21.500 -297.470 ;
        RECT -25.155 -298.280 -22.015 -298.110 ;
        RECT -25.155 -298.500 -24.945 -298.280 ;
        RECT -25.130 -299.000 -24.960 -298.500 ;
        RECT -24.640 -298.915 -24.470 -298.460 ;
        RECT -24.155 -298.550 -23.975 -298.280 ;
        RECT -23.185 -298.460 -23.005 -298.280 ;
        RECT -27.360 -299.075 -27.190 -299.055 ;
        RECT -24.665 -299.170 -24.455 -298.915 ;
        RECT -24.150 -299.000 -23.980 -298.550 ;
        RECT -23.660 -298.890 -23.490 -298.460 ;
        RECT -23.185 -298.550 -23.000 -298.460 ;
        RECT -23.685 -299.170 -23.475 -298.890 ;
        RECT -23.170 -299.000 -23.000 -298.550 ;
        RECT -22.680 -298.895 -22.510 -298.460 ;
        RECT -22.195 -298.540 -22.015 -298.280 ;
        RECT -22.715 -299.170 -22.505 -298.895 ;
        RECT -22.190 -299.000 -22.020 -298.540 ;
        RECT -21.735 -298.575 -21.500 -297.840 ;
        RECT -21.275 -297.560 -20.405 -297.400 ;
        RECT -19.655 -297.560 -19.425 -297.095 ;
        RECT -19.135 -297.175 -18.965 -296.380 ;
        RECT -18.645 -297.095 -18.475 -296.635 ;
        RECT -18.675 -297.560 -18.445 -297.095 ;
        RECT -18.155 -297.175 -17.985 -296.380 ;
        RECT -16.550 -297.455 -16.250 -296.880 ;
        RECT -15.820 -297.095 -15.650 -296.635 ;
        RECT -15.850 -297.400 -15.620 -297.095 ;
        RECT -15.330 -297.175 -15.160 -296.380 ;
        RECT -14.840 -297.095 -14.670 -296.635 ;
        RECT -16.000 -297.455 -15.620 -297.400 ;
        RECT -21.275 -297.750 -18.445 -297.560 ;
        RECT -21.275 -297.870 -20.910 -297.750 ;
        RECT -21.700 -298.945 -21.530 -298.575 ;
        RECT -21.280 -298.710 -20.910 -297.870 ;
        RECT -20.635 -297.790 -18.445 -297.750 ;
        RECT -20.635 -298.115 -20.405 -297.790 ;
        RECT -19.655 -298.115 -19.425 -297.790 ;
        RECT -21.705 -299.170 -21.525 -298.945 ;
        RECT -20.605 -299.075 -20.435 -298.115 ;
        RECT -19.625 -299.075 -19.455 -298.115 ;
        RECT -18.675 -299.055 -18.445 -297.790 ;
        RECT -16.575 -297.560 -15.620 -297.455 ;
        RECT -14.870 -297.560 -14.640 -297.095 ;
        RECT -14.350 -297.175 -14.180 -296.380 ;
        RECT -13.860 -297.095 -13.690 -296.635 ;
        RECT -13.890 -297.560 -13.660 -297.095 ;
        RECT -13.370 -297.175 -13.200 -296.380 ;
        RECT -11.645 -296.855 -11.415 -296.245 ;
        RECT -11.170 -296.445 -10.950 -296.155 ;
        RECT -11.650 -296.905 -11.415 -296.855 ;
        RECT -11.650 -297.070 -11.445 -296.905 ;
        RECT -11.140 -296.925 -10.970 -296.445 ;
        RECT -10.650 -296.860 -10.480 -296.385 ;
        RECT -10.185 -296.500 -9.965 -296.155 ;
        RECT -11.655 -297.105 -11.445 -297.070 ;
        RECT -10.665 -297.105 -10.460 -296.860 ;
        RECT -10.160 -296.925 -9.990 -296.500 ;
        RECT -9.670 -296.860 -9.500 -296.385 ;
        RECT -9.205 -296.500 -8.985 -296.155 ;
        RECT -9.695 -297.105 -9.490 -296.860 ;
        RECT -9.180 -296.925 -9.010 -296.500 ;
        RECT -8.690 -296.900 -8.520 -296.385 ;
        RECT -8.225 -296.445 -8.005 -296.155 ;
        RECT -7.110 -296.380 -0.030 -296.040 ;
        RECT -8.200 -296.795 -8.030 -296.445 ;
        RECT -8.705 -297.105 -8.500 -296.900 ;
        RECT -11.655 -297.275 -8.500 -297.105 ;
        RECT -16.575 -297.680 -13.660 -297.560 ;
        RECT -17.655 -298.350 -17.370 -298.145 ;
        RECT -16.575 -298.350 -16.350 -297.680 ;
        RECT -16.000 -297.750 -13.660 -297.680 ;
        RECT -13.480 -297.385 -12.640 -297.345 ;
        RECT -11.655 -297.385 -10.780 -297.275 ;
        RECT -13.480 -297.670 -10.780 -297.385 ;
        RECT -8.235 -297.470 -8.000 -296.795 ;
        RECT -7.105 -297.095 -6.935 -296.635 ;
        RECT -7.135 -297.400 -6.905 -297.095 ;
        RECT -6.615 -297.175 -6.445 -296.380 ;
        RECT -6.125 -297.095 -5.955 -296.635 ;
        RECT -13.480 -297.715 -12.640 -297.670 ;
        RECT -15.850 -297.790 -13.660 -297.750 ;
        RECT -15.850 -298.115 -15.620 -297.790 ;
        RECT -14.870 -298.115 -14.640 -297.790 ;
        RECT -17.655 -298.575 -16.350 -298.350 ;
        RECT -17.655 -298.965 -17.370 -298.575 ;
        RECT -18.645 -299.075 -18.475 -299.055 ;
        RECT -15.820 -299.075 -15.650 -298.115 ;
        RECT -14.840 -299.075 -14.670 -298.115 ;
        RECT -13.890 -299.055 -13.660 -297.790 ;
        RECT -11.655 -298.110 -10.780 -297.670 ;
        RECT -8.860 -297.840 -8.000 -297.470 ;
        RECT -11.655 -298.280 -8.515 -298.110 ;
        RECT -11.655 -298.500 -11.445 -298.280 ;
        RECT -11.630 -299.000 -11.460 -298.500 ;
        RECT -11.140 -298.915 -10.970 -298.460 ;
        RECT -10.655 -298.550 -10.475 -298.280 ;
        RECT -9.685 -298.460 -9.505 -298.280 ;
        RECT -13.860 -299.075 -13.690 -299.055 ;
        RECT -24.665 -299.340 -21.525 -299.170 ;
        RECT -11.165 -299.170 -10.955 -298.915 ;
        RECT -10.650 -299.000 -10.480 -298.550 ;
        RECT -10.160 -298.890 -9.990 -298.460 ;
        RECT -9.685 -298.550 -9.500 -298.460 ;
        RECT -10.185 -299.170 -9.975 -298.890 ;
        RECT -9.670 -299.000 -9.500 -298.550 ;
        RECT -9.180 -298.895 -9.010 -298.460 ;
        RECT -8.695 -298.540 -8.515 -298.280 ;
        RECT -9.215 -299.170 -9.005 -298.895 ;
        RECT -8.690 -299.000 -8.520 -298.540 ;
        RECT -8.235 -298.575 -8.000 -297.840 ;
        RECT -7.775 -297.560 -6.905 -297.400 ;
        RECT -6.155 -297.560 -5.925 -297.095 ;
        RECT -5.635 -297.175 -5.465 -296.380 ;
        RECT -5.145 -297.095 -4.975 -296.635 ;
        RECT -5.175 -297.560 -4.945 -297.095 ;
        RECT -4.655 -297.175 -4.485 -296.380 ;
        RECT -7.775 -297.750 -4.945 -297.560 ;
        RECT -4.765 -297.370 -3.925 -297.345 ;
        RECT -4.765 -297.430 -3.750 -297.370 ;
        RECT -3.465 -297.430 -3.165 -297.000 ;
        RECT -2.695 -297.095 -2.525 -296.635 ;
        RECT -2.725 -297.400 -2.495 -297.095 ;
        RECT -2.205 -297.175 -2.035 -296.380 ;
        RECT -1.715 -297.095 -1.545 -296.635 ;
        RECT -2.875 -297.430 -2.495 -297.400 ;
        RECT -4.765 -297.560 -2.495 -297.430 ;
        RECT -1.745 -297.560 -1.515 -297.095 ;
        RECT -1.225 -297.175 -1.055 -296.380 ;
        RECT -0.735 -297.095 -0.565 -296.635 ;
        RECT -0.765 -297.560 -0.535 -297.095 ;
        RECT -0.245 -297.175 -0.075 -296.380 ;
        RECT 1.955 -296.675 2.125 -294.410 ;
        RECT 2.445 -295.450 2.615 -293.470 ;
        RECT 4.510 -293.920 6.715 -293.750 ;
        RECT 4.020 -296.270 4.190 -294.410 ;
        RECT 4.510 -295.950 4.680 -293.920 ;
        RECT 5.560 -293.935 6.715 -293.920 ;
        RECT 5.000 -296.270 5.170 -294.410 ;
        RECT 5.560 -294.465 5.735 -293.935 ;
        RECT 5.565 -295.950 5.735 -294.465 ;
        RECT 6.055 -295.950 6.225 -294.410 ;
        RECT 6.540 -294.455 6.715 -293.935 ;
        RECT 6.545 -295.950 6.715 -294.455 ;
        RECT 6.050 -296.265 6.225 -295.950 ;
        RECT 7.115 -296.265 7.285 -294.415 ;
        RECT 7.605 -295.955 7.775 -293.470 ;
        RECT 11.925 -294.220 12.680 -291.820 ;
        RECT 13.810 -294.130 14.430 -291.820 ;
        RECT 15.460 -294.130 16.080 -291.820 ;
        RECT 17.495 -294.030 18.175 -293.800 ;
        RECT 13.810 -294.220 16.385 -294.130 ;
        RECT 6.050 -296.270 7.285 -296.265 ;
        RECT 8.095 -296.270 8.265 -294.415 ;
        RECT 4.020 -296.440 5.185 -296.270 ;
        RECT 6.050 -296.440 8.265 -296.270 ;
        RECT 11.925 -294.435 16.385 -294.220 ;
        RECT 11.925 -294.525 14.175 -294.435 ;
        RECT 1.200 -296.940 2.125 -296.675 ;
        RECT -4.765 -297.640 -0.535 -297.560 ;
        RECT -4.765 -297.660 -3.750 -297.640 ;
        RECT -3.465 -297.660 -3.165 -297.640 ;
        RECT -4.765 -297.715 -3.925 -297.660 ;
        RECT -2.875 -297.750 -0.535 -297.640 ;
        RECT -7.775 -297.870 -7.410 -297.750 ;
        RECT -8.200 -298.945 -8.030 -298.575 ;
        RECT -7.780 -298.710 -7.410 -297.870 ;
        RECT -7.135 -297.790 -4.945 -297.750 ;
        RECT -7.135 -298.115 -6.905 -297.790 ;
        RECT -6.155 -298.115 -5.925 -297.790 ;
        RECT -8.205 -299.170 -8.025 -298.945 ;
        RECT -7.105 -299.075 -6.935 -298.115 ;
        RECT -6.125 -299.075 -5.955 -298.115 ;
        RECT -5.175 -299.055 -4.945 -297.790 ;
        RECT -2.725 -297.790 -0.535 -297.750 ;
        RECT -2.725 -298.115 -2.495 -297.790 ;
        RECT -1.745 -298.115 -1.515 -297.790 ;
        RECT -4.155 -298.965 -3.870 -298.145 ;
        RECT -5.145 -299.075 -4.975 -299.055 ;
        RECT -2.695 -299.075 -2.525 -298.115 ;
        RECT -1.715 -299.075 -1.545 -298.115 ;
        RECT -0.765 -299.055 -0.535 -297.790 ;
        RECT 1.955 -298.990 2.125 -296.940 ;
        RECT 2.300 -296.710 2.975 -296.675 ;
        RECT 5.000 -296.710 5.185 -296.440 ;
        RECT 11.925 -296.560 12.230 -294.525 ;
        RECT 15.625 -294.695 15.800 -294.435 ;
        RECT 14.155 -296.235 14.325 -294.695 ;
        RECT 14.645 -296.235 14.815 -294.695 ;
        RECT 15.135 -296.235 15.305 -294.695 ;
        RECT 15.625 -296.235 15.795 -294.695 ;
        RECT 16.115 -296.235 16.285 -294.695 ;
        RECT 14.015 -296.450 14.385 -296.420 ;
        RECT 16.090 -296.450 16.445 -296.445 ;
        RECT 14.015 -296.455 16.445 -296.450 ;
        RECT 2.300 -296.895 5.185 -296.710 ;
        RECT 2.300 -296.945 2.975 -296.895 ;
        RECT 5.000 -297.585 5.185 -296.895 ;
        RECT 5.355 -296.720 6.030 -296.685 ;
        RECT 5.355 -296.890 10.135 -296.720 ;
        RECT 5.355 -296.955 6.030 -296.890 ;
        RECT 6.295 -297.110 6.970 -297.075 ;
        RECT 9.110 -297.110 9.790 -297.075 ;
        RECT 6.295 -297.300 9.790 -297.110 ;
        RECT 6.295 -297.345 6.970 -297.300 ;
        RECT 9.110 -297.305 9.790 -297.300 ;
        RECT 5.000 -297.770 7.775 -297.585 ;
        RECT 7.975 -297.755 8.935 -297.485 ;
        RECT 9.965 -297.715 10.135 -296.890 ;
        RECT 10.375 -296.990 13.450 -296.560 ;
        RECT 14.015 -296.645 17.350 -296.455 ;
        RECT 14.015 -296.775 14.385 -296.645 ;
        RECT 16.440 -296.655 17.350 -296.645 ;
        RECT 16.035 -296.925 16.710 -296.895 ;
        RECT 16.035 -296.945 16.860 -296.925 ;
        RECT 5.645 -298.990 5.815 -297.770 ;
        RECT 6.625 -298.990 6.795 -297.770 ;
        RECT 7.605 -298.990 7.775 -297.770 ;
        RECT 8.705 -298.175 8.935 -297.755 ;
        RECT 9.935 -298.065 10.790 -297.715 ;
        RECT 11.110 -297.770 11.280 -297.230 ;
        RECT 11.600 -297.770 11.770 -296.990 ;
        RECT 12.090 -297.770 12.260 -297.230 ;
        RECT 12.580 -297.770 12.750 -296.990 ;
        RECT 13.700 -297.050 15.795 -297.010 ;
        RECT 13.645 -297.200 15.795 -297.050 ;
        RECT 16.035 -297.125 16.970 -296.945 ;
        RECT 16.035 -297.165 16.925 -297.125 ;
        RECT 10.620 -298.925 10.790 -298.065 ;
        RECT 12.975 -297.945 13.340 -297.915 ;
        RECT 13.645 -297.945 13.950 -297.200 ;
        RECT 12.975 -298.010 13.950 -297.945 ;
        RECT 12.975 -298.150 13.840 -298.010 ;
        RECT 12.975 -298.215 13.340 -298.150 ;
        RECT 11.600 -298.925 11.770 -298.385 ;
        RECT 12.580 -298.925 12.750 -298.385 ;
        RECT 14.645 -298.920 14.815 -297.200 ;
        RECT 15.625 -298.920 15.795 -297.200 ;
        RECT -0.735 -299.075 -0.565 -299.055 ;
        RECT -11.165 -299.340 -8.025 -299.170 ;
        RECT 16.745 -300.915 16.925 -297.165 ;
        RECT -30.975 -301.190 -30.295 -300.960 ;
        RECT 16.150 -301.145 16.925 -300.915 ;
        RECT -103.175 -307.945 -101.940 -307.940 ;
        RECT -101.130 -307.945 -100.960 -306.090 ;
        RECT -83.940 -306.115 -83.265 -306.085 ;
        RECT -84.040 -306.125 -83.265 -306.115 ;
        RECT -89.350 -306.250 -88.700 -306.165 ;
        RECT -88.480 -306.250 -88.115 -306.185 ;
        RECT -92.025 -306.280 -91.735 -306.275 ;
        RECT -89.350 -306.280 -88.115 -306.250 ;
        RECT -92.025 -306.455 -88.115 -306.280 ;
        RECT -85.075 -306.305 -83.265 -306.125 ;
        RECT -83.025 -306.200 -80.875 -306.050 ;
        RECT -83.025 -306.240 -80.930 -306.200 ;
        RECT -79.980 -306.260 -79.810 -305.480 ;
        RECT -79.490 -306.020 -79.320 -305.480 ;
        RECT -79.000 -306.260 -78.830 -305.480 ;
        RECT -78.510 -306.020 -78.340 -305.480 ;
        RECT -78.020 -305.535 -76.160 -305.185 ;
        RECT -84.040 -306.315 -83.265 -306.305 ;
        RECT -83.940 -306.355 -83.265 -306.315 ;
        RECT -92.025 -306.620 -88.700 -306.455 ;
        RECT -88.480 -306.485 -88.115 -306.455 ;
        RECT -92.025 -306.960 -91.735 -306.620 ;
        RECT -89.350 -306.915 -88.700 -306.620 ;
        RECT -86.415 -306.605 -83.670 -306.595 ;
        RECT -81.615 -306.605 -81.245 -306.475 ;
        RECT -86.415 -306.625 -81.245 -306.605 ;
        RECT -105.205 -308.115 -104.040 -307.945 ;
        RECT -103.175 -308.115 -100.960 -307.945 ;
        RECT -106.925 -308.385 -106.250 -308.350 ;
        RECT -104.225 -308.385 -104.040 -308.115 ;
        RECT -106.925 -308.570 -104.040 -308.385 ;
        RECT -106.925 -308.620 -106.250 -308.570 ;
        RECT -104.225 -309.260 -104.040 -308.570 ;
        RECT -103.870 -308.395 -103.195 -308.360 ;
        RECT -100.725 -308.395 -100.435 -307.880 ;
        RECT -87.890 -307.905 -87.720 -306.625 ;
        RECT -87.400 -307.665 -87.230 -306.625 ;
        RECT -86.910 -307.905 -86.740 -306.625 ;
        RECT -86.420 -306.795 -81.245 -306.625 ;
        RECT -80.680 -306.690 -76.755 -306.260 ;
        RECT -86.420 -307.665 -86.250 -306.795 ;
        RECT -83.675 -306.800 -81.245 -306.795 ;
        RECT -83.675 -306.805 -83.320 -306.800 ;
        RECT -81.615 -306.830 -81.245 -306.800 ;
        RECT -103.870 -308.565 -100.435 -308.395 ;
        RECT -103.870 -308.630 -103.195 -308.565 ;
        RECT -102.930 -308.785 -102.255 -308.750 ;
        RECT -97.075 -308.785 -96.785 -308.290 ;
        RECT -88.590 -308.335 -83.900 -307.905 ;
        RECT -102.930 -308.975 -96.785 -308.785 ;
        RECT -102.930 -309.020 -102.255 -308.975 ;
        RECT -101.250 -309.205 -100.575 -309.160 ;
        RECT -92.450 -309.205 -92.160 -308.720 ;
        RECT -84.330 -308.740 -83.900 -308.335 ;
        RECT -83.515 -308.555 -83.345 -307.015 ;
        RECT -83.025 -308.555 -82.855 -307.015 ;
        RECT -82.535 -308.555 -82.365 -307.015 ;
        RECT -82.045 -308.555 -81.875 -307.015 ;
        RECT -81.555 -308.555 -81.385 -307.015 ;
        RECT -83.030 -308.740 -82.855 -308.555 ;
        RECT -79.460 -308.725 -79.155 -306.690 ;
        RECT -81.405 -308.740 -79.155 -308.725 ;
        RECT -84.330 -309.030 -79.155 -308.740 ;
        RECT -30.775 -308.845 -30.605 -301.190 ;
        RECT -18.575 -301.555 -17.895 -301.325 ;
        RECT 17.150 -301.335 17.350 -296.655 ;
        RECT 17.825 -297.705 18.175 -294.030 ;
        RECT 19.950 -294.210 20.705 -291.820 ;
        RECT 22.160 -294.120 22.915 -291.820 ;
        RECT 23.625 -294.120 24.380 -291.820 ;
        RECT 26.825 -293.190 27.555 -291.820 ;
        RECT 29.050 -293.190 29.780 -291.820 ;
        RECT 30.380 -293.190 31.110 -291.820 ;
        RECT 32.180 -293.190 32.910 -291.820 ;
        RECT 25.335 -293.470 26.015 -293.240 ;
        RECT 22.160 -294.210 24.410 -294.120 ;
        RECT 19.950 -294.425 24.410 -294.210 ;
        RECT 19.950 -294.515 22.200 -294.425 ;
        RECT 19.950 -296.550 20.255 -294.515 ;
        RECT 23.650 -294.685 23.825 -294.425 ;
        RECT 22.180 -296.225 22.350 -294.685 ;
        RECT 22.670 -296.225 22.840 -294.685 ;
        RECT 23.160 -296.225 23.330 -294.685 ;
        RECT 23.650 -296.225 23.820 -294.685 ;
        RECT 24.140 -296.225 24.310 -294.685 ;
        RECT 25.685 -295.745 26.010 -293.470 ;
        RECT 26.705 -293.515 33.075 -293.190 ;
        RECT 26.765 -295.745 26.935 -294.455 ;
        RECT 27.255 -295.495 27.425 -293.515 ;
        RECT 29.320 -293.965 31.525 -293.795 ;
        RECT 25.685 -296.035 26.935 -295.745 ;
        RECT 22.040 -296.440 22.410 -296.410 ;
        RECT 24.115 -296.440 24.470 -296.435 ;
        RECT 22.040 -296.445 24.470 -296.440 ;
        RECT 18.400 -296.980 21.475 -296.550 ;
        RECT 22.040 -296.635 25.490 -296.445 ;
        RECT 22.040 -296.765 22.410 -296.635 ;
        RECT 24.465 -296.645 25.490 -296.635 ;
        RECT 24.060 -296.925 24.735 -296.885 ;
        RECT 24.060 -296.935 24.995 -296.925 ;
        RECT 17.825 -298.055 18.815 -297.705 ;
        RECT 19.135 -297.760 19.305 -297.220 ;
        RECT 19.625 -297.760 19.795 -296.980 ;
        RECT 20.115 -297.760 20.285 -297.220 ;
        RECT 20.605 -297.760 20.775 -296.980 ;
        RECT 21.725 -297.040 23.820 -297.000 ;
        RECT 21.670 -297.190 23.820 -297.040 ;
        RECT 24.060 -297.125 25.095 -296.935 ;
        RECT 24.060 -297.155 24.735 -297.125 ;
        RECT 18.645 -298.915 18.815 -298.055 ;
        RECT 21.000 -297.935 21.365 -297.905 ;
        RECT 21.670 -297.935 21.975 -297.190 ;
        RECT 21.000 -298.000 21.975 -297.935 ;
        RECT 21.000 -298.140 21.865 -298.000 ;
        RECT 21.000 -298.205 21.365 -298.140 ;
        RECT 19.625 -298.915 19.795 -298.375 ;
        RECT 20.605 -298.915 20.775 -298.375 ;
        RECT 22.670 -298.910 22.840 -297.190 ;
        RECT 23.650 -298.910 23.820 -297.190 ;
        RECT -18.575 -302.820 -18.375 -301.555 ;
        RECT 16.670 -301.565 17.350 -301.335 ;
        RECT -18.590 -303.500 -18.360 -302.820 ;
        RECT 24.915 -303.760 25.095 -297.125 ;
        RECT 17.490 -303.940 25.095 -303.760 ;
        RECT 17.490 -304.500 17.670 -303.940 ;
        RECT 25.290 -304.110 25.490 -296.645 ;
        RECT 26.765 -299.035 26.935 -296.035 ;
        RECT 28.830 -296.315 29.000 -294.455 ;
        RECT 29.320 -295.995 29.490 -293.965 ;
        RECT 30.370 -293.980 31.525 -293.965 ;
        RECT 29.810 -296.315 29.980 -294.455 ;
        RECT 30.370 -294.510 30.545 -293.980 ;
        RECT 30.375 -295.995 30.545 -294.510 ;
        RECT 30.865 -295.995 31.035 -294.455 ;
        RECT 31.350 -294.500 31.525 -293.980 ;
        RECT 31.355 -295.995 31.525 -294.500 ;
        RECT 30.860 -296.310 31.035 -295.995 ;
        RECT 31.925 -296.310 32.095 -294.460 ;
        RECT 32.415 -296.000 32.585 -293.515 ;
        RECT 35.000 -294.090 35.985 -291.820 ;
        RECT 37.665 -294.090 38.650 -291.820 ;
        RECT 40.230 -294.045 41.215 -291.820 ;
        RECT 42.745 -294.045 43.730 -291.820 ;
        RECT 44.720 -293.955 46.025 -291.820 ;
        RECT 52.445 -291.505 52.765 -291.390 ;
        RECT 79.270 -291.505 79.685 -290.530 ;
        RECT 83.555 -290.640 84.660 -290.530 ;
        RECT 52.445 -291.920 79.685 -291.505 ;
        RECT 52.445 -291.980 52.765 -291.920 ;
        RECT 98.970 -292.310 99.715 -279.635 ;
        RECT 101.775 -282.285 102.695 -279.635 ;
        RECT 104.895 -279.805 105.105 -279.585 ;
        RECT 105.410 -279.625 105.580 -279.170 ;
        RECT 105.900 -279.535 106.070 -279.085 ;
        RECT 106.365 -279.195 106.575 -278.915 ;
        RECT 105.895 -279.805 106.075 -279.535 ;
        RECT 106.390 -279.625 106.560 -279.195 ;
        RECT 106.880 -279.535 107.050 -279.085 ;
        RECT 107.335 -279.190 107.545 -278.915 ;
        RECT 106.865 -279.625 107.050 -279.535 ;
        RECT 107.370 -279.625 107.540 -279.190 ;
        RECT 107.860 -279.545 108.030 -279.085 ;
        RECT 108.345 -279.140 108.525 -278.915 ;
        RECT 118.885 -278.915 122.025 -278.745 ;
        RECT 108.350 -279.510 108.520 -279.140 ;
        RECT 106.865 -279.805 107.045 -279.625 ;
        RECT 107.855 -279.805 108.035 -279.545 ;
        RECT 104.895 -279.975 108.035 -279.805 ;
        RECT 104.895 -280.520 105.770 -279.975 ;
        RECT 108.315 -280.245 108.550 -279.510 ;
        RECT 108.770 -280.215 109.140 -279.375 ;
        RECT 109.445 -279.970 109.615 -279.010 ;
        RECT 110.425 -279.970 110.595 -279.010 ;
        RECT 111.405 -279.030 111.575 -279.010 ;
        RECT 104.520 -280.810 105.770 -280.520 ;
        RECT 107.690 -280.615 108.550 -280.245 ;
        RECT 104.520 -280.820 108.050 -280.810 ;
        RECT 104.895 -280.980 108.050 -280.820 ;
        RECT 104.895 -281.015 105.105 -280.980 ;
        RECT 104.900 -281.230 105.105 -281.015 ;
        RECT 104.920 -281.700 105.090 -281.230 ;
        RECT 105.410 -281.640 105.580 -281.160 ;
        RECT 105.885 -281.225 106.090 -280.980 ;
        RECT 105.380 -281.930 105.600 -281.640 ;
        RECT 105.900 -281.700 106.070 -281.225 ;
        RECT 106.390 -281.585 106.560 -281.160 ;
        RECT 106.855 -281.225 107.060 -280.980 ;
        RECT 106.365 -281.930 106.585 -281.585 ;
        RECT 106.880 -281.700 107.050 -281.225 ;
        RECT 107.370 -281.585 107.540 -281.160 ;
        RECT 107.845 -281.185 108.050 -280.980 ;
        RECT 107.345 -281.930 107.565 -281.585 ;
        RECT 107.860 -281.700 108.030 -281.185 ;
        RECT 108.315 -281.290 108.550 -280.615 ;
        RECT 108.775 -280.335 109.140 -280.215 ;
        RECT 109.415 -280.295 109.645 -279.970 ;
        RECT 110.395 -280.295 110.625 -279.970 ;
        RECT 111.375 -280.295 111.605 -279.030 ;
        RECT 112.395 -279.380 112.680 -279.120 ;
        RECT 112.395 -279.690 113.420 -279.380 ;
        RECT 112.395 -279.940 112.680 -279.690 ;
        RECT 109.415 -280.335 111.605 -280.295 ;
        RECT 108.775 -280.525 111.605 -280.335 ;
        RECT 108.775 -280.685 109.645 -280.525 ;
        RECT 109.415 -280.990 109.645 -280.685 ;
        RECT 108.350 -281.640 108.520 -281.290 ;
        RECT 109.445 -281.450 109.615 -280.990 ;
        RECT 108.325 -281.930 108.545 -281.640 ;
        RECT 109.935 -281.705 110.105 -280.910 ;
        RECT 110.395 -280.990 110.625 -280.525 ;
        RECT 110.425 -281.450 110.595 -280.990 ;
        RECT 110.915 -281.705 111.085 -280.910 ;
        RECT 111.375 -280.990 111.605 -280.525 ;
        RECT 113.110 -280.335 113.420 -279.690 ;
        RECT 113.630 -279.970 113.800 -279.010 ;
        RECT 114.610 -279.970 114.780 -279.010 ;
        RECT 115.590 -279.030 115.760 -279.010 ;
        RECT 113.600 -280.295 113.830 -279.970 ;
        RECT 114.580 -280.295 114.810 -279.970 ;
        RECT 115.560 -280.295 115.790 -279.030 ;
        RECT 118.420 -279.585 118.590 -279.085 ;
        RECT 118.885 -279.170 119.095 -278.915 ;
        RECT 113.600 -280.335 115.790 -280.295 ;
        RECT 113.110 -280.525 115.790 -280.335 ;
        RECT 118.395 -279.805 118.605 -279.585 ;
        RECT 118.910 -279.625 119.080 -279.170 ;
        RECT 119.400 -279.535 119.570 -279.085 ;
        RECT 119.865 -279.195 120.075 -278.915 ;
        RECT 119.395 -279.805 119.575 -279.535 ;
        RECT 119.890 -279.625 120.060 -279.195 ;
        RECT 120.380 -279.535 120.550 -279.085 ;
        RECT 120.835 -279.190 121.045 -278.915 ;
        RECT 120.365 -279.625 120.550 -279.535 ;
        RECT 120.870 -279.625 121.040 -279.190 ;
        RECT 121.360 -279.545 121.530 -279.085 ;
        RECT 121.845 -279.140 122.025 -278.915 ;
        RECT 147.150 -278.930 147.320 -277.210 ;
        RECT 148.130 -278.930 148.300 -277.210 ;
        RECT 148.995 -277.955 149.300 -277.210 ;
        RECT 150.195 -277.780 150.365 -277.000 ;
        RECT 150.685 -277.780 150.855 -277.240 ;
        RECT 151.175 -277.780 151.345 -277.000 ;
        RECT 183.025 -277.065 184.260 -276.860 ;
        RECT 188.435 -277.000 189.110 -276.960 ;
        RECT 188.335 -277.010 189.110 -277.000 ;
        RECT 183.025 -277.150 183.675 -277.065 ;
        RECT 183.895 -277.130 184.260 -277.065 ;
        RECT 187.300 -277.190 189.110 -277.010 ;
        RECT 191.695 -277.055 195.620 -276.625 ;
        RECT 227.340 -277.055 227.990 -276.595 ;
        RECT 228.800 -276.885 228.970 -275.605 ;
        RECT 229.290 -276.885 229.460 -275.845 ;
        RECT 229.780 -276.885 229.950 -275.605 ;
        RECT 230.270 -276.715 230.440 -275.845 ;
        RECT 233.175 -276.495 233.345 -274.955 ;
        RECT 233.665 -276.495 233.835 -274.955 ;
        RECT 234.155 -276.495 234.325 -274.955 ;
        RECT 234.645 -276.495 234.815 -274.955 ;
        RECT 235.135 -276.495 235.305 -274.955 ;
        RECT 233.015 -276.710 233.370 -276.705 ;
        RECT 235.075 -276.710 235.445 -276.680 ;
        RECT 233.015 -276.715 235.445 -276.710 ;
        RECT 230.270 -276.885 235.445 -276.715 ;
        RECT 237.230 -276.820 237.535 -274.785 ;
        RECT 261.005 -274.625 262.135 -274.580 ;
        RECT 269.270 -274.625 270.500 -274.225 ;
        RECT 261.005 -275.290 270.500 -274.625 ;
        RECT 278.350 -274.310 281.675 -274.170 ;
        RECT 278.350 -274.600 283.525 -274.310 ;
        RECT 278.350 -275.005 278.780 -274.600 ;
        RECT 279.650 -274.785 279.825 -274.600 ;
        RECT 281.275 -274.615 283.525 -274.600 ;
        RECT 261.005 -275.750 262.135 -275.290 ;
        RECT 269.270 -275.325 270.500 -275.290 ;
        RECT 274.090 -275.435 278.780 -275.005 ;
        RECT 230.275 -276.905 235.445 -276.885 ;
        RECT 230.275 -276.915 233.020 -276.905 ;
        RECT 228.210 -277.055 228.575 -277.025 ;
        RECT 235.075 -277.035 235.445 -276.905 ;
        RECT 188.335 -277.200 189.110 -277.190 ;
        RECT 188.435 -277.230 189.110 -277.200 ;
        RECT 189.350 -277.115 191.445 -277.075 ;
        RECT 151.665 -277.780 151.835 -277.240 ;
        RECT 189.350 -277.265 191.500 -277.115 ;
        RECT 149.605 -277.955 149.970 -277.925 ;
        RECT 148.995 -278.020 149.970 -277.955 ;
        RECT 149.105 -278.160 149.970 -278.020 ;
        RECT 149.605 -278.225 149.970 -278.160 ;
        RECT 152.155 -278.075 154.015 -277.725 ;
        RECT 150.195 -278.935 150.365 -278.395 ;
        RECT 151.175 -278.935 151.345 -278.395 ;
        RECT 152.155 -278.935 152.325 -278.075 ;
        RECT 121.850 -279.510 122.020 -279.140 ;
        RECT 120.365 -279.805 120.545 -279.625 ;
        RECT 121.355 -279.805 121.535 -279.545 ;
        RECT 118.395 -279.975 121.535 -279.805 ;
        RECT 113.110 -280.685 113.830 -280.525 ;
        RECT 111.405 -281.450 111.575 -280.990 ;
        RECT 111.895 -281.705 112.065 -280.910 ;
        RECT 113.600 -280.990 113.830 -280.685 ;
        RECT 113.630 -281.450 113.800 -280.990 ;
        RECT 114.120 -281.705 114.290 -280.910 ;
        RECT 114.580 -280.990 114.810 -280.525 ;
        RECT 114.610 -281.450 114.780 -280.990 ;
        RECT 115.100 -281.705 115.270 -280.910 ;
        RECT 115.560 -280.990 115.790 -280.525 ;
        RECT 115.970 -280.405 116.810 -280.370 ;
        RECT 115.970 -280.705 116.920 -280.405 ;
        RECT 118.395 -280.510 119.270 -279.975 ;
        RECT 121.815 -280.245 122.050 -279.510 ;
        RECT 122.270 -280.215 122.640 -279.375 ;
        RECT 122.945 -279.970 123.115 -279.010 ;
        RECT 123.925 -279.970 124.095 -279.010 ;
        RECT 124.905 -279.030 125.075 -279.010 ;
        RECT 115.970 -280.740 116.810 -280.705 ;
        RECT 117.940 -280.810 119.270 -280.510 ;
        RECT 121.190 -280.615 122.050 -280.245 ;
        RECT 115.590 -281.450 115.760 -280.990 ;
        RECT 116.080 -281.705 116.250 -280.910 ;
        RECT 118.395 -280.980 121.550 -280.810 ;
        RECT 118.395 -281.015 118.605 -280.980 ;
        RECT 118.400 -281.230 118.605 -281.015 ;
        RECT 118.420 -281.700 118.590 -281.230 ;
        RECT 118.910 -281.640 119.080 -281.160 ;
        RECT 119.385 -281.225 119.590 -280.980 ;
        RECT 105.380 -282.100 108.545 -281.930 ;
        RECT 109.440 -281.715 112.110 -281.705 ;
        RECT 113.625 -281.715 116.295 -281.705 ;
        RECT 109.440 -282.045 116.295 -281.715 ;
        RECT 118.880 -281.930 119.100 -281.640 ;
        RECT 119.400 -281.700 119.570 -281.225 ;
        RECT 119.890 -281.585 120.060 -281.160 ;
        RECT 120.355 -281.225 120.560 -280.980 ;
        RECT 119.865 -281.930 120.085 -281.585 ;
        RECT 120.380 -281.700 120.550 -281.225 ;
        RECT 120.870 -281.585 121.040 -281.160 ;
        RECT 121.345 -281.185 121.550 -280.980 ;
        RECT 120.845 -281.930 121.065 -281.585 ;
        RECT 121.360 -281.700 121.530 -281.185 ;
        RECT 121.815 -281.290 122.050 -280.615 ;
        RECT 122.275 -280.335 122.640 -280.215 ;
        RECT 122.915 -280.295 123.145 -279.970 ;
        RECT 123.895 -280.295 124.125 -279.970 ;
        RECT 124.875 -280.295 125.105 -279.030 ;
        RECT 125.895 -279.440 126.180 -279.120 ;
        RECT 125.895 -279.685 126.895 -279.440 ;
        RECT 125.895 -279.940 126.180 -279.685 ;
        RECT 122.915 -280.335 125.105 -280.295 ;
        RECT 122.275 -280.525 125.105 -280.335 ;
        RECT 126.665 -280.335 126.895 -279.685 ;
        RECT 127.130 -279.970 127.300 -279.010 ;
        RECT 128.110 -279.970 128.280 -279.010 ;
        RECT 129.090 -279.030 129.260 -279.010 ;
        RECT 127.100 -280.295 127.330 -279.970 ;
        RECT 128.080 -280.295 128.310 -279.970 ;
        RECT 129.060 -280.295 129.290 -279.030 ;
        RECT 127.100 -280.335 129.290 -280.295 ;
        RECT 122.275 -280.685 123.145 -280.525 ;
        RECT 122.915 -280.990 123.145 -280.685 ;
        RECT 121.850 -281.640 122.020 -281.290 ;
        RECT 122.945 -281.450 123.115 -280.990 ;
        RECT 121.825 -281.930 122.045 -281.640 ;
        RECT 123.435 -281.705 123.605 -280.910 ;
        RECT 123.895 -280.990 124.125 -280.525 ;
        RECT 123.925 -281.450 124.095 -280.990 ;
        RECT 124.415 -281.705 124.585 -280.910 ;
        RECT 124.875 -280.990 125.105 -280.525 ;
        RECT 125.285 -280.425 126.125 -280.370 ;
        RECT 125.285 -280.430 126.300 -280.425 ;
        RECT 125.285 -280.740 126.485 -280.430 ;
        RECT 126.665 -280.525 129.290 -280.335 ;
        RECT 126.665 -280.685 127.330 -280.525 ;
        RECT 124.905 -281.450 125.075 -280.990 ;
        RECT 125.395 -281.705 125.565 -280.910 ;
        RECT 126.185 -281.460 126.485 -280.740 ;
        RECT 127.100 -280.990 127.330 -280.685 ;
        RECT 127.130 -281.450 127.300 -280.990 ;
        RECT 127.620 -281.705 127.790 -280.910 ;
        RECT 128.080 -280.990 128.310 -280.525 ;
        RECT 128.110 -281.450 128.280 -280.990 ;
        RECT 128.600 -281.705 128.770 -280.910 ;
        RECT 129.060 -280.990 129.290 -280.525 ;
        RECT 129.470 -280.520 130.310 -280.370 ;
        RECT 129.470 -280.740 130.345 -280.520 ;
        RECT 129.090 -281.450 129.260 -280.990 ;
        RECT 129.580 -281.705 129.750 -280.910 ;
        RECT 110.565 -282.285 111.120 -282.045 ;
        RECT 111.995 -282.055 114.595 -282.045 ;
        RECT 114.955 -282.275 115.510 -282.045 ;
        RECT 118.880 -282.100 122.045 -281.930 ;
        RECT 122.940 -282.045 129.795 -281.705 ;
        RECT 114.940 -282.285 115.625 -282.275 ;
        RECT 123.945 -282.285 124.500 -282.045 ;
        RECT 128.000 -282.245 128.555 -282.045 ;
        RECT 127.925 -282.285 128.610 -282.245 ;
        RECT 101.770 -282.480 128.695 -282.285 ;
        RECT 101.775 -282.575 102.435 -282.480 ;
        RECT 114.940 -282.575 115.625 -282.480 ;
        RECT 127.925 -282.545 128.610 -282.480 ;
        RECT 130.105 -282.600 130.345 -280.740 ;
        RECT 150.425 -281.275 151.625 -281.105 ;
        RECT 103.390 -283.175 104.050 -283.125 ;
        RECT 126.005 -283.175 126.665 -283.135 ;
        RECT 103.390 -283.370 128.695 -283.175 ;
        RECT 130.050 -283.285 130.350 -282.600 ;
        RECT 103.390 -283.425 104.050 -283.370 ;
        RECT 126.005 -283.435 126.665 -283.370 ;
        RECT 100.460 -283.945 107.540 -283.605 ;
        RECT 108.435 -283.720 111.600 -283.550 ;
        RECT 100.505 -284.740 100.675 -283.945 ;
        RECT 100.995 -284.660 101.165 -284.200 ;
        RECT 100.965 -285.125 101.195 -284.660 ;
        RECT 101.485 -284.740 101.655 -283.945 ;
        RECT 101.975 -284.660 102.145 -284.200 ;
        RECT 101.945 -285.125 102.175 -284.660 ;
        RECT 102.465 -284.740 102.635 -283.945 ;
        RECT 102.955 -284.660 103.125 -284.200 ;
        RECT 102.925 -284.965 103.155 -284.660 ;
        RECT 102.925 -284.995 103.305 -284.965 ;
        RECT 103.595 -284.995 103.895 -284.565 ;
        RECT 104.915 -284.740 105.085 -283.945 ;
        RECT 105.405 -284.660 105.575 -284.200 ;
        RECT 104.355 -284.935 105.195 -284.910 ;
        RECT 104.180 -284.995 105.195 -284.935 ;
        RECT 102.925 -285.125 105.195 -284.995 ;
        RECT 100.965 -285.205 105.195 -285.125 ;
        RECT 100.965 -285.315 103.305 -285.205 ;
        RECT 103.595 -285.225 103.895 -285.205 ;
        RECT 104.180 -285.225 105.195 -285.205 ;
        RECT 104.355 -285.280 105.195 -285.225 ;
        RECT 105.375 -285.125 105.605 -284.660 ;
        RECT 105.895 -284.740 106.065 -283.945 ;
        RECT 106.385 -284.660 106.555 -284.200 ;
        RECT 106.355 -285.125 106.585 -284.660 ;
        RECT 106.875 -284.740 107.045 -283.945 ;
        RECT 108.435 -284.010 108.655 -283.720 ;
        RECT 107.365 -284.660 107.535 -284.200 ;
        RECT 108.460 -284.360 108.630 -284.010 ;
        RECT 107.335 -284.965 107.565 -284.660 ;
        RECT 107.335 -285.125 108.205 -284.965 ;
        RECT 105.375 -285.315 108.205 -285.125 ;
        RECT 100.965 -285.355 103.155 -285.315 ;
        RECT 100.965 -286.620 101.195 -285.355 ;
        RECT 101.945 -285.680 102.175 -285.355 ;
        RECT 102.925 -285.680 103.155 -285.355 ;
        RECT 105.375 -285.355 107.565 -285.315 ;
        RECT 100.995 -286.640 101.165 -286.620 ;
        RECT 101.975 -286.640 102.145 -285.680 ;
        RECT 102.955 -286.640 103.125 -285.680 ;
        RECT 104.300 -286.530 104.585 -285.710 ;
        RECT 105.375 -286.620 105.605 -285.355 ;
        RECT 106.355 -285.680 106.585 -285.355 ;
        RECT 107.335 -285.680 107.565 -285.355 ;
        RECT 107.840 -285.435 108.205 -285.315 ;
        RECT 108.430 -285.035 108.665 -284.360 ;
        RECT 108.950 -284.465 109.120 -283.950 ;
        RECT 109.415 -284.065 109.635 -283.720 ;
        RECT 108.930 -284.670 109.135 -284.465 ;
        RECT 109.440 -284.490 109.610 -284.065 ;
        RECT 109.930 -284.425 110.100 -283.950 ;
        RECT 110.395 -284.065 110.615 -283.720 ;
        RECT 109.920 -284.670 110.125 -284.425 ;
        RECT 110.420 -284.490 110.590 -284.065 ;
        RECT 110.910 -284.425 111.080 -283.950 ;
        RECT 111.380 -284.010 111.600 -283.720 ;
        RECT 110.890 -284.670 111.095 -284.425 ;
        RECT 111.400 -284.490 111.570 -284.010 ;
        RECT 111.845 -284.420 112.075 -283.810 ;
        RECT 113.585 -283.945 121.040 -283.605 ;
        RECT 121.935 -283.720 125.100 -283.550 ;
        RECT 111.845 -284.470 112.080 -284.420 ;
        RECT 111.875 -284.635 112.080 -284.470 ;
        RECT 111.875 -284.670 112.085 -284.635 ;
        RECT 108.930 -284.840 112.085 -284.670 ;
        RECT 113.630 -284.740 113.800 -283.945 ;
        RECT 114.120 -284.660 114.290 -284.200 ;
        RECT 111.210 -284.950 112.085 -284.840 ;
        RECT 113.070 -284.950 113.910 -284.910 ;
        RECT 108.430 -285.405 109.290 -285.035 ;
        RECT 111.210 -285.235 113.910 -284.950 ;
        RECT 105.405 -286.640 105.575 -286.620 ;
        RECT 106.385 -286.640 106.555 -285.680 ;
        RECT 107.365 -286.640 107.535 -285.680 ;
        RECT 107.840 -286.275 108.210 -285.435 ;
        RECT 108.430 -286.140 108.665 -285.405 ;
        RECT 111.210 -285.675 112.085 -285.235 ;
        RECT 113.070 -285.280 113.910 -285.235 ;
        RECT 114.090 -285.125 114.320 -284.660 ;
        RECT 114.610 -284.740 114.780 -283.945 ;
        RECT 115.100 -284.660 115.270 -284.200 ;
        RECT 115.070 -285.125 115.300 -284.660 ;
        RECT 115.590 -284.740 115.760 -283.945 ;
        RECT 116.080 -284.660 116.250 -284.200 ;
        RECT 116.050 -284.965 116.280 -284.660 ;
        RECT 116.050 -285.020 116.430 -284.965 ;
        RECT 116.680 -285.020 116.980 -284.445 ;
        RECT 118.415 -284.740 118.585 -283.945 ;
        RECT 118.905 -284.660 119.075 -284.200 ;
        RECT 116.050 -285.125 117.005 -285.020 ;
        RECT 114.090 -285.245 117.005 -285.125 ;
        RECT 108.945 -285.845 112.085 -285.675 ;
        RECT 108.945 -286.105 109.125 -285.845 ;
        RECT 109.935 -286.025 110.115 -285.845 ;
        RECT 108.460 -286.510 108.630 -286.140 ;
        RECT 108.455 -286.735 108.635 -286.510 ;
        RECT 108.950 -286.565 109.120 -286.105 ;
        RECT 109.440 -286.460 109.610 -286.025 ;
        RECT 109.930 -286.115 110.115 -286.025 ;
        RECT 109.435 -286.735 109.645 -286.460 ;
        RECT 109.930 -286.565 110.100 -286.115 ;
        RECT 110.420 -286.455 110.590 -286.025 ;
        RECT 110.905 -286.115 111.085 -285.845 ;
        RECT 110.405 -286.735 110.615 -286.455 ;
        RECT 110.910 -286.565 111.080 -286.115 ;
        RECT 111.400 -286.480 111.570 -286.025 ;
        RECT 111.875 -286.065 112.085 -285.845 ;
        RECT 114.090 -285.315 116.430 -285.245 ;
        RECT 114.090 -285.355 116.280 -285.315 ;
        RECT 111.385 -286.735 111.595 -286.480 ;
        RECT 111.890 -286.565 112.060 -286.065 ;
        RECT 114.090 -286.620 114.320 -285.355 ;
        RECT 115.070 -285.680 115.300 -285.355 ;
        RECT 116.050 -285.680 116.280 -285.355 ;
        RECT 114.120 -286.640 114.290 -286.620 ;
        RECT 115.100 -286.640 115.270 -285.680 ;
        RECT 116.080 -286.640 116.250 -285.680 ;
        RECT 116.780 -285.915 117.005 -285.245 ;
        RECT 118.875 -285.125 119.105 -284.660 ;
        RECT 119.395 -284.740 119.565 -283.945 ;
        RECT 119.885 -284.660 120.055 -284.200 ;
        RECT 119.855 -285.125 120.085 -284.660 ;
        RECT 120.375 -284.740 120.545 -283.945 ;
        RECT 121.935 -284.010 122.155 -283.720 ;
        RECT 120.865 -284.660 121.035 -284.200 ;
        RECT 121.960 -284.360 122.130 -284.010 ;
        RECT 120.835 -284.965 121.065 -284.660 ;
        RECT 120.835 -285.125 121.705 -284.965 ;
        RECT 118.875 -285.315 121.705 -285.125 ;
        RECT 118.875 -285.355 121.065 -285.315 ;
        RECT 117.800 -285.915 118.085 -285.710 ;
        RECT 116.780 -286.140 118.085 -285.915 ;
        RECT 117.800 -286.530 118.085 -286.140 ;
        RECT 118.875 -286.620 119.105 -285.355 ;
        RECT 119.855 -285.680 120.085 -285.355 ;
        RECT 120.835 -285.680 121.065 -285.355 ;
        RECT 121.340 -285.435 121.705 -285.315 ;
        RECT 121.930 -285.035 122.165 -284.360 ;
        RECT 122.450 -284.465 122.620 -283.950 ;
        RECT 122.915 -284.065 123.135 -283.720 ;
        RECT 122.430 -284.670 122.635 -284.465 ;
        RECT 122.940 -284.490 123.110 -284.065 ;
        RECT 123.430 -284.425 123.600 -283.950 ;
        RECT 123.895 -284.065 124.115 -283.720 ;
        RECT 123.420 -284.670 123.625 -284.425 ;
        RECT 123.920 -284.490 124.090 -284.065 ;
        RECT 124.410 -284.425 124.580 -283.950 ;
        RECT 124.880 -284.010 125.100 -283.720 ;
        RECT 127.085 -283.945 129.755 -283.605 ;
        RECT 124.390 -284.670 124.595 -284.425 ;
        RECT 124.900 -284.490 125.070 -284.010 ;
        RECT 125.390 -284.420 125.560 -283.950 ;
        RECT 125.375 -284.635 125.580 -284.420 ;
        RECT 125.375 -284.670 125.585 -284.635 ;
        RECT 122.430 -284.840 125.585 -284.670 ;
        RECT 127.130 -284.740 127.300 -283.945 ;
        RECT 127.620 -284.660 127.790 -284.200 ;
        RECT 124.710 -284.985 125.585 -284.840 ;
        RECT 126.570 -284.985 127.410 -284.910 ;
        RECT 121.930 -285.405 122.790 -285.035 ;
        RECT 124.710 -285.250 127.410 -284.985 ;
        RECT 118.905 -286.640 119.075 -286.620 ;
        RECT 119.885 -286.640 120.055 -285.680 ;
        RECT 120.865 -286.640 121.035 -285.680 ;
        RECT 121.340 -286.275 121.710 -285.435 ;
        RECT 121.930 -286.140 122.165 -285.405 ;
        RECT 124.710 -285.675 125.585 -285.250 ;
        RECT 126.570 -285.280 127.410 -285.250 ;
        RECT 127.590 -285.125 127.820 -284.660 ;
        RECT 128.110 -284.740 128.280 -283.945 ;
        RECT 128.600 -284.660 128.770 -284.200 ;
        RECT 128.570 -285.125 128.800 -284.660 ;
        RECT 129.090 -284.740 129.260 -283.945 ;
        RECT 129.580 -284.660 129.750 -284.200 ;
        RECT 129.550 -284.965 129.780 -284.660 ;
        RECT 129.550 -285.075 129.930 -284.965 ;
        RECT 130.105 -285.075 130.345 -283.285 ;
        RECT 142.155 -283.610 142.325 -281.890 ;
        RECT 143.135 -283.610 143.305 -281.890 ;
        RECT 145.200 -282.425 145.370 -281.885 ;
        RECT 146.180 -282.425 146.350 -281.885 ;
        RECT 144.610 -282.660 144.975 -282.595 ;
        RECT 144.110 -282.800 144.975 -282.660 ;
        RECT 144.000 -282.865 144.975 -282.800 ;
        RECT 144.000 -283.610 144.305 -282.865 ;
        RECT 144.610 -282.895 144.975 -282.865 ;
        RECT 147.160 -282.745 147.330 -281.885 ;
        RECT 142.155 -283.760 144.305 -283.610 ;
        RECT 142.155 -283.800 144.250 -283.760 ;
        RECT 145.200 -283.820 145.370 -283.040 ;
        RECT 145.690 -283.580 145.860 -283.040 ;
        RECT 146.180 -283.820 146.350 -283.040 ;
        RECT 146.670 -283.580 146.840 -283.040 ;
        RECT 147.160 -283.095 148.550 -282.745 ;
        RECT 140.375 -284.165 141.510 -284.155 ;
        RECT 143.565 -284.165 143.935 -284.035 ;
        RECT 140.375 -284.355 143.935 -284.165 ;
        RECT 144.500 -284.250 147.575 -283.820 ;
        RECT 129.550 -285.125 130.345 -285.075 ;
        RECT 127.590 -285.260 130.345 -285.125 ;
        RECT 127.590 -285.270 130.340 -285.260 ;
        RECT 122.445 -285.845 125.585 -285.675 ;
        RECT 122.445 -286.105 122.625 -285.845 ;
        RECT 123.435 -286.025 123.615 -285.845 ;
        RECT 121.960 -286.510 122.130 -286.140 ;
        RECT 108.455 -286.905 111.595 -286.735 ;
        RECT 121.955 -286.735 122.135 -286.510 ;
        RECT 122.450 -286.565 122.620 -286.105 ;
        RECT 122.940 -286.460 123.110 -286.025 ;
        RECT 123.430 -286.115 123.615 -286.025 ;
        RECT 122.935 -286.735 123.145 -286.460 ;
        RECT 123.430 -286.565 123.600 -286.115 ;
        RECT 123.920 -286.455 124.090 -286.025 ;
        RECT 124.405 -286.115 124.585 -285.845 ;
        RECT 123.905 -286.735 124.115 -286.455 ;
        RECT 124.410 -286.565 124.580 -286.115 ;
        RECT 124.900 -286.480 125.070 -286.025 ;
        RECT 125.375 -286.065 125.585 -285.845 ;
        RECT 127.590 -285.315 129.930 -285.270 ;
        RECT 127.590 -285.355 129.780 -285.315 ;
        RECT 124.885 -286.735 125.095 -286.480 ;
        RECT 125.390 -286.565 125.560 -286.065 ;
        RECT 127.590 -286.620 127.820 -285.355 ;
        RECT 128.570 -285.680 128.800 -285.355 ;
        RECT 129.550 -285.680 129.780 -285.355 ;
        RECT 127.620 -286.640 127.790 -286.620 ;
        RECT 128.600 -286.640 128.770 -285.680 ;
        RECT 129.580 -286.640 129.750 -285.680 ;
        RECT 121.955 -286.905 125.095 -286.735 ;
        RECT 110.620 -288.410 111.420 -287.750 ;
        RECT 110.655 -289.325 111.330 -288.410 ;
        RECT 115.410 -289.020 130.030 -288.535 ;
        RECT 110.605 -289.985 111.405 -289.325 ;
        RECT 113.220 -291.580 113.390 -289.360 ;
        RECT 114.200 -291.580 114.370 -289.360 ;
        RECT 113.220 -291.585 114.370 -291.580 ;
        RECT 110.090 -291.650 110.750 -291.600 ;
        RECT 112.305 -291.645 112.980 -291.615 ;
        RECT 112.205 -291.650 112.980 -291.645 ;
        RECT 110.090 -291.830 112.980 -291.650 ;
        RECT 113.220 -291.770 114.440 -291.585 ;
        RECT 110.090 -291.900 110.750 -291.830 ;
        RECT 112.205 -291.845 112.980 -291.830 ;
        RECT 112.305 -291.885 112.980 -291.845 ;
        RECT 114.270 -291.945 114.440 -291.770 ;
        RECT 114.920 -291.945 115.220 -291.645 ;
        RECT 102.945 -292.310 110.925 -292.095 ;
        RECT 93.700 -292.420 110.925 -292.310 ;
        RECT 111.855 -292.110 112.650 -292.105 ;
        RECT 111.855 -292.135 112.655 -292.110 ;
        RECT 113.395 -292.135 114.070 -292.105 ;
        RECT 111.855 -292.330 114.070 -292.135 ;
        RECT 111.855 -292.335 112.925 -292.330 ;
        RECT 111.855 -292.400 112.655 -292.335 ;
        RECT 113.395 -292.375 114.070 -292.330 ;
        RECT 114.270 -292.250 115.220 -291.945 ;
        RECT 111.855 -292.405 112.650 -292.400 ;
        RECT 93.700 -292.755 103.845 -292.420 ;
        RECT 50.840 -293.025 51.135 -292.990 ;
        RECT 50.840 -293.440 70.720 -293.025 ;
        RECT 50.840 -293.465 51.135 -293.440 ;
        RECT 40.230 -294.090 43.975 -294.045 ;
        RECT 34.810 -294.355 43.975 -294.090 ;
        RECT 30.860 -296.315 32.095 -296.310 ;
        RECT 32.905 -296.315 33.075 -294.460 ;
        RECT 34.810 -294.970 35.005 -294.355 ;
        RECT 40.815 -294.525 43.975 -294.355 ;
        RECT 35.320 -294.725 40.360 -294.545 ;
        RECT 34.830 -295.915 35.000 -294.970 ;
        RECT 28.830 -296.485 29.995 -296.315 ;
        RECT 30.860 -296.485 33.075 -296.315 ;
        RECT 34.820 -296.330 35.005 -295.915 ;
        RECT 35.320 -295.950 35.490 -294.725 ;
        RECT 36.900 -295.920 37.070 -294.910 ;
        RECT 37.390 -295.905 37.560 -294.910 ;
        RECT 38.710 -295.905 38.880 -294.910 ;
        RECT 36.885 -296.025 37.070 -295.920 ;
        RECT 36.290 -296.210 37.070 -296.025 ;
        RECT 37.380 -296.100 38.880 -295.905 ;
        RECT 36.290 -296.330 36.475 -296.210 ;
        RECT 27.110 -296.755 27.785 -296.720 ;
        RECT 29.810 -296.755 29.995 -296.485 ;
        RECT 34.820 -296.515 36.475 -296.330 ;
        RECT 39.200 -296.365 39.370 -294.910 ;
        RECT 40.180 -294.995 40.360 -294.725 ;
        RECT 40.180 -295.950 40.350 -294.995 ;
        RECT 40.670 -296.365 40.840 -294.910 ;
        RECT 41.730 -295.865 41.900 -294.910 ;
        RECT 42.195 -294.945 42.410 -294.525 ;
        RECT 41.705 -296.090 41.920 -295.865 ;
        RECT 42.220 -295.950 42.390 -294.945 ;
        RECT 43.275 -295.855 43.445 -294.910 ;
        RECT 43.740 -294.955 43.955 -294.525 ;
        RECT 41.225 -296.320 41.920 -296.090 ;
        RECT 38.035 -296.535 40.840 -296.365 ;
        RECT 27.110 -296.940 29.995 -296.755 ;
        RECT 27.110 -296.990 27.785 -296.940 ;
        RECT 29.810 -297.630 29.995 -296.940 ;
        RECT 30.165 -296.765 30.840 -296.730 ;
        RECT 30.165 -296.935 34.260 -296.765 ;
        RECT 38.035 -296.845 38.205 -296.535 ;
        RECT 30.165 -297.000 30.840 -296.935 ;
        RECT 31.105 -297.155 31.780 -297.120 ;
        RECT 31.105 -297.345 33.910 -297.155 ;
        RECT 31.105 -297.390 31.780 -297.345 ;
        RECT 32.780 -297.575 33.460 -297.530 ;
        RECT 29.810 -297.815 32.585 -297.630 ;
        RECT 32.780 -297.760 33.555 -297.575 ;
        RECT 32.785 -297.800 33.460 -297.760 ;
        RECT 30.455 -299.035 30.625 -297.815 ;
        RECT 31.435 -299.035 31.605 -297.815 ;
        RECT 32.415 -299.035 32.585 -297.815 ;
        RECT -4.590 -304.680 17.670 -304.500 ;
        RECT 17.980 -304.280 25.490 -304.110 ;
        RECT 33.740 -304.190 33.910 -297.345 ;
        RECT -4.590 -304.920 -4.345 -304.680 ;
        RECT 7.460 -304.900 8.140 -304.855 ;
        RECT 17.980 -304.900 18.150 -304.280 ;
        RECT 32.210 -304.360 33.910 -304.190 ;
        RECT 18.375 -304.555 19.055 -304.540 ;
        RECT 32.210 -304.555 32.380 -304.360 ;
        RECT 18.375 -304.725 32.380 -304.555 ;
        RECT 32.900 -304.650 33.580 -304.620 ;
        RECT 34.090 -304.650 34.260 -296.935 ;
        RECT 34.825 -297.190 35.520 -296.920 ;
        RECT 37.475 -297.015 38.205 -296.845 ;
        RECT 37.475 -297.590 37.645 -297.015 ;
        RECT 38.570 -297.040 39.265 -296.770 ;
        RECT 34.575 -297.760 37.645 -297.590 ;
        RECT 37.950 -297.395 40.350 -297.225 ;
        RECT 34.830 -299.500 35.000 -297.940 ;
        RECT 35.320 -298.980 35.490 -297.760 ;
        RECT 35.810 -299.500 35.980 -297.940 ;
        RECT 36.410 -299.155 36.580 -297.940 ;
        RECT 36.900 -298.980 37.070 -297.760 ;
        RECT 37.390 -299.155 37.560 -297.940 ;
        RECT 37.950 -299.155 38.120 -297.395 ;
        RECT 36.410 -299.325 38.120 -299.155 ;
        RECT 38.300 -297.765 39.370 -297.595 ;
        RECT 38.300 -299.500 38.470 -297.765 ;
        RECT 39.200 -298.980 39.370 -297.765 ;
        RECT 40.180 -298.980 40.350 -297.395 ;
        RECT 40.615 -297.410 41.310 -297.140 ;
        RECT 41.705 -298.015 41.920 -296.320 ;
        RECT 43.255 -296.810 43.470 -295.855 ;
        RECT 43.765 -295.950 43.935 -294.955 ;
        RECT 44.720 -295.260 50.495 -293.955 ;
        RECT 67.405 -294.385 68.830 -294.095 ;
        RECT 70.305 -294.385 70.720 -293.440 ;
        RECT 94.345 -293.515 94.565 -292.755 ;
        RECT 94.365 -294.310 94.535 -293.515 ;
        RECT 94.855 -294.265 95.025 -293.270 ;
        RECT 95.315 -293.510 95.535 -292.755 ;
        RECT 67.405 -294.525 92.205 -294.385 ;
        RECT 93.895 -294.525 94.625 -294.485 ;
        RECT 67.405 -294.705 94.625 -294.525 ;
        RECT 94.830 -294.510 95.055 -294.265 ;
        RECT 95.345 -294.310 95.515 -293.510 ;
        RECT 99.075 -293.515 99.295 -292.755 ;
        RECT 99.095 -294.310 99.265 -293.515 ;
        RECT 99.585 -294.265 99.755 -293.270 ;
        RECT 100.045 -293.510 100.265 -292.755 ;
        RECT 94.830 -294.515 96.800 -294.510 ;
        RECT 94.830 -294.690 97.045 -294.515 ;
        RECT 98.625 -294.525 99.355 -294.485 ;
        RECT 67.405 -294.855 92.205 -294.705 ;
        RECT 93.895 -294.785 94.625 -294.705 ;
        RECT 96.105 -294.735 97.045 -294.690 ;
        RECT 98.330 -294.705 99.355 -294.525 ;
        RECT 99.560 -294.510 99.785 -294.265 ;
        RECT 100.075 -294.310 100.245 -293.510 ;
        RECT 99.560 -294.690 102.910 -294.510 ;
        RECT 96.385 -294.815 97.045 -294.735 ;
        RECT 98.625 -294.785 99.355 -294.705 ;
        RECT 100.835 -294.735 102.910 -294.690 ;
        RECT 67.405 -295.190 68.830 -294.855 ;
        RECT 95.010 -294.970 95.725 -294.885 ;
        RECT 92.720 -295.150 95.725 -294.970 ;
        RECT 42.755 -297.040 43.470 -296.810 ;
        RECT 41.730 -298.980 41.900 -298.015 ;
        RECT 43.255 -298.025 43.470 -297.040 ;
        RECT 43.690 -297.380 44.385 -297.110 ;
        RECT 43.275 -298.980 43.445 -298.025 ;
        RECT 34.830 -299.670 38.470 -299.500 ;
        RECT 18.375 -304.770 19.055 -304.725 ;
        RECT 32.900 -304.820 34.260 -304.650 ;
        RECT 32.900 -304.850 33.580 -304.820 ;
        RECT -5.025 -305.150 -4.345 -304.920 ;
        RECT 7.295 -305.070 18.150 -304.900 ;
        RECT 7.460 -305.085 8.140 -305.070 ;
        RECT 44.720 -305.235 46.025 -295.260 ;
        RECT 49.190 -299.230 50.495 -295.260 ;
        RECT 92.720 -295.415 92.900 -295.150 ;
        RECT 95.010 -295.185 95.725 -295.150 ;
        RECT 72.315 -296.225 92.900 -295.415 ;
        RECT 94.360 -295.560 96.100 -295.380 ;
        RECT 94.360 -295.755 94.540 -295.560 ;
        RECT 51.605 -297.040 51.950 -296.950 ;
        RECT 77.670 -297.040 78.225 -296.225 ;
        RECT 51.605 -297.595 78.225 -297.040 ;
        RECT 51.605 -297.645 51.950 -297.595 ;
        RECT 94.365 -297.770 94.535 -295.755 ;
        RECT 95.420 -297.630 95.590 -295.730 ;
        RECT 95.875 -295.780 96.100 -295.560 ;
        RECT 95.385 -297.950 95.615 -297.630 ;
        RECT 95.910 -297.770 96.080 -295.780 ;
        RECT 96.385 -295.960 96.635 -294.815 ;
        RECT 99.740 -294.970 100.455 -294.885 ;
        RECT 98.325 -295.150 100.455 -294.970 ;
        RECT 99.740 -295.185 100.455 -295.150 ;
        RECT 99.090 -295.560 100.830 -295.380 ;
        RECT 99.090 -295.755 99.270 -295.560 ;
        RECT 96.400 -297.630 96.570 -295.960 ;
        RECT 96.375 -297.950 96.605 -297.630 ;
        RECT 99.095 -297.770 99.265 -295.755 ;
        RECT 100.150 -297.630 100.320 -295.730 ;
        RECT 100.605 -295.780 100.830 -295.560 ;
        RECT 95.385 -298.140 96.605 -297.950 ;
        RECT 100.115 -297.950 100.345 -297.630 ;
        RECT 100.640 -297.770 100.810 -295.780 ;
        RECT 101.115 -295.960 101.365 -294.735 ;
        RECT 101.130 -297.630 101.300 -295.960 ;
        RECT 101.565 -296.060 101.865 -295.230 ;
        RECT 102.740 -295.670 102.910 -294.735 ;
        RECT 103.185 -295.220 103.355 -293.365 ;
        RECT 103.675 -294.905 103.845 -292.755 ;
        RECT 104.735 -292.870 106.940 -292.700 ;
        RECT 104.735 -292.885 105.890 -292.870 ;
        RECT 104.165 -295.215 104.335 -293.365 ;
        RECT 104.735 -293.405 104.910 -292.885 ;
        RECT 104.735 -294.900 104.905 -293.405 ;
        RECT 105.225 -294.900 105.395 -293.360 ;
        RECT 105.715 -293.415 105.890 -292.885 ;
        RECT 105.715 -294.900 105.885 -293.415 ;
        RECT 105.225 -295.215 105.400 -294.900 ;
        RECT 104.165 -295.220 105.400 -295.215 ;
        RECT 106.280 -295.220 106.450 -293.360 ;
        RECT 106.770 -294.900 106.940 -292.870 ;
        RECT 107.260 -295.220 107.430 -293.360 ;
        RECT 108.835 -294.400 109.005 -292.420 ;
        RECT 109.345 -292.500 110.925 -292.420 ;
        RECT 109.345 -292.675 110.920 -292.500 ;
        RECT 103.185 -295.390 105.400 -295.220 ;
        RECT 106.265 -295.390 107.430 -295.220 ;
        RECT 109.325 -295.325 109.495 -293.360 ;
        RECT 110.515 -294.205 110.920 -292.675 ;
        RECT 112.730 -294.190 112.900 -292.630 ;
        RECT 113.220 -293.770 113.390 -292.630 ;
        RECT 113.780 -293.770 113.950 -292.630 ;
        RECT 114.270 -293.670 114.440 -292.250 ;
        RECT 114.920 -292.315 115.220 -292.250 ;
        RECT 113.220 -293.945 113.950 -293.770 ;
        RECT 112.565 -294.205 114.960 -294.190 ;
        RECT 115.410 -294.205 115.760 -289.020 ;
        RECT 110.515 -294.995 115.760 -294.205 ;
        RECT 112.435 -295.210 115.760 -294.995 ;
        RECT 116.045 -293.415 116.395 -289.745 ;
        RECT 116.880 -293.125 117.050 -289.020 ;
        RECT 117.370 -293.405 117.540 -289.585 ;
        RECT 118.880 -293.125 119.050 -289.020 ;
        RECT 118.530 -293.405 119.200 -293.340 ;
        RECT 116.045 -293.685 117.190 -293.415 ;
        RECT 117.370 -293.575 119.200 -293.405 ;
        RECT 105.420 -295.670 106.095 -295.635 ;
        RECT 102.715 -295.840 106.095 -295.670 ;
        RECT 105.420 -295.905 106.095 -295.840 ;
        RECT 106.265 -295.660 106.450 -295.390 ;
        RECT 109.325 -295.505 110.710 -295.325 ;
        RECT 108.475 -295.660 109.150 -295.625 ;
        RECT 106.265 -295.845 109.150 -295.660 ;
        RECT 104.480 -296.060 105.155 -296.025 ;
        RECT 101.565 -296.250 105.155 -296.060 ;
        RECT 104.480 -296.295 105.155 -296.250 ;
        RECT 102.800 -296.480 103.475 -296.435 ;
        RECT 102.140 -296.655 103.475 -296.480 ;
        RECT 106.265 -296.535 106.450 -295.845 ;
        RECT 108.475 -295.895 109.150 -295.845 ;
        RECT 102.140 -297.140 102.440 -296.655 ;
        RECT 102.705 -296.665 103.475 -296.655 ;
        RECT 102.800 -296.705 103.475 -296.665 ;
        RECT 103.675 -296.720 106.450 -296.535 ;
        RECT 101.105 -297.950 101.335 -297.630 ;
        RECT 103.675 -297.940 103.845 -296.720 ;
        RECT 104.655 -297.940 104.825 -296.720 ;
        RECT 105.635 -297.940 105.805 -296.720 ;
        RECT 109.325 -297.940 109.495 -295.505 ;
        RECT 110.055 -295.625 110.710 -295.505 ;
        RECT 112.480 -296.005 112.650 -295.210 ;
        RECT 112.970 -295.925 113.140 -295.465 ;
        RECT 111.920 -296.545 112.760 -296.175 ;
        RECT 112.940 -296.390 113.170 -295.925 ;
        RECT 113.460 -296.005 113.630 -295.210 ;
        RECT 113.950 -295.925 114.120 -295.465 ;
        RECT 113.920 -296.390 114.150 -295.925 ;
        RECT 114.440 -296.005 114.610 -295.210 ;
        RECT 114.930 -295.925 115.100 -295.465 ;
        RECT 114.900 -296.230 115.130 -295.925 ;
        RECT 116.045 -296.230 116.395 -293.685 ;
        RECT 114.900 -296.390 116.395 -296.230 ;
        RECT 112.940 -296.580 116.395 -296.390 ;
        RECT 112.940 -296.620 115.130 -296.580 ;
        RECT 112.940 -297.885 113.170 -296.620 ;
        RECT 113.920 -296.945 114.150 -296.620 ;
        RECT 114.900 -296.945 115.130 -296.620 ;
        RECT 112.970 -297.905 113.140 -297.885 ;
        RECT 113.950 -297.905 114.120 -296.945 ;
        RECT 114.930 -297.905 115.100 -296.945 ;
        RECT 117.370 -297.550 117.540 -293.575 ;
        RECT 118.530 -293.610 119.200 -293.575 ;
        RECT 119.370 -293.355 119.540 -289.585 ;
        RECT 119.910 -293.355 120.500 -293.295 ;
        RECT 119.370 -293.525 120.500 -293.355 ;
        RECT 119.370 -297.550 119.540 -293.525 ;
        RECT 119.910 -293.585 120.500 -293.525 ;
        RECT 121.265 -293.405 121.615 -292.500 ;
        RECT 121.880 -293.125 122.050 -289.020 ;
        RECT 121.265 -293.675 122.135 -293.405 ;
        RECT 122.370 -293.455 122.540 -289.585 ;
        RECT 123.880 -293.125 124.050 -289.020 ;
        RECT 123.530 -293.455 124.200 -293.415 ;
        RECT 122.370 -293.650 124.200 -293.455 ;
        RECT 122.370 -297.550 122.540 -293.650 ;
        RECT 123.530 -293.685 124.200 -293.650 ;
        RECT 124.370 -293.490 124.540 -289.585 ;
        RECT 125.295 -293.490 125.885 -293.430 ;
        RECT 124.370 -293.660 125.885 -293.490 ;
        RECT 124.370 -297.550 124.540 -293.660 ;
        RECT 125.295 -293.720 125.885 -293.660 ;
        RECT 126.220 -293.440 126.570 -292.505 ;
        RECT 126.880 -293.125 127.050 -289.020 ;
        RECT 126.220 -293.710 127.135 -293.440 ;
        RECT 127.370 -293.460 127.540 -289.585 ;
        RECT 128.880 -293.125 129.050 -289.020 ;
        RECT 129.370 -293.410 129.540 -289.585 ;
        RECT 140.430 -289.715 140.810 -284.355 ;
        RECT 141.505 -284.360 143.935 -284.355 ;
        RECT 141.505 -284.365 141.860 -284.360 ;
        RECT 143.565 -284.390 143.935 -284.360 ;
        RECT 141.665 -286.115 141.835 -284.575 ;
        RECT 142.155 -286.115 142.325 -284.575 ;
        RECT 142.645 -286.115 142.815 -284.575 ;
        RECT 143.135 -286.115 143.305 -284.575 ;
        RECT 143.625 -286.115 143.795 -284.575 ;
        RECT 142.150 -286.375 142.325 -286.115 ;
        RECT 145.720 -286.285 146.025 -284.250 ;
        RECT 148.170 -285.070 148.520 -283.095 ;
        RECT 149.390 -284.365 149.560 -281.445 ;
        RECT 150.425 -281.485 150.635 -281.275 ;
        RECT 149.370 -284.660 149.580 -284.365 ;
        RECT 150.445 -284.395 150.615 -281.485 ;
        RECT 150.935 -284.385 151.105 -281.445 ;
        RECT 151.415 -281.495 151.625 -281.275 ;
        RECT 150.430 -284.660 150.640 -284.395 ;
        RECT 149.370 -284.840 150.640 -284.660 ;
        RECT 150.915 -284.655 151.125 -284.385 ;
        RECT 151.425 -284.485 151.595 -281.495 ;
        RECT 152.485 -284.415 152.655 -281.445 ;
        RECT 150.915 -284.850 151.620 -284.655 ;
        RECT 151.405 -284.910 151.620 -284.850 ;
        RECT 150.195 -285.070 150.970 -285.020 ;
        RECT 148.170 -285.250 150.970 -285.070 ;
        RECT 148.170 -285.260 148.520 -285.250 ;
        RECT 150.195 -285.295 150.970 -285.250 ;
        RECT 151.405 -285.185 152.310 -284.910 ;
        RECT 151.405 -285.535 151.620 -285.185 ;
        RECT 148.845 -285.605 149.620 -285.560 ;
        RECT 148.660 -285.775 149.620 -285.605 ;
        RECT 148.845 -285.835 149.620 -285.775 ;
        RECT 149.850 -285.735 151.620 -285.535 ;
        RECT 152.480 -285.635 152.695 -284.415 ;
        RECT 153.665 -284.760 154.015 -278.075 ;
        RECT 184.485 -278.340 184.655 -277.300 ;
        RECT 185.465 -278.340 185.635 -277.300 ;
        RECT 186.445 -278.340 186.615 -277.300 ;
        RECT 189.350 -278.985 189.520 -277.265 ;
        RECT 190.330 -278.985 190.500 -277.265 ;
        RECT 191.195 -278.010 191.500 -277.265 ;
        RECT 192.395 -277.835 192.565 -277.055 ;
        RECT 192.885 -277.835 193.055 -277.295 ;
        RECT 193.375 -277.835 193.545 -277.055 ;
        RECT 227.340 -277.260 228.575 -277.055 ;
        RECT 232.750 -277.195 233.425 -277.155 ;
        RECT 232.650 -277.205 233.425 -277.195 ;
        RECT 193.865 -277.835 194.035 -277.295 ;
        RECT 227.340 -277.345 227.990 -277.260 ;
        RECT 228.210 -277.325 228.575 -277.260 ;
        RECT 231.615 -277.385 233.425 -277.205 ;
        RECT 236.010 -277.250 239.935 -276.820 ;
        RECT 273.330 -276.885 273.980 -276.425 ;
        RECT 274.790 -276.715 274.960 -275.435 ;
        RECT 275.280 -276.715 275.450 -275.675 ;
        RECT 275.770 -276.715 275.940 -275.435 ;
        RECT 276.260 -276.545 276.430 -275.675 ;
        RECT 279.165 -276.325 279.335 -274.785 ;
        RECT 279.655 -276.325 279.825 -274.785 ;
        RECT 280.145 -276.325 280.315 -274.785 ;
        RECT 280.635 -276.325 280.805 -274.785 ;
        RECT 281.125 -276.325 281.295 -274.785 ;
        RECT 279.005 -276.540 279.360 -276.535 ;
        RECT 281.065 -276.540 281.435 -276.510 ;
        RECT 279.005 -276.545 281.435 -276.540 ;
        RECT 276.260 -276.715 281.435 -276.545 ;
        RECT 283.220 -276.650 283.525 -274.615 ;
        RECT 306.460 -274.765 315.715 -274.010 ;
        RECT 322.120 -273.980 325.445 -273.840 ;
        RECT 322.120 -274.270 327.295 -273.980 ;
        RECT 322.120 -274.675 322.550 -274.270 ;
        RECT 323.420 -274.455 323.595 -274.270 ;
        RECT 325.045 -274.285 327.295 -274.270 ;
        RECT 306.460 -275.105 308.340 -274.765 ;
        RECT 314.465 -275.020 315.715 -274.765 ;
        RECT 317.860 -275.105 322.550 -274.675 ;
        RECT 317.100 -276.555 317.750 -276.095 ;
        RECT 318.560 -276.385 318.730 -275.105 ;
        RECT 319.050 -276.385 319.220 -275.345 ;
        RECT 319.540 -276.385 319.710 -275.105 ;
        RECT 320.030 -276.215 320.200 -275.345 ;
        RECT 322.935 -275.995 323.105 -274.455 ;
        RECT 323.425 -275.995 323.595 -274.455 ;
        RECT 323.915 -275.995 324.085 -274.455 ;
        RECT 324.405 -275.995 324.575 -274.455 ;
        RECT 324.895 -275.995 325.065 -274.455 ;
        RECT 322.775 -276.210 323.130 -276.205 ;
        RECT 324.835 -276.210 325.205 -276.180 ;
        RECT 322.775 -276.215 325.205 -276.210 ;
        RECT 320.030 -276.385 325.205 -276.215 ;
        RECT 326.990 -276.320 327.295 -274.285 ;
        RECT 350.340 -274.040 352.030 -273.560 ;
        RECT 369.220 -273.755 370.920 -271.785 ;
        RECT 396.490 -273.735 397.840 -273.130 ;
        RECT 406.555 -273.735 408.030 -273.525 ;
        RECT 415.900 -273.565 416.955 -271.785 ;
        RECT 360.280 -274.040 361.620 -273.835 ;
        RECT 350.340 -274.695 361.620 -274.040 ;
        RECT 367.885 -273.895 371.210 -273.755 ;
        RECT 367.885 -274.185 373.060 -273.895 ;
        RECT 367.885 -274.590 368.315 -274.185 ;
        RECT 369.185 -274.370 369.360 -274.185 ;
        RECT 370.810 -274.200 373.060 -274.185 ;
        RECT 350.340 -275.015 352.030 -274.695 ;
        RECT 360.280 -275.035 361.620 -274.695 ;
        RECT 363.625 -275.020 368.315 -274.590 ;
        RECT 320.035 -276.405 325.205 -276.385 ;
        RECT 320.035 -276.415 322.780 -276.405 ;
        RECT 317.970 -276.555 318.335 -276.525 ;
        RECT 324.835 -276.535 325.205 -276.405 ;
        RECT 276.265 -276.735 281.435 -276.715 ;
        RECT 276.265 -276.745 279.010 -276.735 ;
        RECT 274.200 -276.885 274.565 -276.855 ;
        RECT 281.065 -276.865 281.435 -276.735 ;
        RECT 273.330 -277.090 274.565 -276.885 ;
        RECT 278.740 -277.025 279.415 -276.985 ;
        RECT 278.640 -277.035 279.415 -277.025 ;
        RECT 273.330 -277.175 273.980 -277.090 ;
        RECT 274.200 -277.155 274.565 -277.090 ;
        RECT 277.605 -277.215 279.415 -277.035 ;
        RECT 282.000 -277.080 285.925 -276.650 ;
        RECT 317.100 -276.760 318.335 -276.555 ;
        RECT 322.510 -276.695 323.185 -276.655 ;
        RECT 322.410 -276.705 323.185 -276.695 ;
        RECT 317.100 -276.845 317.750 -276.760 ;
        RECT 317.970 -276.825 318.335 -276.760 ;
        RECT 321.375 -276.885 323.185 -276.705 ;
        RECT 325.770 -276.750 329.695 -276.320 ;
        RECT 362.865 -276.470 363.515 -276.010 ;
        RECT 364.325 -276.300 364.495 -275.020 ;
        RECT 364.815 -276.300 364.985 -275.260 ;
        RECT 365.305 -276.300 365.475 -275.020 ;
        RECT 365.795 -276.130 365.965 -275.260 ;
        RECT 368.700 -275.910 368.870 -274.370 ;
        RECT 369.190 -275.910 369.360 -274.370 ;
        RECT 369.680 -275.910 369.850 -274.370 ;
        RECT 370.170 -275.910 370.340 -274.370 ;
        RECT 370.660 -275.910 370.830 -274.370 ;
        RECT 368.540 -276.125 368.895 -276.120 ;
        RECT 370.600 -276.125 370.970 -276.095 ;
        RECT 368.540 -276.130 370.970 -276.125 ;
        RECT 365.795 -276.300 370.970 -276.130 ;
        RECT 372.755 -276.235 373.060 -274.200 ;
        RECT 396.490 -274.430 408.030 -273.735 ;
        RECT 414.705 -273.705 418.030 -273.565 ;
        RECT 414.705 -273.995 419.880 -273.705 ;
        RECT 414.705 -274.400 415.135 -273.995 ;
        RECT 416.005 -274.180 416.180 -273.995 ;
        RECT 417.630 -274.010 419.880 -273.995 ;
        RECT 396.490 -274.555 397.840 -274.430 ;
        RECT 406.555 -274.890 408.030 -274.430 ;
        RECT 410.445 -274.830 415.135 -274.400 ;
        RECT 365.800 -276.320 370.970 -276.300 ;
        RECT 365.800 -276.330 368.545 -276.320 ;
        RECT 363.735 -276.470 364.100 -276.440 ;
        RECT 370.600 -276.450 370.970 -276.320 ;
        RECT 362.865 -276.675 364.100 -276.470 ;
        RECT 368.275 -276.610 368.950 -276.570 ;
        RECT 368.175 -276.620 368.950 -276.610 ;
        RECT 322.410 -276.895 323.185 -276.885 ;
        RECT 322.510 -276.925 323.185 -276.895 ;
        RECT 323.425 -276.810 325.520 -276.770 ;
        RECT 323.425 -276.960 325.575 -276.810 ;
        RECT 278.640 -277.225 279.415 -277.215 ;
        RECT 232.650 -277.395 233.425 -277.385 ;
        RECT 232.750 -277.425 233.425 -277.395 ;
        RECT 233.665 -277.310 235.760 -277.270 ;
        RECT 233.665 -277.460 235.815 -277.310 ;
        RECT 191.805 -278.010 192.170 -277.980 ;
        RECT 191.195 -278.075 192.170 -278.010 ;
        RECT 191.305 -278.215 192.170 -278.075 ;
        RECT 191.805 -278.280 192.170 -278.215 ;
        RECT 194.355 -278.130 196.215 -277.780 ;
        RECT 192.395 -278.990 192.565 -278.450 ;
        RECT 193.375 -278.990 193.545 -278.450 ;
        RECT 194.355 -278.990 194.525 -278.130 ;
        RECT 160.245 -280.555 161.850 -280.385 ;
        RECT 159.350 -283.235 159.520 -280.735 ;
        RECT 159.345 -283.465 159.520 -283.235 ;
        RECT 160.245 -283.465 160.445 -280.555 ;
        RECT 160.690 -280.755 160.865 -280.555 ;
        RECT 160.695 -283.275 160.865 -280.755 ;
        RECT 161.185 -283.240 161.355 -280.735 ;
        RECT 161.675 -280.750 161.850 -280.555 ;
        RECT 159.345 -283.665 160.445 -283.465 ;
        RECT 161.170 -283.840 161.360 -283.240 ;
        RECT 161.675 -283.275 161.845 -280.750 ;
        RECT 162.325 -283.655 162.495 -280.735 ;
        RECT 163.955 -283.305 164.125 -280.735 ;
        RECT 165.095 -282.185 165.265 -280.735 ;
        RECT 192.625 -281.330 193.825 -281.160 ;
        RECT 165.090 -282.650 165.275 -282.185 ;
        RECT 165.090 -282.835 165.775 -282.650 ;
        RECT 163.955 -283.475 164.750 -283.305 ;
        RECT 163.070 -283.655 163.760 -283.600 ;
        RECT 159.350 -284.030 161.360 -283.840 ;
        RECT 161.695 -283.825 163.760 -283.655 ;
        RECT 158.165 -284.085 158.855 -284.035 ;
        RECT 156.215 -284.255 158.855 -284.085 ;
        RECT 153.610 -285.120 154.135 -284.760 ;
        RECT 156.215 -285.635 156.430 -284.255 ;
        RECT 158.165 -284.305 158.855 -284.255 ;
        RECT 158.445 -284.760 159.135 -284.715 ;
        RECT 157.395 -284.930 159.135 -284.760 ;
        RECT 157.395 -285.565 157.755 -284.930 ;
        RECT 158.445 -284.985 159.135 -284.930 ;
        RECT 157.395 -285.610 157.815 -285.565 ;
        RECT 143.775 -286.375 146.025 -286.285 ;
        RECT 141.565 -286.590 146.025 -286.375 ;
        RECT 141.565 -286.680 143.810 -286.590 ;
        RECT 145.720 -288.065 146.025 -286.590 ;
        RECT 149.390 -287.475 149.560 -286.005 ;
        RECT 149.850 -286.085 150.075 -285.735 ;
        RECT 151.810 -285.835 156.430 -285.635 ;
        RECT 152.050 -285.850 156.430 -285.835 ;
        RECT 149.355 -288.065 149.590 -287.475 ;
        RECT 149.880 -287.545 150.050 -286.085 ;
        RECT 150.370 -287.470 150.540 -286.005 ;
        RECT 151.580 -287.420 151.750 -286.005 ;
        RECT 152.050 -286.050 152.270 -285.850 ;
        RECT 157.420 -285.960 157.815 -285.610 ;
        RECT 150.335 -288.065 150.570 -287.470 ;
        RECT 151.545 -288.065 151.780 -287.420 ;
        RECT 152.070 -287.545 152.240 -286.050 ;
        RECT 158.860 -287.170 159.030 -285.715 ;
        RECT 158.850 -287.725 159.035 -287.170 ;
        RECT 159.350 -287.255 159.520 -284.030 ;
        RECT 160.495 -284.380 160.685 -284.030 ;
        RECT 161.695 -284.220 161.865 -283.825 ;
        RECT 163.070 -283.870 163.760 -283.825 ;
        RECT 160.445 -285.070 160.715 -284.380 ;
        RECT 161.210 -284.390 161.865 -284.220 ;
        RECT 162.195 -284.305 162.885 -284.035 ;
        RECT 164.120 -284.380 164.390 -283.690 ;
        RECT 164.580 -283.695 164.750 -283.475 ;
        RECT 164.580 -283.965 165.410 -283.695 ;
        RECT 161.210 -287.255 161.380 -284.390 ;
        RECT 164.580 -284.540 164.750 -283.965 ;
        RECT 165.010 -284.540 165.280 -284.455 ;
        RECT 161.700 -284.735 162.495 -284.560 ;
        RECT 164.580 -284.565 165.280 -284.540 ;
        RECT 164.440 -284.710 165.280 -284.565 ;
        RECT 161.700 -287.255 161.870 -284.735 ;
        RECT 162.325 -287.255 162.495 -284.735 ;
        RECT 162.815 -287.170 162.985 -284.715 ;
        RECT 163.465 -287.165 163.635 -284.715 ;
        RECT 156.165 -287.745 159.220 -287.725 ;
        RECT 162.810 -287.745 162.995 -287.170 ;
        RECT 163.450 -287.745 163.635 -287.165 ;
        RECT 163.955 -287.255 164.125 -284.715 ;
        RECT 164.440 -284.735 164.750 -284.710 ;
        RECT 164.445 -287.255 164.615 -284.735 ;
        RECT 165.010 -284.750 165.280 -284.710 ;
        RECT 165.585 -285.300 165.775 -282.835 ;
        RECT 184.355 -283.665 184.525 -281.945 ;
        RECT 185.335 -283.665 185.505 -281.945 ;
        RECT 187.400 -282.480 187.570 -281.940 ;
        RECT 188.380 -282.480 188.550 -281.940 ;
        RECT 186.810 -282.715 187.175 -282.650 ;
        RECT 186.310 -282.855 187.175 -282.715 ;
        RECT 186.200 -282.920 187.175 -282.855 ;
        RECT 186.200 -283.665 186.505 -282.920 ;
        RECT 186.810 -282.950 187.175 -282.920 ;
        RECT 189.360 -282.800 189.530 -281.940 ;
        RECT 184.355 -283.815 186.505 -283.665 ;
        RECT 184.355 -283.855 186.450 -283.815 ;
        RECT 187.400 -283.875 187.570 -283.095 ;
        RECT 187.890 -283.635 188.060 -283.095 ;
        RECT 188.380 -283.875 188.550 -283.095 ;
        RECT 188.870 -283.635 189.040 -283.095 ;
        RECT 189.360 -283.150 190.750 -282.800 ;
        RECT 182.575 -284.220 183.710 -284.210 ;
        RECT 185.765 -284.220 186.135 -284.090 ;
        RECT 182.575 -284.410 186.135 -284.220 ;
        RECT 186.700 -284.305 189.775 -283.875 ;
        RECT 165.585 -285.490 167.045 -285.300 ;
        RECT 165.095 -287.160 165.265 -285.715 ;
        RECT 165.585 -285.740 165.775 -285.490 ;
        RECT 165.085 -287.745 165.270 -287.160 ;
        RECT 165.585 -287.255 165.755 -285.740 ;
        RECT 156.165 -288.065 165.835 -287.745 ;
        RECT 145.720 -288.290 165.835 -288.065 ;
        RECT 145.720 -288.630 156.730 -288.290 ;
        RECT 158.470 -288.550 165.835 -288.290 ;
        RECT 136.450 -289.995 140.810 -289.715 ;
        RECT 166.855 -289.965 167.045 -285.490 ;
        RECT 182.630 -288.660 183.010 -284.410 ;
        RECT 183.705 -284.415 186.135 -284.410 ;
        RECT 183.705 -284.420 184.060 -284.415 ;
        RECT 185.765 -284.445 186.135 -284.415 ;
        RECT 183.865 -286.170 184.035 -284.630 ;
        RECT 184.355 -286.170 184.525 -284.630 ;
        RECT 184.845 -286.170 185.015 -284.630 ;
        RECT 185.335 -286.170 185.505 -284.630 ;
        RECT 185.825 -286.170 185.995 -284.630 ;
        RECT 184.350 -286.430 184.525 -286.170 ;
        RECT 187.920 -286.340 188.225 -284.305 ;
        RECT 190.370 -285.125 190.720 -283.150 ;
        RECT 191.590 -284.420 191.760 -281.500 ;
        RECT 192.625 -281.540 192.835 -281.330 ;
        RECT 191.570 -284.715 191.780 -284.420 ;
        RECT 192.645 -284.450 192.815 -281.540 ;
        RECT 193.135 -284.440 193.305 -281.500 ;
        RECT 193.615 -281.550 193.825 -281.330 ;
        RECT 192.630 -284.715 192.840 -284.450 ;
        RECT 191.570 -284.895 192.840 -284.715 ;
        RECT 193.115 -284.710 193.325 -284.440 ;
        RECT 193.625 -284.540 193.795 -281.550 ;
        RECT 194.685 -284.470 194.855 -281.500 ;
        RECT 193.115 -284.905 193.820 -284.710 ;
        RECT 193.605 -284.965 193.820 -284.905 ;
        RECT 192.395 -285.125 193.170 -285.075 ;
        RECT 190.370 -285.305 193.170 -285.125 ;
        RECT 190.370 -285.315 190.720 -285.305 ;
        RECT 192.395 -285.350 193.170 -285.305 ;
        RECT 193.605 -285.240 194.510 -284.965 ;
        RECT 193.605 -285.590 193.820 -285.240 ;
        RECT 191.045 -285.660 191.820 -285.615 ;
        RECT 190.860 -285.830 191.820 -285.660 ;
        RECT 191.045 -285.890 191.820 -285.830 ;
        RECT 192.050 -285.790 193.820 -285.590 ;
        RECT 194.680 -285.690 194.895 -284.470 ;
        RECT 195.865 -284.815 196.215 -278.130 ;
        RECT 228.800 -278.535 228.970 -277.495 ;
        RECT 229.780 -278.535 229.950 -277.495 ;
        RECT 230.760 -278.535 230.930 -277.495 ;
        RECT 233.665 -279.180 233.835 -277.460 ;
        RECT 234.645 -279.180 234.815 -277.460 ;
        RECT 235.510 -278.205 235.815 -277.460 ;
        RECT 236.710 -278.030 236.880 -277.250 ;
        RECT 237.200 -278.030 237.370 -277.490 ;
        RECT 237.690 -278.030 237.860 -277.250 ;
        RECT 278.740 -277.255 279.415 -277.225 ;
        RECT 279.655 -277.140 281.750 -277.100 ;
        RECT 279.655 -277.290 281.805 -277.140 ;
        RECT 238.180 -278.030 238.350 -277.490 ;
        RECT 236.120 -278.205 236.485 -278.175 ;
        RECT 235.510 -278.270 236.485 -278.205 ;
        RECT 235.620 -278.410 236.485 -278.270 ;
        RECT 236.120 -278.475 236.485 -278.410 ;
        RECT 238.670 -278.325 240.530 -277.975 ;
        RECT 236.710 -279.185 236.880 -278.645 ;
        RECT 237.690 -279.185 237.860 -278.645 ;
        RECT 238.670 -279.185 238.840 -278.325 ;
        RECT 202.445 -280.610 204.050 -280.440 ;
        RECT 201.550 -283.290 201.720 -280.790 ;
        RECT 201.545 -283.520 201.720 -283.290 ;
        RECT 202.445 -283.520 202.645 -280.610 ;
        RECT 202.890 -280.810 203.065 -280.610 ;
        RECT 202.895 -283.330 203.065 -280.810 ;
        RECT 203.385 -283.295 203.555 -280.790 ;
        RECT 203.875 -280.805 204.050 -280.610 ;
        RECT 201.545 -283.720 202.645 -283.520 ;
        RECT 203.370 -283.895 203.560 -283.295 ;
        RECT 203.875 -283.330 204.045 -280.805 ;
        RECT 204.525 -283.710 204.695 -280.790 ;
        RECT 206.155 -283.360 206.325 -280.790 ;
        RECT 207.295 -282.240 207.465 -280.790 ;
        RECT 236.940 -281.525 238.140 -281.355 ;
        RECT 207.290 -282.705 207.475 -282.240 ;
        RECT 207.290 -282.890 207.975 -282.705 ;
        RECT 206.155 -283.530 206.950 -283.360 ;
        RECT 205.270 -283.710 205.960 -283.655 ;
        RECT 201.550 -284.085 203.560 -283.895 ;
        RECT 203.895 -283.880 205.960 -283.710 ;
        RECT 200.365 -284.140 201.055 -284.090 ;
        RECT 198.415 -284.310 201.055 -284.140 ;
        RECT 195.810 -285.175 196.335 -284.815 ;
        RECT 198.415 -285.690 198.630 -284.310 ;
        RECT 200.365 -284.360 201.055 -284.310 ;
        RECT 200.645 -284.815 201.335 -284.770 ;
        RECT 199.595 -284.985 201.335 -284.815 ;
        RECT 199.595 -285.620 199.955 -284.985 ;
        RECT 200.645 -285.040 201.335 -284.985 ;
        RECT 199.595 -285.665 200.015 -285.620 ;
        RECT 185.975 -286.430 188.225 -286.340 ;
        RECT 183.765 -286.645 188.225 -286.430 ;
        RECT 183.765 -286.735 186.010 -286.645 ;
        RECT 136.450 -290.375 156.980 -289.995 ;
        RECT 136.450 -290.445 140.810 -290.375 ;
        RECT 129.775 -293.410 130.365 -293.370 ;
        RECT 128.495 -293.460 129.165 -293.425 ;
        RECT 127.370 -293.655 129.165 -293.460 ;
        RECT 127.370 -297.550 127.540 -293.655 ;
        RECT 128.495 -293.695 129.165 -293.655 ;
        RECT 129.370 -293.580 130.380 -293.410 ;
        RECT 129.370 -297.550 129.540 -293.580 ;
        RECT 129.775 -293.660 130.365 -293.580 ;
        RECT 100.115 -298.140 101.335 -297.950 ;
        RECT 49.190 -300.535 54.040 -299.230 ;
        RECT 49.930 -302.750 50.670 -302.510 ;
        RECT 49.150 -303.425 49.765 -303.205 ;
        RECT -24.235 -305.345 -21.075 -305.300 ;
        RECT -11.735 -305.345 -8.575 -305.300 ;
        RECT 0.765 -305.345 3.925 -305.300 ;
        RECT 13.265 -305.345 16.425 -305.300 ;
        RECT 25.765 -305.345 28.925 -305.300 ;
        RECT 40.685 -305.345 46.025 -305.235 ;
        RECT -30.240 -305.350 -21.075 -305.345 ;
        RECT -17.740 -305.350 46.025 -305.345 ;
        RECT -30.240 -305.610 46.025 -305.350 ;
        RECT -30.240 -306.225 -30.045 -305.610 ;
        RECT -24.235 -305.780 -17.545 -305.610 ;
        RECT -11.735 -305.780 -8.575 -305.610 ;
        RECT -29.730 -305.980 -24.690 -305.800 ;
        RECT -30.220 -307.170 -30.050 -306.225 ;
        RECT -30.230 -307.585 -30.045 -307.170 ;
        RECT -29.730 -307.205 -29.560 -305.980 ;
        RECT -28.150 -307.175 -27.980 -306.165 ;
        RECT -27.660 -307.160 -27.490 -306.165 ;
        RECT -26.340 -307.160 -26.170 -306.165 ;
        RECT -28.165 -307.280 -27.980 -307.175 ;
        RECT -28.760 -307.465 -27.980 -307.280 ;
        RECT -27.670 -307.355 -26.170 -307.160 ;
        RECT -28.760 -307.585 -28.575 -307.465 ;
        RECT -30.230 -307.770 -28.575 -307.585 ;
        RECT -25.850 -307.620 -25.680 -306.165 ;
        RECT -24.870 -306.250 -24.690 -305.980 ;
        RECT -24.870 -307.205 -24.700 -306.250 ;
        RECT -24.380 -307.620 -24.210 -306.165 ;
        RECT -23.320 -307.120 -23.150 -306.165 ;
        RECT -22.855 -306.200 -22.640 -305.780 ;
        RECT -21.680 -305.785 -17.545 -305.780 ;
        RECT -23.345 -307.345 -23.130 -307.120 ;
        RECT -22.830 -307.205 -22.660 -306.200 ;
        RECT -21.775 -307.110 -21.605 -306.165 ;
        RECT -21.310 -306.210 -21.095 -305.785 ;
        RECT -23.825 -307.575 -23.130 -307.345 ;
        RECT -27.015 -307.790 -24.210 -307.620 ;
        RECT -27.015 -308.100 -26.845 -307.790 ;
        RECT -30.225 -308.445 -29.530 -308.175 ;
        RECT -27.575 -308.270 -26.845 -308.100 ;
        RECT -27.575 -308.845 -27.405 -308.270 ;
        RECT -26.480 -308.295 -25.785 -308.025 ;
        RECT -30.775 -309.015 -27.405 -308.845 ;
        RECT -27.100 -308.650 -24.700 -308.480 ;
        RECT -84.330 -309.170 -81.005 -309.030 ;
        RECT -104.225 -309.445 -101.450 -309.260 ;
        RECT -101.250 -309.380 -92.160 -309.205 ;
        RECT -101.250 -309.390 -100.480 -309.380 ;
        RECT -101.250 -309.430 -100.575 -309.390 ;
        RECT -92.450 -309.405 -92.160 -309.380 ;
        RECT -103.580 -310.665 -103.410 -309.445 ;
        RECT -102.600 -310.665 -102.430 -309.445 ;
        RECT -101.620 -310.665 -101.450 -309.445 ;
        RECT -38.725 -309.985 -37.725 -309.865 ;
        RECT -90.630 -310.665 -37.725 -309.985 ;
        RECT -38.725 -310.720 -37.725 -310.665 ;
        RECT -30.220 -310.755 -30.050 -309.195 ;
        RECT -29.730 -310.235 -29.560 -309.015 ;
        RECT -29.240 -310.755 -29.070 -309.195 ;
        RECT -28.640 -310.410 -28.470 -309.195 ;
        RECT -28.150 -310.235 -27.980 -309.015 ;
        RECT -27.660 -310.410 -27.490 -309.195 ;
        RECT -27.100 -310.410 -26.930 -308.650 ;
        RECT -28.640 -310.580 -26.930 -310.410 ;
        RECT -26.750 -309.020 -25.680 -308.850 ;
        RECT -26.750 -310.755 -26.580 -309.020 ;
        RECT -25.850 -310.235 -25.680 -309.020 ;
        RECT -24.870 -310.235 -24.700 -308.650 ;
        RECT -24.435 -308.665 -23.740 -308.395 ;
        RECT -23.345 -309.270 -23.130 -307.575 ;
        RECT -21.795 -308.065 -21.580 -307.110 ;
        RECT -21.285 -307.205 -21.115 -306.210 ;
        RECT -17.740 -306.225 -17.545 -305.785 ;
        RECT -17.230 -305.980 -12.190 -305.800 ;
        RECT -18.590 -307.030 -18.360 -306.350 ;
        RECT -22.295 -308.295 -21.580 -308.065 ;
        RECT -23.320 -310.235 -23.150 -309.270 ;
        RECT -21.795 -309.280 -21.580 -308.295 ;
        RECT -21.360 -308.635 -20.665 -308.365 ;
        RECT -18.560 -308.845 -18.390 -307.030 ;
        RECT -17.720 -307.170 -17.550 -306.225 ;
        RECT -17.730 -307.585 -17.545 -307.170 ;
        RECT -17.230 -307.205 -17.060 -305.980 ;
        RECT -15.650 -307.175 -15.480 -306.165 ;
        RECT -15.160 -307.160 -14.990 -306.165 ;
        RECT -13.840 -307.160 -13.670 -306.165 ;
        RECT -15.665 -307.280 -15.480 -307.175 ;
        RECT -16.260 -307.465 -15.480 -307.280 ;
        RECT -15.170 -307.355 -13.670 -307.160 ;
        RECT -16.260 -307.585 -16.075 -307.465 ;
        RECT -17.730 -307.770 -16.075 -307.585 ;
        RECT -13.350 -307.620 -13.180 -306.165 ;
        RECT -12.370 -306.250 -12.190 -305.980 ;
        RECT -12.370 -307.205 -12.200 -306.250 ;
        RECT -11.880 -307.620 -11.710 -306.165 ;
        RECT -10.820 -307.120 -10.650 -306.165 ;
        RECT -10.355 -306.200 -10.140 -305.780 ;
        RECT -10.845 -307.345 -10.630 -307.120 ;
        RECT -10.330 -307.205 -10.160 -306.200 ;
        RECT -9.275 -307.110 -9.105 -306.165 ;
        RECT -8.810 -306.210 -8.595 -305.780 ;
        RECT -11.325 -307.575 -10.630 -307.345 ;
        RECT -15.815 -307.925 -15.120 -307.655 ;
        RECT -14.515 -307.790 -11.710 -307.620 ;
        RECT -14.515 -308.100 -14.345 -307.790 ;
        RECT -17.725 -308.445 -17.030 -308.175 ;
        RECT -15.075 -308.270 -14.345 -308.100 ;
        RECT -15.075 -308.845 -14.905 -308.270 ;
        RECT -13.980 -308.295 -13.285 -308.025 ;
        RECT -18.560 -309.015 -14.905 -308.845 ;
        RECT -14.600 -308.650 -12.200 -308.480 ;
        RECT -21.775 -310.235 -21.605 -309.280 ;
        RECT -30.220 -310.925 -26.580 -310.755 ;
        RECT -17.720 -310.755 -17.550 -309.195 ;
        RECT -17.230 -310.235 -17.060 -309.015 ;
        RECT -16.740 -310.755 -16.570 -309.195 ;
        RECT -16.140 -310.410 -15.970 -309.195 ;
        RECT -15.650 -310.235 -15.480 -309.015 ;
        RECT -15.160 -310.410 -14.990 -309.195 ;
        RECT -14.600 -310.410 -14.430 -308.650 ;
        RECT -16.140 -310.580 -14.430 -310.410 ;
        RECT -14.250 -309.020 -13.180 -308.850 ;
        RECT -14.250 -310.755 -14.080 -309.020 ;
        RECT -13.350 -310.235 -13.180 -309.020 ;
        RECT -12.370 -310.235 -12.200 -308.650 ;
        RECT -11.935 -308.665 -11.240 -308.395 ;
        RECT -10.845 -309.270 -10.630 -307.575 ;
        RECT -10.425 -307.895 -9.730 -307.625 ;
        RECT -9.295 -308.065 -9.080 -307.110 ;
        RECT -8.785 -307.205 -8.615 -306.210 ;
        RECT -5.240 -306.225 -5.045 -305.610 ;
        RECT 0.765 -305.780 3.925 -305.610 ;
        RECT -4.730 -305.980 0.310 -305.800 ;
        RECT -5.850 -307.010 -5.620 -306.330 ;
        RECT -9.795 -308.295 -9.080 -308.065 ;
        RECT -10.820 -310.235 -10.650 -309.270 ;
        RECT -9.295 -309.280 -9.080 -308.295 ;
        RECT -8.860 -308.635 -8.165 -308.365 ;
        RECT -5.820 -308.845 -5.650 -307.010 ;
        RECT -5.220 -307.170 -5.050 -306.225 ;
        RECT -5.230 -307.585 -5.045 -307.170 ;
        RECT -4.730 -307.205 -4.560 -305.980 ;
        RECT -3.150 -307.175 -2.980 -306.165 ;
        RECT -2.660 -307.160 -2.490 -306.165 ;
        RECT -1.340 -307.160 -1.170 -306.165 ;
        RECT -3.165 -307.280 -2.980 -307.175 ;
        RECT -3.760 -307.465 -2.980 -307.280 ;
        RECT -2.670 -307.355 -1.170 -307.160 ;
        RECT -3.760 -307.585 -3.575 -307.465 ;
        RECT -5.230 -307.770 -3.575 -307.585 ;
        RECT -0.850 -307.620 -0.680 -306.165 ;
        RECT 0.130 -306.250 0.310 -305.980 ;
        RECT 0.130 -307.205 0.300 -306.250 ;
        RECT 0.620 -307.620 0.790 -306.165 ;
        RECT 1.680 -307.120 1.850 -306.165 ;
        RECT 2.145 -306.200 2.360 -305.780 ;
        RECT 1.655 -307.345 1.870 -307.120 ;
        RECT 2.170 -307.205 2.340 -306.200 ;
        RECT 3.225 -307.110 3.395 -306.165 ;
        RECT 3.690 -306.210 3.905 -305.780 ;
        RECT 1.175 -307.575 1.870 -307.345 ;
        RECT -3.315 -307.925 -2.620 -307.655 ;
        RECT -2.015 -307.790 0.790 -307.620 ;
        RECT -2.015 -308.100 -1.845 -307.790 ;
        RECT -5.225 -308.445 -4.530 -308.175 ;
        RECT -2.575 -308.270 -1.845 -308.100 ;
        RECT -2.575 -308.845 -2.405 -308.270 ;
        RECT -1.480 -308.295 -0.785 -308.025 ;
        RECT -5.820 -309.015 -2.405 -308.845 ;
        RECT -2.100 -308.650 0.300 -308.480 ;
        RECT -9.275 -310.235 -9.105 -309.280 ;
        RECT -17.720 -310.925 -14.080 -310.755 ;
        RECT -5.220 -310.755 -5.050 -309.195 ;
        RECT -4.730 -310.235 -4.560 -309.015 ;
        RECT -4.240 -310.755 -4.070 -309.195 ;
        RECT -3.640 -310.410 -3.470 -309.195 ;
        RECT -3.150 -310.235 -2.980 -309.015 ;
        RECT -2.660 -310.410 -2.490 -309.195 ;
        RECT -2.100 -310.410 -1.930 -308.650 ;
        RECT -3.640 -310.580 -1.930 -310.410 ;
        RECT -1.750 -309.020 -0.680 -308.850 ;
        RECT -1.750 -310.755 -1.580 -309.020 ;
        RECT -0.850 -310.235 -0.680 -309.020 ;
        RECT 0.130 -310.235 0.300 -308.650 ;
        RECT 0.565 -308.665 1.260 -308.395 ;
        RECT 1.655 -309.270 1.870 -307.575 ;
        RECT 2.075 -307.895 2.770 -307.625 ;
        RECT 3.205 -308.065 3.420 -307.110 ;
        RECT 3.715 -307.205 3.885 -306.210 ;
        RECT 7.260 -306.225 7.455 -305.610 ;
        RECT 13.265 -305.780 16.425 -305.610 ;
        RECT 7.770 -305.980 12.810 -305.800 ;
        RECT 6.550 -307.010 6.780 -306.330 ;
        RECT 2.705 -308.295 3.420 -308.065 ;
        RECT 1.680 -310.235 1.850 -309.270 ;
        RECT 3.205 -309.280 3.420 -308.295 ;
        RECT 3.640 -308.635 4.335 -308.365 ;
        RECT 6.580 -308.845 6.750 -307.010 ;
        RECT 7.280 -307.170 7.450 -306.225 ;
        RECT 7.270 -307.585 7.455 -307.170 ;
        RECT 7.770 -307.205 7.940 -305.980 ;
        RECT 9.350 -307.175 9.520 -306.165 ;
        RECT 9.840 -307.160 10.010 -306.165 ;
        RECT 11.160 -307.160 11.330 -306.165 ;
        RECT 9.335 -307.280 9.520 -307.175 ;
        RECT 8.740 -307.465 9.520 -307.280 ;
        RECT 9.830 -307.355 11.330 -307.160 ;
        RECT 8.740 -307.585 8.925 -307.465 ;
        RECT 7.270 -307.770 8.925 -307.585 ;
        RECT 11.650 -307.620 11.820 -306.165 ;
        RECT 12.630 -306.250 12.810 -305.980 ;
        RECT 12.630 -307.205 12.800 -306.250 ;
        RECT 13.120 -307.620 13.290 -306.165 ;
        RECT 14.180 -307.120 14.350 -306.165 ;
        RECT 14.645 -306.200 14.860 -305.780 ;
        RECT 14.155 -307.345 14.370 -307.120 ;
        RECT 14.670 -307.205 14.840 -306.200 ;
        RECT 15.725 -307.110 15.895 -306.165 ;
        RECT 16.190 -306.210 16.405 -305.780 ;
        RECT 13.675 -307.575 14.370 -307.345 ;
        RECT 9.185 -307.925 9.880 -307.655 ;
        RECT 10.485 -307.790 13.290 -307.620 ;
        RECT 10.485 -308.100 10.655 -307.790 ;
        RECT 7.275 -308.445 7.970 -308.175 ;
        RECT 9.925 -308.270 10.655 -308.100 ;
        RECT 9.925 -308.845 10.095 -308.270 ;
        RECT 11.020 -308.295 11.715 -308.025 ;
        RECT 6.580 -309.015 10.095 -308.845 ;
        RECT 10.400 -308.650 12.800 -308.480 ;
        RECT 6.580 -309.020 6.750 -309.015 ;
        RECT 3.225 -310.235 3.395 -309.280 ;
        RECT -5.220 -310.925 -1.580 -310.755 ;
        RECT 7.280 -310.755 7.450 -309.195 ;
        RECT 7.770 -310.235 7.940 -309.015 ;
        RECT 8.260 -310.755 8.430 -309.195 ;
        RECT 8.860 -310.410 9.030 -309.195 ;
        RECT 9.350 -310.235 9.520 -309.015 ;
        RECT 9.840 -310.410 10.010 -309.195 ;
        RECT 10.400 -310.410 10.570 -308.650 ;
        RECT 8.860 -310.580 10.570 -310.410 ;
        RECT 10.750 -309.020 11.820 -308.850 ;
        RECT 10.750 -310.755 10.920 -309.020 ;
        RECT 11.650 -310.235 11.820 -309.020 ;
        RECT 12.630 -310.235 12.800 -308.650 ;
        RECT 13.065 -308.665 13.760 -308.395 ;
        RECT 14.155 -309.270 14.370 -307.575 ;
        RECT 14.575 -307.895 15.270 -307.625 ;
        RECT 15.705 -308.065 15.920 -307.110 ;
        RECT 16.215 -307.205 16.385 -306.210 ;
        RECT 19.760 -306.225 19.955 -305.610 ;
        RECT 25.765 -305.780 28.925 -305.610 ;
        RECT 20.270 -305.980 25.310 -305.800 ;
        RECT 18.635 -307.010 18.865 -306.330 ;
        RECT 18.660 -307.015 18.835 -307.010 ;
        RECT 15.205 -308.295 15.920 -308.065 ;
        RECT 14.180 -310.235 14.350 -309.270 ;
        RECT 15.705 -309.280 15.920 -308.295 ;
        RECT 16.140 -308.635 16.835 -308.365 ;
        RECT 18.660 -308.845 18.830 -307.015 ;
        RECT 19.780 -307.170 19.950 -306.225 ;
        RECT 19.770 -307.585 19.955 -307.170 ;
        RECT 20.270 -307.205 20.440 -305.980 ;
        RECT 21.850 -307.175 22.020 -306.165 ;
        RECT 22.340 -307.160 22.510 -306.165 ;
        RECT 23.660 -307.160 23.830 -306.165 ;
        RECT 21.835 -307.280 22.020 -307.175 ;
        RECT 21.240 -307.465 22.020 -307.280 ;
        RECT 22.330 -307.355 23.830 -307.160 ;
        RECT 21.240 -307.585 21.425 -307.465 ;
        RECT 19.770 -307.770 21.425 -307.585 ;
        RECT 24.150 -307.620 24.320 -306.165 ;
        RECT 25.130 -306.250 25.310 -305.980 ;
        RECT 25.130 -307.205 25.300 -306.250 ;
        RECT 25.620 -307.620 25.790 -306.165 ;
        RECT 26.680 -307.120 26.850 -306.165 ;
        RECT 27.145 -306.200 27.360 -305.780 ;
        RECT 26.655 -307.345 26.870 -307.120 ;
        RECT 27.170 -307.205 27.340 -306.200 ;
        RECT 28.225 -307.110 28.395 -306.165 ;
        RECT 28.690 -306.210 28.905 -305.780 ;
        RECT 26.175 -307.575 26.870 -307.345 ;
        RECT 22.985 -307.790 25.790 -307.620 ;
        RECT 22.985 -308.100 23.155 -307.790 ;
        RECT 19.775 -308.445 20.470 -308.175 ;
        RECT 22.425 -308.270 23.155 -308.100 ;
        RECT 22.425 -308.845 22.595 -308.270 ;
        RECT 23.520 -308.295 24.215 -308.025 ;
        RECT 18.660 -309.015 22.595 -308.845 ;
        RECT 22.900 -308.650 25.300 -308.480 ;
        RECT 15.725 -310.235 15.895 -309.280 ;
        RECT 7.280 -310.925 10.920 -310.755 ;
        RECT 19.780 -310.755 19.950 -309.195 ;
        RECT 20.270 -310.235 20.440 -309.015 ;
        RECT 20.760 -310.755 20.930 -309.195 ;
        RECT 21.360 -310.410 21.530 -309.195 ;
        RECT 21.850 -310.235 22.020 -309.015 ;
        RECT 22.340 -310.410 22.510 -309.195 ;
        RECT 22.900 -310.410 23.070 -308.650 ;
        RECT 21.360 -310.580 23.070 -310.410 ;
        RECT 23.250 -309.020 24.320 -308.850 ;
        RECT 23.250 -310.755 23.420 -309.020 ;
        RECT 24.150 -310.235 24.320 -309.020 ;
        RECT 25.130 -310.235 25.300 -308.650 ;
        RECT 25.565 -308.665 26.260 -308.395 ;
        RECT 26.655 -309.270 26.870 -307.575 ;
        RECT 28.205 -308.065 28.420 -307.110 ;
        RECT 28.715 -307.205 28.885 -306.210 ;
        RECT 34.760 -306.225 34.955 -305.610 ;
        RECT 35.270 -305.980 40.310 -305.800 ;
        RECT 40.685 -305.870 46.025 -305.610 ;
        RECT 48.355 -304.060 49.140 -303.860 ;
        RECT 33.160 -307.010 33.390 -306.330 ;
        RECT 27.705 -308.295 28.420 -308.065 ;
        RECT 26.680 -310.235 26.850 -309.270 ;
        RECT 28.205 -309.280 28.420 -308.295 ;
        RECT 28.640 -308.635 29.335 -308.365 ;
        RECT 33.190 -308.845 33.360 -307.010 ;
        RECT 34.780 -307.170 34.950 -306.225 ;
        RECT 34.770 -307.585 34.955 -307.170 ;
        RECT 35.270 -307.205 35.440 -305.980 ;
        RECT 36.850 -307.175 37.020 -306.165 ;
        RECT 37.340 -307.160 37.510 -306.165 ;
        RECT 38.660 -307.160 38.830 -306.165 ;
        RECT 36.835 -307.280 37.020 -307.175 ;
        RECT 36.240 -307.465 37.020 -307.280 ;
        RECT 37.330 -307.355 38.830 -307.160 ;
        RECT 36.240 -307.585 36.425 -307.465 ;
        RECT 34.770 -307.770 36.425 -307.585 ;
        RECT 39.150 -307.620 39.320 -306.165 ;
        RECT 40.130 -306.250 40.310 -305.980 ;
        RECT 40.130 -307.205 40.300 -306.250 ;
        RECT 40.620 -307.620 40.790 -306.165 ;
        RECT 41.680 -307.120 41.850 -306.165 ;
        RECT 42.145 -306.200 42.360 -305.870 ;
        RECT 41.655 -307.345 41.870 -307.120 ;
        RECT 42.170 -307.205 42.340 -306.200 ;
        RECT 43.225 -307.110 43.395 -306.165 ;
        RECT 43.690 -306.210 43.905 -305.870 ;
        RECT 41.175 -307.575 41.870 -307.345 ;
        RECT 37.985 -307.790 40.790 -307.620 ;
        RECT 37.985 -308.100 38.155 -307.790 ;
        RECT 34.775 -308.445 35.470 -308.175 ;
        RECT 37.425 -308.270 38.155 -308.100 ;
        RECT 37.425 -308.845 37.595 -308.270 ;
        RECT 38.520 -308.295 39.215 -308.025 ;
        RECT 33.190 -309.015 37.595 -308.845 ;
        RECT 37.900 -308.650 40.300 -308.480 ;
        RECT 28.225 -310.235 28.395 -309.280 ;
        RECT 19.780 -310.925 23.420 -310.755 ;
        RECT 34.780 -310.755 34.950 -309.195 ;
        RECT 35.270 -310.235 35.440 -309.015 ;
        RECT 35.760 -310.755 35.930 -309.195 ;
        RECT 36.360 -310.410 36.530 -309.195 ;
        RECT 36.850 -310.235 37.020 -309.015 ;
        RECT 37.340 -310.410 37.510 -309.195 ;
        RECT 37.900 -310.410 38.070 -308.650 ;
        RECT 36.360 -310.580 38.070 -310.410 ;
        RECT 38.250 -309.020 39.320 -308.850 ;
        RECT 38.250 -310.755 38.420 -309.020 ;
        RECT 39.150 -310.235 39.320 -309.020 ;
        RECT 40.130 -310.235 40.300 -308.650 ;
        RECT 40.565 -308.665 41.260 -308.395 ;
        RECT 41.655 -309.270 41.870 -307.575 ;
        RECT 43.205 -308.065 43.420 -307.110 ;
        RECT 43.715 -307.205 43.885 -306.210 ;
        RECT 42.705 -308.295 43.420 -308.065 ;
        RECT 41.680 -310.235 41.850 -309.270 ;
        RECT 43.205 -309.280 43.420 -308.295 ;
        RECT 43.640 -308.635 44.335 -308.365 ;
        RECT 43.225 -310.235 43.395 -309.280 ;
        RECT 34.780 -310.925 38.420 -310.755 ;
        RECT -33.040 -311.255 -32.225 -311.155 ;
        RECT -117.245 -311.555 -114.550 -311.360 ;
        RECT -140.735 -312.240 -114.550 -311.555 ;
        RECT -91.515 -311.935 -32.225 -311.255 ;
        RECT 48.355 -311.715 48.625 -304.060 ;
        RECT 49.425 -305.580 49.695 -303.425 ;
        RECT 48.930 -305.850 49.695 -305.580 ;
        RECT 48.930 -311.715 49.200 -305.850 ;
        RECT 49.650 -311.240 49.920 -311.090 ;
        RECT 50.140 -311.240 50.410 -302.750 ;
        RECT 52.735 -309.435 54.040 -300.535 ;
        RECT 67.815 -301.695 70.955 -301.525 ;
        RECT 60.355 -301.810 60.525 -301.790 ;
        RECT 60.325 -303.075 60.555 -301.810 ;
        RECT 61.335 -302.750 61.505 -301.790 ;
        RECT 62.315 -302.750 62.485 -301.790 ;
        RECT 64.765 -301.810 64.935 -301.790 ;
        RECT 63.660 -302.720 63.945 -301.900 ;
        RECT 61.305 -303.075 61.535 -302.750 ;
        RECT 62.285 -303.075 62.515 -302.750 ;
        RECT 60.325 -303.115 62.515 -303.075 ;
        RECT 64.735 -303.075 64.965 -301.810 ;
        RECT 65.745 -302.750 65.915 -301.790 ;
        RECT 66.725 -302.750 66.895 -301.790 ;
        RECT 67.815 -301.920 67.995 -301.695 ;
        RECT 65.715 -303.075 65.945 -302.750 ;
        RECT 66.695 -303.075 66.925 -302.750 ;
        RECT 64.735 -303.115 66.925 -303.075 ;
        RECT 67.200 -302.995 67.570 -302.155 ;
        RECT 67.820 -302.290 67.990 -301.920 ;
        RECT 67.200 -303.115 67.565 -302.995 ;
        RECT 60.325 -303.225 62.665 -303.115 ;
        RECT 63.715 -303.205 64.555 -303.150 ;
        RECT 62.955 -303.225 63.255 -303.205 ;
        RECT 63.540 -303.225 64.555 -303.205 ;
        RECT 60.325 -303.305 64.555 -303.225 ;
        RECT 59.865 -304.485 60.035 -303.690 ;
        RECT 60.325 -303.770 60.555 -303.305 ;
        RECT 60.355 -304.230 60.525 -303.770 ;
        RECT 60.845 -304.485 61.015 -303.690 ;
        RECT 61.305 -303.770 61.535 -303.305 ;
        RECT 62.285 -303.435 64.555 -303.305 ;
        RECT 62.285 -303.465 62.665 -303.435 ;
        RECT 61.335 -304.230 61.505 -303.770 ;
        RECT 61.825 -304.485 61.995 -303.690 ;
        RECT 62.285 -303.770 62.515 -303.465 ;
        RECT 62.315 -304.230 62.485 -303.770 ;
        RECT 62.955 -303.865 63.255 -303.435 ;
        RECT 63.540 -303.495 64.555 -303.435 ;
        RECT 63.715 -303.520 64.555 -303.495 ;
        RECT 64.735 -303.305 67.565 -303.115 ;
        RECT 64.275 -304.485 64.445 -303.690 ;
        RECT 64.735 -303.770 64.965 -303.305 ;
        RECT 64.765 -304.230 64.935 -303.770 ;
        RECT 65.255 -304.485 65.425 -303.690 ;
        RECT 65.715 -303.770 65.945 -303.305 ;
        RECT 66.695 -303.465 67.565 -303.305 ;
        RECT 67.790 -303.025 68.025 -302.290 ;
        RECT 68.310 -302.325 68.480 -301.865 ;
        RECT 68.795 -301.970 69.005 -301.695 ;
        RECT 68.305 -302.585 68.485 -302.325 ;
        RECT 68.800 -302.405 68.970 -301.970 ;
        RECT 69.290 -302.315 69.460 -301.865 ;
        RECT 69.765 -301.975 69.975 -301.695 ;
        RECT 69.290 -302.405 69.475 -302.315 ;
        RECT 69.780 -302.405 69.950 -301.975 ;
        RECT 70.270 -302.315 70.440 -301.865 ;
        RECT 70.745 -301.950 70.955 -301.695 ;
        RECT 81.315 -301.695 84.455 -301.525 ;
        RECT 73.480 -301.810 73.650 -301.790 ;
        RECT 69.295 -302.585 69.475 -302.405 ;
        RECT 70.265 -302.585 70.445 -302.315 ;
        RECT 70.760 -302.405 70.930 -301.950 ;
        RECT 71.250 -302.365 71.420 -301.865 ;
        RECT 71.235 -302.585 71.445 -302.365 ;
        RECT 68.305 -302.755 71.445 -302.585 ;
        RECT 67.790 -303.395 68.650 -303.025 ;
        RECT 70.570 -303.195 71.445 -302.755 ;
        RECT 73.450 -303.075 73.680 -301.810 ;
        RECT 74.460 -302.750 74.630 -301.790 ;
        RECT 75.440 -302.750 75.610 -301.790 ;
        RECT 78.265 -301.810 78.435 -301.790 ;
        RECT 77.160 -302.290 77.445 -301.900 ;
        RECT 76.140 -302.515 77.445 -302.290 ;
        RECT 74.430 -303.075 74.660 -302.750 ;
        RECT 75.410 -303.075 75.640 -302.750 ;
        RECT 73.450 -303.115 75.640 -303.075 ;
        RECT 72.430 -303.195 73.270 -303.150 ;
        RECT 65.745 -304.230 65.915 -303.770 ;
        RECT 66.235 -304.485 66.405 -303.690 ;
        RECT 66.695 -303.770 66.925 -303.465 ;
        RECT 66.725 -304.230 66.895 -303.770 ;
        RECT 67.790 -304.070 68.025 -303.395 ;
        RECT 70.570 -303.480 73.270 -303.195 ;
        RECT 70.570 -303.590 71.445 -303.480 ;
        RECT 72.430 -303.520 73.270 -303.480 ;
        RECT 73.450 -303.185 75.790 -303.115 ;
        RECT 76.140 -303.185 76.365 -302.515 ;
        RECT 77.160 -302.720 77.445 -302.515 ;
        RECT 73.450 -303.305 76.365 -303.185 ;
        RECT 68.290 -303.760 71.445 -303.590 ;
        RECT 68.290 -303.965 68.495 -303.760 ;
        RECT 67.820 -304.420 67.990 -304.070 ;
        RECT 59.820 -304.825 66.900 -304.485 ;
        RECT 67.795 -304.710 68.015 -304.420 ;
        RECT 68.310 -304.480 68.480 -303.965 ;
        RECT 68.800 -304.365 68.970 -303.940 ;
        RECT 69.280 -304.005 69.485 -303.760 ;
        RECT 68.775 -304.710 68.995 -304.365 ;
        RECT 69.290 -304.480 69.460 -304.005 ;
        RECT 69.780 -304.365 69.950 -303.940 ;
        RECT 70.250 -304.005 70.455 -303.760 ;
        RECT 71.235 -303.795 71.445 -303.760 ;
        RECT 69.755 -304.710 69.975 -304.365 ;
        RECT 70.270 -304.480 70.440 -304.005 ;
        RECT 70.760 -304.420 70.930 -303.940 ;
        RECT 71.235 -303.960 71.440 -303.795 ;
        RECT 71.205 -304.010 71.440 -303.960 ;
        RECT 70.740 -304.710 70.960 -304.420 ;
        RECT 71.205 -304.620 71.435 -304.010 ;
        RECT 72.990 -304.485 73.160 -303.690 ;
        RECT 73.450 -303.770 73.680 -303.305 ;
        RECT 73.480 -304.230 73.650 -303.770 ;
        RECT 73.970 -304.485 74.140 -303.690 ;
        RECT 74.430 -303.770 74.660 -303.305 ;
        RECT 75.410 -303.410 76.365 -303.305 ;
        RECT 78.235 -303.075 78.465 -301.810 ;
        RECT 79.245 -302.750 79.415 -301.790 ;
        RECT 80.225 -302.750 80.395 -301.790 ;
        RECT 81.315 -301.920 81.495 -301.695 ;
        RECT 79.215 -303.075 79.445 -302.750 ;
        RECT 80.195 -303.075 80.425 -302.750 ;
        RECT 78.235 -303.115 80.425 -303.075 ;
        RECT 80.700 -302.995 81.070 -302.155 ;
        RECT 81.320 -302.290 81.490 -301.920 ;
        RECT 80.700 -303.115 81.065 -302.995 ;
        RECT 78.235 -303.305 81.065 -303.115 ;
        RECT 75.410 -303.465 75.790 -303.410 ;
        RECT 74.460 -304.230 74.630 -303.770 ;
        RECT 74.950 -304.485 75.120 -303.690 ;
        RECT 75.410 -303.770 75.640 -303.465 ;
        RECT 75.440 -304.230 75.610 -303.770 ;
        RECT 76.040 -303.985 76.340 -303.410 ;
        RECT 77.775 -304.485 77.945 -303.690 ;
        RECT 78.235 -303.770 78.465 -303.305 ;
        RECT 78.265 -304.230 78.435 -303.770 ;
        RECT 78.755 -304.485 78.925 -303.690 ;
        RECT 79.215 -303.770 79.445 -303.305 ;
        RECT 80.195 -303.465 81.065 -303.305 ;
        RECT 81.290 -303.025 81.525 -302.290 ;
        RECT 81.810 -302.325 81.980 -301.865 ;
        RECT 82.295 -301.970 82.505 -301.695 ;
        RECT 81.805 -302.585 81.985 -302.325 ;
        RECT 82.300 -302.405 82.470 -301.970 ;
        RECT 82.790 -302.315 82.960 -301.865 ;
        RECT 83.265 -301.975 83.475 -301.695 ;
        RECT 82.790 -302.405 82.975 -302.315 ;
        RECT 83.280 -302.405 83.450 -301.975 ;
        RECT 83.770 -302.315 83.940 -301.865 ;
        RECT 84.245 -301.950 84.455 -301.695 ;
        RECT 86.980 -301.810 87.150 -301.790 ;
        RECT 82.795 -302.585 82.975 -302.405 ;
        RECT 83.765 -302.585 83.945 -302.315 ;
        RECT 84.260 -302.405 84.430 -301.950 ;
        RECT 84.750 -302.365 84.920 -301.865 ;
        RECT 84.735 -302.585 84.945 -302.365 ;
        RECT 81.805 -302.755 84.945 -302.585 ;
        RECT 81.290 -303.395 82.150 -303.025 ;
        RECT 84.070 -303.180 84.945 -302.755 ;
        RECT 86.950 -303.075 87.180 -301.810 ;
        RECT 87.960 -302.750 88.130 -301.790 ;
        RECT 88.940 -302.750 89.110 -301.790 ;
        RECT 87.930 -303.075 88.160 -302.750 ;
        RECT 88.910 -303.075 89.140 -302.750 ;
        RECT 86.950 -303.115 89.140 -303.075 ;
        RECT 85.930 -303.180 86.770 -303.150 ;
        RECT 79.245 -304.230 79.415 -303.770 ;
        RECT 79.735 -304.485 79.905 -303.690 ;
        RECT 80.195 -303.770 80.425 -303.465 ;
        RECT 80.225 -304.230 80.395 -303.770 ;
        RECT 81.290 -304.070 81.525 -303.395 ;
        RECT 84.070 -303.445 86.770 -303.180 ;
        RECT 84.070 -303.590 84.945 -303.445 ;
        RECT 85.930 -303.520 86.770 -303.445 ;
        RECT 86.950 -303.160 89.290 -303.115 ;
        RECT 86.950 -303.170 89.700 -303.160 ;
        RECT 86.950 -303.305 89.705 -303.170 ;
        RECT 81.790 -303.760 84.945 -303.590 ;
        RECT 81.790 -303.965 81.995 -303.760 ;
        RECT 81.320 -304.420 81.490 -304.070 ;
        RECT 67.795 -304.880 70.960 -304.710 ;
        RECT 72.945 -304.825 80.400 -304.485 ;
        RECT 81.295 -304.710 81.515 -304.420 ;
        RECT 81.810 -304.480 81.980 -303.965 ;
        RECT 82.300 -304.365 82.470 -303.940 ;
        RECT 82.780 -304.005 82.985 -303.760 ;
        RECT 82.275 -304.710 82.495 -304.365 ;
        RECT 82.790 -304.480 82.960 -304.005 ;
        RECT 83.280 -304.365 83.450 -303.940 ;
        RECT 83.750 -304.005 83.955 -303.760 ;
        RECT 84.735 -303.795 84.945 -303.760 ;
        RECT 83.255 -304.710 83.475 -304.365 ;
        RECT 83.770 -304.480 83.940 -304.005 ;
        RECT 84.260 -304.420 84.430 -303.940 ;
        RECT 84.735 -304.010 84.940 -303.795 ;
        RECT 84.240 -304.710 84.460 -304.420 ;
        RECT 84.750 -304.480 84.920 -304.010 ;
        RECT 86.490 -304.485 86.660 -303.690 ;
        RECT 86.950 -303.770 87.180 -303.305 ;
        RECT 86.980 -304.230 87.150 -303.770 ;
        RECT 87.470 -304.485 87.640 -303.690 ;
        RECT 87.930 -303.770 88.160 -303.305 ;
        RECT 88.910 -303.355 89.705 -303.305 ;
        RECT 88.910 -303.465 89.290 -303.355 ;
        RECT 87.960 -304.230 88.130 -303.770 ;
        RECT 88.450 -304.485 88.620 -303.690 ;
        RECT 88.910 -303.770 89.140 -303.465 ;
        RECT 88.940 -304.230 89.110 -303.770 ;
        RECT 81.295 -304.880 84.460 -304.710 ;
        RECT 86.445 -304.825 89.115 -304.485 ;
        RECT 62.750 -305.060 63.410 -305.005 ;
        RECT 85.365 -305.060 86.025 -304.995 ;
        RECT 62.750 -305.255 88.055 -305.060 ;
        RECT 89.465 -305.145 89.705 -303.355 ;
        RECT 62.750 -305.305 63.410 -305.255 ;
        RECT 85.365 -305.295 86.025 -305.255 ;
        RECT 89.410 -305.830 89.710 -305.145 ;
        RECT 61.135 -305.950 61.795 -305.855 ;
        RECT 74.300 -305.950 74.985 -305.855 ;
        RECT 87.285 -305.950 87.970 -305.885 ;
        RECT 61.130 -306.145 88.055 -305.950 ;
        RECT 61.135 -306.155 62.960 -306.145 ;
        RECT 61.655 -309.435 62.960 -306.155 ;
        RECT 64.740 -306.500 67.905 -306.330 ;
        RECT 69.925 -306.385 70.480 -306.145 ;
        RECT 74.300 -306.155 74.985 -306.145 ;
        RECT 71.355 -306.385 73.955 -306.375 ;
        RECT 74.315 -306.385 74.870 -306.155 ;
        RECT 64.280 -307.200 64.450 -306.730 ;
        RECT 64.740 -306.790 64.960 -306.500 ;
        RECT 64.260 -307.415 64.465 -307.200 ;
        RECT 64.770 -307.270 64.940 -306.790 ;
        RECT 65.260 -307.205 65.430 -306.730 ;
        RECT 65.725 -306.845 65.945 -306.500 ;
        RECT 64.255 -307.450 64.465 -307.415 ;
        RECT 65.245 -307.450 65.450 -307.205 ;
        RECT 65.750 -307.270 65.920 -306.845 ;
        RECT 66.240 -307.205 66.410 -306.730 ;
        RECT 66.705 -306.845 66.925 -306.500 ;
        RECT 66.215 -307.450 66.420 -307.205 ;
        RECT 66.730 -307.270 66.900 -306.845 ;
        RECT 67.220 -307.245 67.390 -306.730 ;
        RECT 67.685 -306.790 67.905 -306.500 ;
        RECT 68.800 -306.715 75.655 -306.385 ;
        RECT 68.800 -306.725 71.470 -306.715 ;
        RECT 72.985 -306.725 75.655 -306.715 ;
        RECT 78.240 -306.500 81.405 -306.330 ;
        RECT 83.305 -306.385 83.860 -306.145 ;
        RECT 87.285 -306.185 87.970 -306.145 ;
        RECT 87.360 -306.385 87.915 -306.185 ;
        RECT 67.710 -307.140 67.880 -306.790 ;
        RECT 67.205 -307.450 67.410 -307.245 ;
        RECT 64.255 -307.610 67.410 -307.450 ;
        RECT 63.880 -307.620 67.410 -307.610 ;
        RECT 63.880 -307.910 65.130 -307.620 ;
        RECT 67.675 -307.815 67.910 -307.140 ;
        RECT 68.805 -307.440 68.975 -306.980 ;
        RECT 68.775 -307.745 69.005 -307.440 ;
        RECT 69.295 -307.520 69.465 -306.725 ;
        RECT 69.785 -307.440 69.955 -306.980 ;
        RECT 64.255 -308.455 65.130 -307.910 ;
        RECT 67.050 -308.185 67.910 -307.815 ;
        RECT 64.255 -308.625 67.395 -308.455 ;
        RECT 64.255 -308.845 64.465 -308.625 ;
        RECT 64.280 -309.345 64.450 -308.845 ;
        RECT 64.770 -309.260 64.940 -308.805 ;
        RECT 65.255 -308.895 65.435 -308.625 ;
        RECT 66.225 -308.805 66.405 -308.625 ;
        RECT 52.735 -310.740 62.960 -309.435 ;
        RECT 64.745 -309.515 64.955 -309.260 ;
        RECT 65.260 -309.345 65.430 -308.895 ;
        RECT 65.750 -309.235 65.920 -308.805 ;
        RECT 66.225 -308.895 66.410 -308.805 ;
        RECT 65.725 -309.515 65.935 -309.235 ;
        RECT 66.240 -309.345 66.410 -308.895 ;
        RECT 66.730 -309.240 66.900 -308.805 ;
        RECT 67.215 -308.885 67.395 -308.625 ;
        RECT 66.695 -309.515 66.905 -309.240 ;
        RECT 67.220 -309.345 67.390 -308.885 ;
        RECT 67.675 -308.920 67.910 -308.185 ;
        RECT 68.135 -307.905 69.005 -307.745 ;
        RECT 69.755 -307.905 69.985 -307.440 ;
        RECT 70.275 -307.520 70.445 -306.725 ;
        RECT 70.765 -307.440 70.935 -306.980 ;
        RECT 70.735 -307.905 70.965 -307.440 ;
        RECT 71.255 -307.520 71.425 -306.725 ;
        RECT 72.990 -307.440 73.160 -306.980 ;
        RECT 72.960 -307.745 73.190 -307.440 ;
        RECT 73.480 -307.520 73.650 -306.725 ;
        RECT 73.970 -307.440 74.140 -306.980 ;
        RECT 68.135 -308.095 70.965 -307.905 ;
        RECT 68.135 -308.215 68.500 -308.095 ;
        RECT 67.710 -309.290 67.880 -308.920 ;
        RECT 68.130 -309.055 68.500 -308.215 ;
        RECT 68.775 -308.135 70.965 -308.095 ;
        RECT 68.775 -308.460 69.005 -308.135 ;
        RECT 69.755 -308.460 69.985 -308.135 ;
        RECT 67.705 -309.515 67.885 -309.290 ;
        RECT 68.805 -309.420 68.975 -308.460 ;
        RECT 69.785 -309.420 69.955 -308.460 ;
        RECT 70.735 -309.400 70.965 -308.135 ;
        RECT 72.470 -307.905 73.190 -307.745 ;
        RECT 73.940 -307.905 74.170 -307.440 ;
        RECT 74.460 -307.520 74.630 -306.725 ;
        RECT 74.950 -307.440 75.120 -306.980 ;
        RECT 74.920 -307.905 75.150 -307.440 ;
        RECT 75.440 -307.520 75.610 -306.725 ;
        RECT 77.780 -307.200 77.950 -306.730 ;
        RECT 78.240 -306.790 78.460 -306.500 ;
        RECT 77.760 -307.415 77.965 -307.200 ;
        RECT 78.270 -307.270 78.440 -306.790 ;
        RECT 78.760 -307.205 78.930 -306.730 ;
        RECT 79.225 -306.845 79.445 -306.500 ;
        RECT 77.755 -307.450 77.965 -307.415 ;
        RECT 78.745 -307.450 78.950 -307.205 ;
        RECT 79.250 -307.270 79.420 -306.845 ;
        RECT 79.740 -307.205 79.910 -306.730 ;
        RECT 80.205 -306.845 80.425 -306.500 ;
        RECT 79.715 -307.450 79.920 -307.205 ;
        RECT 80.230 -307.270 80.400 -306.845 ;
        RECT 80.720 -307.245 80.890 -306.730 ;
        RECT 81.185 -306.790 81.405 -306.500 ;
        RECT 82.300 -306.725 89.155 -306.385 ;
        RECT 81.210 -307.140 81.380 -306.790 ;
        RECT 80.705 -307.450 80.910 -307.245 ;
        RECT 77.755 -307.620 80.910 -307.450 ;
        RECT 72.470 -308.095 75.150 -307.905 ;
        RECT 75.330 -307.725 76.170 -307.690 ;
        RECT 75.330 -308.025 76.280 -307.725 ;
        RECT 77.300 -307.920 78.630 -307.620 ;
        RECT 81.175 -307.815 81.410 -307.140 ;
        RECT 82.305 -307.440 82.475 -306.980 ;
        RECT 82.275 -307.745 82.505 -307.440 ;
        RECT 82.795 -307.520 82.965 -306.725 ;
        RECT 83.285 -307.440 83.455 -306.980 ;
        RECT 75.330 -308.060 76.170 -308.025 ;
        RECT 71.755 -308.740 72.040 -308.490 ;
        RECT 72.470 -308.740 72.780 -308.095 ;
        RECT 72.960 -308.135 75.150 -308.095 ;
        RECT 72.960 -308.460 73.190 -308.135 ;
        RECT 73.940 -308.460 74.170 -308.135 ;
        RECT 71.755 -309.050 72.780 -308.740 ;
        RECT 71.755 -309.310 72.040 -309.050 ;
        RECT 70.765 -309.420 70.935 -309.400 ;
        RECT 72.990 -309.420 73.160 -308.460 ;
        RECT 73.970 -309.420 74.140 -308.460 ;
        RECT 74.920 -309.400 75.150 -308.135 ;
        RECT 77.755 -308.455 78.630 -307.920 ;
        RECT 80.550 -308.185 81.410 -307.815 ;
        RECT 77.755 -308.625 80.895 -308.455 ;
        RECT 77.755 -308.845 77.965 -308.625 ;
        RECT 77.780 -309.345 77.950 -308.845 ;
        RECT 78.270 -309.260 78.440 -308.805 ;
        RECT 78.755 -308.895 78.935 -308.625 ;
        RECT 79.725 -308.805 79.905 -308.625 ;
        RECT 74.950 -309.420 75.120 -309.400 ;
        RECT 64.745 -309.685 67.885 -309.515 ;
        RECT 78.245 -309.515 78.455 -309.260 ;
        RECT 78.760 -309.345 78.930 -308.895 ;
        RECT 79.250 -309.235 79.420 -308.805 ;
        RECT 79.725 -308.895 79.910 -308.805 ;
        RECT 79.225 -309.515 79.435 -309.235 ;
        RECT 79.740 -309.345 79.910 -308.895 ;
        RECT 80.230 -309.240 80.400 -308.805 ;
        RECT 80.715 -308.885 80.895 -308.625 ;
        RECT 80.195 -309.515 80.405 -309.240 ;
        RECT 80.720 -309.345 80.890 -308.885 ;
        RECT 81.175 -308.920 81.410 -308.185 ;
        RECT 81.635 -307.905 82.505 -307.745 ;
        RECT 83.255 -307.905 83.485 -307.440 ;
        RECT 83.775 -307.520 83.945 -306.725 ;
        RECT 84.265 -307.440 84.435 -306.980 ;
        RECT 84.235 -307.905 84.465 -307.440 ;
        RECT 84.755 -307.520 84.925 -306.725 ;
        RECT 85.545 -307.690 85.845 -306.970 ;
        RECT 86.490 -307.440 86.660 -306.980 ;
        RECT 81.635 -308.095 84.465 -307.905 ;
        RECT 84.645 -308.000 85.845 -307.690 ;
        RECT 86.460 -307.745 86.690 -307.440 ;
        RECT 86.980 -307.520 87.150 -306.725 ;
        RECT 87.470 -307.440 87.640 -306.980 ;
        RECT 86.025 -307.905 86.690 -307.745 ;
        RECT 87.440 -307.905 87.670 -307.440 ;
        RECT 87.960 -307.520 88.130 -306.725 ;
        RECT 88.450 -307.440 88.620 -306.980 ;
        RECT 88.420 -307.905 88.650 -307.440 ;
        RECT 88.940 -307.520 89.110 -306.725 ;
        RECT 89.465 -307.690 89.705 -305.830 ;
        RECT 84.645 -308.005 85.660 -308.000 ;
        RECT 84.645 -308.060 85.485 -308.005 ;
        RECT 81.635 -308.215 82.000 -308.095 ;
        RECT 81.210 -309.290 81.380 -308.920 ;
        RECT 81.630 -309.055 82.000 -308.215 ;
        RECT 82.275 -308.135 84.465 -308.095 ;
        RECT 82.275 -308.460 82.505 -308.135 ;
        RECT 83.255 -308.460 83.485 -308.135 ;
        RECT 81.205 -309.515 81.385 -309.290 ;
        RECT 82.305 -309.420 82.475 -308.460 ;
        RECT 83.285 -309.420 83.455 -308.460 ;
        RECT 84.235 -309.400 84.465 -308.135 ;
        RECT 86.025 -308.095 88.650 -307.905 ;
        RECT 88.830 -307.910 89.705 -307.690 ;
        RECT 88.830 -308.060 89.670 -307.910 ;
        RECT 85.255 -308.745 85.540 -308.490 ;
        RECT 86.025 -308.745 86.255 -308.095 ;
        RECT 86.460 -308.135 88.650 -308.095 ;
        RECT 86.460 -308.460 86.690 -308.135 ;
        RECT 87.440 -308.460 87.670 -308.135 ;
        RECT 85.255 -308.990 86.255 -308.745 ;
        RECT 85.255 -309.310 85.540 -308.990 ;
        RECT 84.265 -309.420 84.435 -309.400 ;
        RECT 86.490 -309.420 86.660 -308.460 ;
        RECT 87.470 -309.420 87.640 -308.460 ;
        RECT 88.420 -309.400 88.650 -308.135 ;
        RECT 136.450 -309.195 137.180 -290.445 ;
        RECT 140.430 -291.285 140.810 -290.445 ;
        RECT 140.430 -291.665 141.140 -291.285 ;
        RECT 140.760 -293.610 141.140 -291.665 ;
        RECT 145.805 -291.495 149.130 -291.355 ;
        RECT 145.805 -291.785 150.980 -291.495 ;
        RECT 154.850 -291.780 155.310 -291.355 ;
        RECT 145.805 -292.190 146.235 -291.785 ;
        RECT 147.105 -291.970 147.280 -291.785 ;
        RECT 148.730 -291.800 150.980 -291.785 ;
        RECT 141.545 -292.620 146.235 -292.190 ;
        RECT 140.760 -294.070 141.435 -293.610 ;
        RECT 142.245 -293.900 142.415 -292.620 ;
        RECT 142.735 -293.900 142.905 -292.860 ;
        RECT 143.225 -293.900 143.395 -292.620 ;
        RECT 143.715 -293.730 143.885 -292.860 ;
        RECT 146.620 -293.510 146.790 -291.970 ;
        RECT 147.110 -293.510 147.280 -291.970 ;
        RECT 147.600 -293.510 147.770 -291.970 ;
        RECT 148.090 -293.510 148.260 -291.970 ;
        RECT 148.580 -293.510 148.750 -291.970 ;
        RECT 146.460 -293.725 146.815 -293.720 ;
        RECT 148.520 -293.725 148.890 -293.695 ;
        RECT 146.460 -293.730 148.890 -293.725 ;
        RECT 143.715 -293.900 148.890 -293.730 ;
        RECT 150.675 -293.835 150.980 -291.800 ;
        RECT 143.720 -293.920 148.890 -293.900 ;
        RECT 143.720 -293.930 146.465 -293.920 ;
        RECT 141.655 -294.070 142.020 -294.040 ;
        RECT 148.520 -294.050 148.890 -293.920 ;
        RECT 140.760 -294.155 142.020 -294.070 ;
        RECT 140.785 -294.275 142.020 -294.155 ;
        RECT 146.195 -294.210 146.870 -294.170 ;
        RECT 146.095 -294.220 146.870 -294.210 ;
        RECT 140.785 -294.360 141.435 -294.275 ;
        RECT 141.655 -294.340 142.020 -294.275 ;
        RECT 145.060 -294.400 146.870 -294.220 ;
        RECT 149.455 -294.265 153.380 -293.835 ;
        RECT 146.095 -294.410 146.870 -294.400 ;
        RECT 146.195 -294.440 146.870 -294.410 ;
        RECT 147.110 -294.325 149.205 -294.285 ;
        RECT 147.110 -294.475 149.260 -294.325 ;
        RECT 142.245 -295.550 142.415 -294.510 ;
        RECT 143.225 -295.550 143.395 -294.510 ;
        RECT 144.205 -295.550 144.375 -294.510 ;
        RECT 147.110 -296.195 147.280 -294.475 ;
        RECT 148.090 -296.195 148.260 -294.475 ;
        RECT 148.955 -295.220 149.260 -294.475 ;
        RECT 150.155 -295.045 150.325 -294.265 ;
        RECT 150.645 -295.045 150.815 -294.505 ;
        RECT 151.135 -295.045 151.305 -294.265 ;
        RECT 151.625 -295.045 151.795 -294.505 ;
        RECT 149.565 -295.220 149.930 -295.190 ;
        RECT 148.955 -295.285 149.930 -295.220 ;
        RECT 149.065 -295.425 149.930 -295.285 ;
        RECT 149.565 -295.490 149.930 -295.425 ;
        RECT 152.115 -295.340 153.975 -294.990 ;
        RECT 150.155 -296.200 150.325 -295.660 ;
        RECT 151.135 -296.200 151.305 -295.660 ;
        RECT 152.115 -296.200 152.285 -295.340 ;
        RECT 150.385 -298.540 151.585 -298.370 ;
        RECT 142.115 -300.875 142.285 -299.155 ;
        RECT 143.095 -300.875 143.265 -299.155 ;
        RECT 145.160 -299.690 145.330 -299.150 ;
        RECT 146.140 -299.690 146.310 -299.150 ;
        RECT 144.570 -299.925 144.935 -299.860 ;
        RECT 144.070 -300.065 144.935 -299.925 ;
        RECT 143.960 -300.130 144.935 -300.065 ;
        RECT 143.960 -300.875 144.265 -300.130 ;
        RECT 144.570 -300.160 144.935 -300.130 ;
        RECT 147.120 -300.010 147.290 -299.150 ;
        RECT 142.115 -301.025 144.265 -300.875 ;
        RECT 142.115 -301.065 144.210 -301.025 ;
        RECT 145.160 -301.085 145.330 -300.305 ;
        RECT 145.650 -300.845 145.820 -300.305 ;
        RECT 146.140 -301.085 146.310 -300.305 ;
        RECT 146.630 -300.845 146.800 -300.305 ;
        RECT 147.120 -300.360 148.510 -300.010 ;
        RECT 140.335 -301.430 141.470 -301.420 ;
        RECT 143.525 -301.430 143.895 -301.300 ;
        RECT 140.335 -301.620 143.895 -301.430 ;
        RECT 144.460 -301.515 147.535 -301.085 ;
        RECT 141.465 -301.625 143.895 -301.620 ;
        RECT 141.465 -301.630 141.820 -301.625 ;
        RECT 143.525 -301.655 143.895 -301.625 ;
        RECT 141.625 -303.380 141.795 -301.840 ;
        RECT 142.115 -303.380 142.285 -301.840 ;
        RECT 142.605 -303.380 142.775 -301.840 ;
        RECT 143.095 -303.380 143.265 -301.840 ;
        RECT 143.585 -303.380 143.755 -301.840 ;
        RECT 142.110 -303.640 142.285 -303.380 ;
        RECT 145.680 -303.550 145.985 -301.515 ;
        RECT 148.130 -302.335 148.480 -300.360 ;
        RECT 149.350 -301.630 149.520 -298.710 ;
        RECT 150.385 -298.750 150.595 -298.540 ;
        RECT 149.330 -301.925 149.540 -301.630 ;
        RECT 150.405 -301.660 150.575 -298.750 ;
        RECT 150.895 -301.650 151.065 -298.710 ;
        RECT 151.375 -298.760 151.585 -298.540 ;
        RECT 150.390 -301.925 150.600 -301.660 ;
        RECT 149.330 -302.105 150.600 -301.925 ;
        RECT 150.875 -301.920 151.085 -301.650 ;
        RECT 151.385 -301.750 151.555 -298.760 ;
        RECT 152.445 -301.680 152.615 -298.710 ;
        RECT 150.875 -302.115 151.580 -301.920 ;
        RECT 151.365 -302.175 151.580 -302.115 ;
        RECT 150.155 -302.335 150.930 -302.285 ;
        RECT 148.130 -302.515 150.930 -302.335 ;
        RECT 148.130 -302.525 148.480 -302.515 ;
        RECT 150.155 -302.560 150.930 -302.515 ;
        RECT 151.365 -302.450 152.270 -302.175 ;
        RECT 151.365 -302.800 151.580 -302.450 ;
        RECT 148.805 -302.870 149.580 -302.825 ;
        RECT 148.620 -303.040 149.580 -302.870 ;
        RECT 148.805 -303.100 149.580 -303.040 ;
        RECT 149.810 -303.000 151.580 -302.800 ;
        RECT 152.440 -302.900 152.655 -301.680 ;
        RECT 153.625 -302.025 153.975 -295.340 ;
        RECT 154.965 -301.655 155.180 -291.780 ;
        RECT 156.600 -293.895 156.980 -290.375 ;
        RECT 158.110 -290.155 167.045 -289.965 ;
        RECT 179.350 -289.390 183.010 -288.660 ;
        RECT 187.920 -288.120 188.225 -286.645 ;
        RECT 191.590 -287.530 191.760 -286.060 ;
        RECT 192.050 -286.140 192.275 -285.790 ;
        RECT 194.010 -285.890 198.630 -285.690 ;
        RECT 194.250 -285.905 198.630 -285.890 ;
        RECT 191.555 -288.120 191.790 -287.530 ;
        RECT 192.080 -287.600 192.250 -286.140 ;
        RECT 192.570 -287.525 192.740 -286.060 ;
        RECT 193.780 -287.475 193.950 -286.060 ;
        RECT 194.250 -286.105 194.470 -285.905 ;
        RECT 199.620 -286.015 200.015 -285.665 ;
        RECT 192.535 -288.120 192.770 -287.525 ;
        RECT 193.745 -288.120 193.980 -287.475 ;
        RECT 194.270 -287.600 194.440 -286.105 ;
        RECT 201.060 -287.225 201.230 -285.770 ;
        RECT 201.050 -287.780 201.235 -287.225 ;
        RECT 201.550 -287.310 201.720 -284.085 ;
        RECT 202.695 -284.435 202.885 -284.085 ;
        RECT 203.895 -284.275 204.065 -283.880 ;
        RECT 205.270 -283.925 205.960 -283.880 ;
        RECT 202.645 -285.125 202.915 -284.435 ;
        RECT 203.410 -284.445 204.065 -284.275 ;
        RECT 204.395 -284.360 205.085 -284.090 ;
        RECT 206.320 -284.435 206.590 -283.745 ;
        RECT 206.780 -283.750 206.950 -283.530 ;
        RECT 206.780 -284.020 207.610 -283.750 ;
        RECT 203.410 -287.310 203.580 -284.445 ;
        RECT 206.780 -284.595 206.950 -284.020 ;
        RECT 207.210 -284.595 207.480 -284.510 ;
        RECT 203.900 -284.790 204.695 -284.615 ;
        RECT 206.780 -284.620 207.480 -284.595 ;
        RECT 206.640 -284.765 207.480 -284.620 ;
        RECT 203.900 -287.310 204.070 -284.790 ;
        RECT 204.525 -287.310 204.695 -284.790 ;
        RECT 205.015 -287.225 205.185 -284.770 ;
        RECT 205.665 -287.220 205.835 -284.770 ;
        RECT 198.365 -287.800 201.420 -287.780 ;
        RECT 205.010 -287.800 205.195 -287.225 ;
        RECT 205.650 -287.800 205.835 -287.220 ;
        RECT 206.155 -287.310 206.325 -284.770 ;
        RECT 206.640 -284.790 206.950 -284.765 ;
        RECT 206.645 -287.310 206.815 -284.790 ;
        RECT 207.210 -284.805 207.480 -284.765 ;
        RECT 207.785 -285.355 207.975 -282.890 ;
        RECT 228.670 -283.860 228.840 -282.140 ;
        RECT 229.650 -283.860 229.820 -282.140 ;
        RECT 231.715 -282.675 231.885 -282.135 ;
        RECT 232.695 -282.675 232.865 -282.135 ;
        RECT 231.125 -282.910 231.490 -282.845 ;
        RECT 230.625 -283.050 231.490 -282.910 ;
        RECT 230.515 -283.115 231.490 -283.050 ;
        RECT 230.515 -283.860 230.820 -283.115 ;
        RECT 231.125 -283.145 231.490 -283.115 ;
        RECT 233.675 -282.995 233.845 -282.135 ;
        RECT 228.670 -284.010 230.820 -283.860 ;
        RECT 228.670 -284.050 230.765 -284.010 ;
        RECT 231.715 -284.070 231.885 -283.290 ;
        RECT 232.205 -283.830 232.375 -283.290 ;
        RECT 232.695 -284.070 232.865 -283.290 ;
        RECT 233.185 -283.830 233.355 -283.290 ;
        RECT 233.675 -283.345 235.065 -282.995 ;
        RECT 226.890 -284.415 228.025 -284.405 ;
        RECT 230.080 -284.415 230.450 -284.285 ;
        RECT 226.890 -284.605 230.450 -284.415 ;
        RECT 231.015 -284.500 234.090 -284.070 ;
        RECT 207.785 -285.545 209.245 -285.355 ;
        RECT 207.295 -287.215 207.465 -285.770 ;
        RECT 207.785 -285.795 207.975 -285.545 ;
        RECT 207.285 -287.800 207.470 -287.215 ;
        RECT 207.785 -287.310 207.955 -285.795 ;
        RECT 198.365 -288.120 208.035 -287.800 ;
        RECT 187.920 -288.345 208.035 -288.120 ;
        RECT 187.920 -288.685 198.930 -288.345 ;
        RECT 200.670 -288.605 208.035 -288.345 ;
        RECT 158.110 -292.045 158.300 -290.155 ;
        RECT 164.145 -291.650 167.470 -291.510 ;
        RECT 164.145 -291.940 169.320 -291.650 ;
        RECT 157.995 -292.315 158.360 -292.045 ;
        RECT 164.145 -292.345 164.575 -291.940 ;
        RECT 165.445 -292.125 165.620 -291.940 ;
        RECT 167.070 -291.955 169.320 -291.940 ;
        RECT 159.885 -292.775 164.575 -292.345 ;
        RECT 159.125 -293.895 159.775 -293.765 ;
        RECT 156.600 -294.225 159.775 -293.895 ;
        RECT 160.585 -294.055 160.755 -292.775 ;
        RECT 161.075 -294.055 161.245 -293.015 ;
        RECT 161.565 -294.055 161.735 -292.775 ;
        RECT 162.055 -293.885 162.225 -293.015 ;
        RECT 164.960 -293.665 165.130 -292.125 ;
        RECT 165.450 -293.665 165.620 -292.125 ;
        RECT 165.940 -293.665 166.110 -292.125 ;
        RECT 166.430 -293.665 166.600 -292.125 ;
        RECT 166.920 -293.665 167.090 -292.125 ;
        RECT 164.800 -293.880 165.155 -293.875 ;
        RECT 166.860 -293.880 167.230 -293.850 ;
        RECT 164.800 -293.885 167.230 -293.880 ;
        RECT 162.055 -294.055 167.230 -293.885 ;
        RECT 169.015 -293.990 169.320 -291.955 ;
        RECT 162.060 -294.075 167.230 -294.055 ;
        RECT 162.060 -294.085 164.805 -294.075 ;
        RECT 159.995 -294.225 160.360 -294.195 ;
        RECT 166.860 -294.205 167.230 -294.075 ;
        RECT 156.600 -294.275 160.360 -294.225 ;
        RECT 159.125 -294.430 160.360 -294.275 ;
        RECT 164.535 -294.365 165.210 -294.325 ;
        RECT 164.435 -294.375 165.210 -294.365 ;
        RECT 159.125 -294.515 159.775 -294.430 ;
        RECT 159.995 -294.495 160.360 -294.430 ;
        RECT 159.260 -294.765 159.640 -294.515 ;
        RECT 163.400 -294.555 165.210 -294.375 ;
        RECT 167.795 -294.420 171.720 -293.990 ;
        RECT 164.435 -294.565 165.210 -294.555 ;
        RECT 164.535 -294.595 165.210 -294.565 ;
        RECT 165.450 -294.480 167.545 -294.440 ;
        RECT 165.450 -294.630 167.600 -294.480 ;
        RECT 160.585 -295.705 160.755 -294.665 ;
        RECT 161.565 -295.705 161.735 -294.665 ;
        RECT 162.545 -295.705 162.715 -294.665 ;
        RECT 165.450 -296.350 165.620 -294.630 ;
        RECT 166.430 -296.350 166.600 -294.630 ;
        RECT 167.295 -295.375 167.600 -294.630 ;
        RECT 168.495 -295.200 168.665 -294.420 ;
        RECT 168.985 -295.200 169.155 -294.660 ;
        RECT 169.475 -295.200 169.645 -294.420 ;
        RECT 169.965 -295.200 170.135 -294.660 ;
        RECT 167.905 -295.375 168.270 -295.345 ;
        RECT 167.295 -295.440 168.270 -295.375 ;
        RECT 167.405 -295.580 168.270 -295.440 ;
        RECT 167.905 -295.645 168.270 -295.580 ;
        RECT 170.455 -295.495 172.315 -295.145 ;
        RECT 168.495 -296.355 168.665 -295.815 ;
        RECT 169.475 -296.355 169.645 -295.815 ;
        RECT 170.455 -296.355 170.625 -295.495 ;
        RECT 168.725 -298.695 169.925 -298.525 ;
        RECT 160.455 -301.030 160.625 -299.310 ;
        RECT 161.435 -301.030 161.605 -299.310 ;
        RECT 163.500 -299.845 163.670 -299.305 ;
        RECT 164.480 -299.845 164.650 -299.305 ;
        RECT 162.910 -300.080 163.275 -300.015 ;
        RECT 162.410 -300.220 163.275 -300.080 ;
        RECT 162.300 -300.285 163.275 -300.220 ;
        RECT 162.300 -301.030 162.605 -300.285 ;
        RECT 162.910 -300.315 163.275 -300.285 ;
        RECT 165.460 -300.165 165.630 -299.305 ;
        RECT 160.455 -301.180 162.605 -301.030 ;
        RECT 160.455 -301.220 162.550 -301.180 ;
        RECT 163.500 -301.240 163.670 -300.460 ;
        RECT 163.990 -301.000 164.160 -300.460 ;
        RECT 164.480 -301.240 164.650 -300.460 ;
        RECT 164.970 -301.000 165.140 -300.460 ;
        RECT 165.460 -300.515 166.850 -300.165 ;
        RECT 158.675 -301.585 159.810 -301.575 ;
        RECT 161.865 -301.585 162.235 -301.455 ;
        RECT 154.965 -301.870 156.390 -301.655 ;
        RECT 158.675 -301.775 162.235 -301.585 ;
        RECT 162.800 -301.670 165.875 -301.240 ;
        RECT 159.805 -301.780 162.235 -301.775 ;
        RECT 159.805 -301.785 160.160 -301.780 ;
        RECT 161.865 -301.810 162.235 -301.780 ;
        RECT 153.570 -302.385 154.095 -302.025 ;
        RECT 156.175 -302.900 156.390 -301.870 ;
        RECT 143.735 -303.640 145.985 -303.550 ;
        RECT 141.525 -303.855 145.985 -303.640 ;
        RECT 141.525 -303.945 143.770 -303.855 ;
        RECT 145.680 -305.330 145.985 -303.855 ;
        RECT 149.350 -304.740 149.520 -303.270 ;
        RECT 149.810 -303.350 150.035 -303.000 ;
        RECT 151.770 -303.100 156.390 -302.900 ;
        RECT 152.010 -303.115 156.390 -303.100 ;
        RECT 149.315 -305.330 149.550 -304.740 ;
        RECT 149.840 -304.810 150.010 -303.350 ;
        RECT 150.330 -304.735 150.500 -303.270 ;
        RECT 151.540 -304.685 151.710 -303.270 ;
        RECT 152.010 -303.315 152.230 -303.115 ;
        RECT 150.295 -305.330 150.530 -304.735 ;
        RECT 151.505 -305.330 151.740 -304.685 ;
        RECT 152.030 -304.810 152.200 -303.315 ;
        RECT 159.965 -303.535 160.135 -301.995 ;
        RECT 160.455 -303.535 160.625 -301.995 ;
        RECT 160.945 -303.535 161.115 -301.995 ;
        RECT 161.435 -303.535 161.605 -301.995 ;
        RECT 161.925 -303.535 162.095 -301.995 ;
        RECT 160.450 -303.795 160.625 -303.535 ;
        RECT 164.020 -303.705 164.325 -301.670 ;
        RECT 166.470 -302.490 166.820 -300.515 ;
        RECT 167.690 -301.785 167.860 -298.865 ;
        RECT 168.725 -298.905 168.935 -298.695 ;
        RECT 167.670 -302.080 167.880 -301.785 ;
        RECT 168.745 -301.815 168.915 -298.905 ;
        RECT 169.235 -301.805 169.405 -298.865 ;
        RECT 169.715 -298.915 169.925 -298.695 ;
        RECT 168.730 -302.080 168.940 -301.815 ;
        RECT 167.670 -302.260 168.940 -302.080 ;
        RECT 169.215 -302.075 169.425 -301.805 ;
        RECT 169.725 -301.905 169.895 -298.915 ;
        RECT 170.785 -301.835 170.955 -298.865 ;
        RECT 169.215 -302.270 169.920 -302.075 ;
        RECT 169.705 -302.330 169.920 -302.270 ;
        RECT 168.495 -302.490 169.270 -302.440 ;
        RECT 166.470 -302.670 169.270 -302.490 ;
        RECT 166.470 -302.680 166.820 -302.670 ;
        RECT 168.495 -302.715 169.270 -302.670 ;
        RECT 169.705 -302.605 170.610 -302.330 ;
        RECT 169.705 -302.955 169.920 -302.605 ;
        RECT 167.145 -303.025 167.920 -302.980 ;
        RECT 166.960 -303.195 167.920 -303.025 ;
        RECT 167.145 -303.255 167.920 -303.195 ;
        RECT 168.150 -303.155 169.920 -302.955 ;
        RECT 170.780 -303.055 170.995 -301.835 ;
        RECT 171.965 -302.180 172.315 -295.495 ;
        RECT 171.910 -302.540 172.435 -302.180 ;
        RECT 174.440 -303.055 175.555 -302.605 ;
        RECT 162.075 -303.795 164.325 -303.705 ;
        RECT 159.865 -304.010 164.325 -303.795 ;
        RECT 159.865 -304.100 162.110 -304.010 ;
        RECT 145.680 -305.895 153.065 -305.330 ;
        RECT 164.020 -305.485 164.325 -304.010 ;
        RECT 167.690 -304.895 167.860 -303.425 ;
        RECT 168.150 -303.505 168.375 -303.155 ;
        RECT 170.110 -303.255 176.120 -303.055 ;
        RECT 170.350 -303.270 176.120 -303.255 ;
        RECT 167.655 -305.485 167.890 -304.895 ;
        RECT 168.180 -304.965 168.350 -303.505 ;
        RECT 168.670 -304.890 168.840 -303.425 ;
        RECT 169.880 -304.840 170.050 -303.425 ;
        RECT 170.350 -303.470 170.570 -303.270 ;
        RECT 174.440 -303.455 175.555 -303.270 ;
        RECT 168.635 -305.485 168.870 -304.890 ;
        RECT 169.845 -305.485 170.080 -304.840 ;
        RECT 170.370 -304.965 170.540 -303.470 ;
        RECT 164.020 -306.050 171.405 -305.485 ;
        RECT 127.120 -309.205 137.180 -309.195 ;
        RECT 88.450 -309.420 88.620 -309.400 ;
        RECT 78.245 -309.685 81.385 -309.515 ;
        RECT 127.120 -310.045 137.275 -309.205 ;
        RECT 179.350 -309.305 180.080 -289.390 ;
        RECT 182.630 -290.050 183.010 -289.390 ;
        RECT 209.055 -290.020 209.245 -285.545 ;
        RECT 226.945 -289.295 227.325 -284.605 ;
        RECT 228.020 -284.610 230.450 -284.605 ;
        RECT 228.020 -284.615 228.375 -284.610 ;
        RECT 230.080 -284.640 230.450 -284.610 ;
        RECT 228.180 -286.365 228.350 -284.825 ;
        RECT 228.670 -286.365 228.840 -284.825 ;
        RECT 229.160 -286.365 229.330 -284.825 ;
        RECT 229.650 -286.365 229.820 -284.825 ;
        RECT 230.140 -286.365 230.310 -284.825 ;
        RECT 228.665 -286.625 228.840 -286.365 ;
        RECT 232.235 -286.535 232.540 -284.500 ;
        RECT 234.685 -285.320 235.035 -283.345 ;
        RECT 235.905 -284.615 236.075 -281.695 ;
        RECT 236.940 -281.735 237.150 -281.525 ;
        RECT 235.885 -284.910 236.095 -284.615 ;
        RECT 236.960 -284.645 237.130 -281.735 ;
        RECT 237.450 -284.635 237.620 -281.695 ;
        RECT 237.930 -281.745 238.140 -281.525 ;
        RECT 236.945 -284.910 237.155 -284.645 ;
        RECT 235.885 -285.090 237.155 -284.910 ;
        RECT 237.430 -284.905 237.640 -284.635 ;
        RECT 237.940 -284.735 238.110 -281.745 ;
        RECT 239.000 -284.665 239.170 -281.695 ;
        RECT 237.430 -285.100 238.135 -284.905 ;
        RECT 237.920 -285.160 238.135 -285.100 ;
        RECT 236.710 -285.320 237.485 -285.270 ;
        RECT 234.685 -285.500 237.485 -285.320 ;
        RECT 234.685 -285.510 235.035 -285.500 ;
        RECT 236.710 -285.545 237.485 -285.500 ;
        RECT 237.920 -285.435 238.825 -285.160 ;
        RECT 237.920 -285.785 238.135 -285.435 ;
        RECT 235.360 -285.855 236.135 -285.810 ;
        RECT 235.175 -286.025 236.135 -285.855 ;
        RECT 235.360 -286.085 236.135 -286.025 ;
        RECT 236.365 -285.985 238.135 -285.785 ;
        RECT 238.995 -285.885 239.210 -284.665 ;
        RECT 240.180 -285.010 240.530 -278.325 ;
        RECT 274.790 -278.365 274.960 -277.325 ;
        RECT 275.770 -278.365 275.940 -277.325 ;
        RECT 276.750 -278.365 276.920 -277.325 ;
        RECT 279.655 -279.010 279.825 -277.290 ;
        RECT 280.635 -279.010 280.805 -277.290 ;
        RECT 281.500 -278.035 281.805 -277.290 ;
        RECT 282.700 -277.860 282.870 -277.080 ;
        RECT 283.190 -277.860 283.360 -277.320 ;
        RECT 283.680 -277.860 283.850 -277.080 ;
        RECT 284.170 -277.860 284.340 -277.320 ;
        RECT 282.110 -278.035 282.475 -278.005 ;
        RECT 281.500 -278.100 282.475 -278.035 ;
        RECT 281.610 -278.240 282.475 -278.100 ;
        RECT 282.110 -278.305 282.475 -278.240 ;
        RECT 284.660 -278.155 286.520 -277.805 ;
        RECT 318.560 -278.035 318.730 -276.995 ;
        RECT 319.540 -278.035 319.710 -276.995 ;
        RECT 320.520 -278.035 320.690 -276.995 ;
        RECT 282.700 -279.015 282.870 -278.475 ;
        RECT 283.680 -279.015 283.850 -278.475 ;
        RECT 284.660 -279.015 284.830 -278.155 ;
        RECT 246.760 -280.805 248.365 -280.635 ;
        RECT 245.865 -283.485 246.035 -280.985 ;
        RECT 245.860 -283.715 246.035 -283.485 ;
        RECT 246.760 -283.715 246.960 -280.805 ;
        RECT 247.205 -281.005 247.380 -280.805 ;
        RECT 247.210 -283.525 247.380 -281.005 ;
        RECT 247.700 -283.490 247.870 -280.985 ;
        RECT 248.190 -281.000 248.365 -280.805 ;
        RECT 245.860 -283.915 246.960 -283.715 ;
        RECT 247.685 -284.090 247.875 -283.490 ;
        RECT 248.190 -283.525 248.360 -281.000 ;
        RECT 248.840 -283.905 249.010 -280.985 ;
        RECT 250.470 -283.555 250.640 -280.985 ;
        RECT 251.610 -282.435 251.780 -280.985 ;
        RECT 282.930 -281.355 284.130 -281.185 ;
        RECT 251.605 -282.900 251.790 -282.435 ;
        RECT 251.605 -283.085 252.290 -282.900 ;
        RECT 250.470 -283.725 251.265 -283.555 ;
        RECT 249.585 -283.905 250.275 -283.850 ;
        RECT 245.865 -284.280 247.875 -284.090 ;
        RECT 248.210 -284.075 250.275 -283.905 ;
        RECT 244.680 -284.335 245.370 -284.285 ;
        RECT 242.730 -284.505 245.370 -284.335 ;
        RECT 240.125 -285.370 240.650 -285.010 ;
        RECT 242.730 -285.885 242.945 -284.505 ;
        RECT 244.680 -284.555 245.370 -284.505 ;
        RECT 244.960 -285.010 245.650 -284.965 ;
        RECT 243.910 -285.180 245.650 -285.010 ;
        RECT 243.910 -285.815 244.270 -285.180 ;
        RECT 244.960 -285.235 245.650 -285.180 ;
        RECT 243.910 -285.860 244.330 -285.815 ;
        RECT 230.290 -286.625 232.540 -286.535 ;
        RECT 228.080 -286.840 232.540 -286.625 ;
        RECT 228.080 -286.930 230.325 -286.840 ;
        RECT 232.235 -288.315 232.540 -286.840 ;
        RECT 235.905 -287.725 236.075 -286.255 ;
        RECT 236.365 -286.335 236.590 -285.985 ;
        RECT 238.325 -286.085 242.945 -285.885 ;
        RECT 238.565 -286.100 242.945 -286.085 ;
        RECT 235.870 -288.315 236.105 -287.725 ;
        RECT 236.395 -287.795 236.565 -286.335 ;
        RECT 236.885 -287.720 237.055 -286.255 ;
        RECT 238.095 -287.670 238.265 -286.255 ;
        RECT 238.565 -286.300 238.785 -286.100 ;
        RECT 243.935 -286.210 244.330 -285.860 ;
        RECT 236.850 -288.315 237.085 -287.720 ;
        RECT 238.060 -288.315 238.295 -287.670 ;
        RECT 238.585 -287.795 238.755 -286.300 ;
        RECT 245.375 -287.420 245.545 -285.965 ;
        RECT 245.365 -287.975 245.550 -287.420 ;
        RECT 245.865 -287.505 246.035 -284.280 ;
        RECT 247.010 -284.630 247.200 -284.280 ;
        RECT 248.210 -284.470 248.380 -284.075 ;
        RECT 249.585 -284.120 250.275 -284.075 ;
        RECT 246.960 -285.320 247.230 -284.630 ;
        RECT 247.725 -284.640 248.380 -284.470 ;
        RECT 248.710 -284.555 249.400 -284.285 ;
        RECT 250.635 -284.630 250.905 -283.940 ;
        RECT 251.095 -283.945 251.265 -283.725 ;
        RECT 251.095 -284.215 251.925 -283.945 ;
        RECT 247.725 -287.505 247.895 -284.640 ;
        RECT 251.095 -284.790 251.265 -284.215 ;
        RECT 251.525 -284.790 251.795 -284.705 ;
        RECT 248.215 -284.985 249.010 -284.810 ;
        RECT 251.095 -284.815 251.795 -284.790 ;
        RECT 250.955 -284.960 251.795 -284.815 ;
        RECT 248.215 -287.505 248.385 -284.985 ;
        RECT 248.840 -287.505 249.010 -284.985 ;
        RECT 249.330 -287.420 249.500 -284.965 ;
        RECT 249.980 -287.415 250.150 -284.965 ;
        RECT 242.680 -287.995 245.735 -287.975 ;
        RECT 249.325 -287.995 249.510 -287.420 ;
        RECT 249.965 -287.995 250.150 -287.415 ;
        RECT 250.470 -287.505 250.640 -284.965 ;
        RECT 250.955 -284.985 251.265 -284.960 ;
        RECT 250.960 -287.505 251.130 -284.985 ;
        RECT 251.525 -285.000 251.795 -284.960 ;
        RECT 252.100 -285.550 252.290 -283.085 ;
        RECT 274.660 -283.690 274.830 -281.970 ;
        RECT 275.640 -283.690 275.810 -281.970 ;
        RECT 277.705 -282.505 277.875 -281.965 ;
        RECT 278.685 -282.505 278.855 -281.965 ;
        RECT 277.115 -282.740 277.480 -282.675 ;
        RECT 276.615 -282.880 277.480 -282.740 ;
        RECT 276.505 -282.945 277.480 -282.880 ;
        RECT 276.505 -283.690 276.810 -282.945 ;
        RECT 277.115 -282.975 277.480 -282.945 ;
        RECT 279.665 -282.825 279.835 -281.965 ;
        RECT 274.660 -283.840 276.810 -283.690 ;
        RECT 274.660 -283.880 276.755 -283.840 ;
        RECT 277.705 -283.900 277.875 -283.120 ;
        RECT 278.195 -283.660 278.365 -283.120 ;
        RECT 278.685 -283.900 278.855 -283.120 ;
        RECT 279.175 -283.660 279.345 -283.120 ;
        RECT 279.665 -283.175 281.055 -282.825 ;
        RECT 272.880 -284.245 274.015 -284.235 ;
        RECT 276.070 -284.245 276.440 -284.115 ;
        RECT 272.880 -284.435 276.440 -284.245 ;
        RECT 277.005 -284.330 280.080 -283.900 ;
        RECT 252.100 -285.740 253.560 -285.550 ;
        RECT 251.610 -287.410 251.780 -285.965 ;
        RECT 252.100 -285.990 252.290 -285.740 ;
        RECT 251.600 -287.995 251.785 -287.410 ;
        RECT 252.100 -287.505 252.270 -285.990 ;
        RECT 242.680 -288.315 252.350 -287.995 ;
        RECT 232.235 -288.540 252.350 -288.315 ;
        RECT 232.235 -288.880 243.245 -288.540 ;
        RECT 244.985 -288.800 252.350 -288.540 ;
        RECT 182.630 -290.430 199.180 -290.050 ;
        RECT 182.630 -291.340 183.010 -290.430 ;
        RECT 182.630 -291.720 183.340 -291.340 ;
        RECT 182.960 -293.665 183.340 -291.720 ;
        RECT 188.005 -291.550 191.330 -291.410 ;
        RECT 188.005 -291.840 193.180 -291.550 ;
        RECT 197.050 -291.835 197.510 -291.410 ;
        RECT 188.005 -292.245 188.435 -291.840 ;
        RECT 189.305 -292.025 189.480 -291.840 ;
        RECT 190.930 -291.855 193.180 -291.840 ;
        RECT 183.745 -292.675 188.435 -292.245 ;
        RECT 182.960 -294.125 183.635 -293.665 ;
        RECT 184.445 -293.955 184.615 -292.675 ;
        RECT 184.935 -293.955 185.105 -292.915 ;
        RECT 185.425 -293.955 185.595 -292.675 ;
        RECT 185.915 -293.785 186.085 -292.915 ;
        RECT 188.820 -293.565 188.990 -292.025 ;
        RECT 189.310 -293.565 189.480 -292.025 ;
        RECT 189.800 -293.565 189.970 -292.025 ;
        RECT 190.290 -293.565 190.460 -292.025 ;
        RECT 190.780 -293.565 190.950 -292.025 ;
        RECT 188.660 -293.780 189.015 -293.775 ;
        RECT 190.720 -293.780 191.090 -293.750 ;
        RECT 188.660 -293.785 191.090 -293.780 ;
        RECT 185.915 -293.955 191.090 -293.785 ;
        RECT 192.875 -293.890 193.180 -291.855 ;
        RECT 185.920 -293.975 191.090 -293.955 ;
        RECT 185.920 -293.985 188.665 -293.975 ;
        RECT 183.855 -294.125 184.220 -294.095 ;
        RECT 190.720 -294.105 191.090 -293.975 ;
        RECT 182.960 -294.210 184.220 -294.125 ;
        RECT 182.985 -294.330 184.220 -294.210 ;
        RECT 188.395 -294.265 189.070 -294.225 ;
        RECT 188.295 -294.275 189.070 -294.265 ;
        RECT 182.985 -294.415 183.635 -294.330 ;
        RECT 183.855 -294.395 184.220 -294.330 ;
        RECT 187.260 -294.455 189.070 -294.275 ;
        RECT 191.655 -294.320 195.580 -293.890 ;
        RECT 188.295 -294.465 189.070 -294.455 ;
        RECT 188.395 -294.495 189.070 -294.465 ;
        RECT 189.310 -294.380 191.405 -294.340 ;
        RECT 189.310 -294.530 191.460 -294.380 ;
        RECT 184.445 -295.605 184.615 -294.565 ;
        RECT 185.425 -295.605 185.595 -294.565 ;
        RECT 186.405 -295.605 186.575 -294.565 ;
        RECT 189.310 -296.250 189.480 -294.530 ;
        RECT 190.290 -296.250 190.460 -294.530 ;
        RECT 191.155 -295.275 191.460 -294.530 ;
        RECT 192.355 -295.100 192.525 -294.320 ;
        RECT 192.845 -295.100 193.015 -294.560 ;
        RECT 193.335 -295.100 193.505 -294.320 ;
        RECT 193.825 -295.100 193.995 -294.560 ;
        RECT 191.765 -295.275 192.130 -295.245 ;
        RECT 191.155 -295.340 192.130 -295.275 ;
        RECT 191.265 -295.480 192.130 -295.340 ;
        RECT 191.765 -295.545 192.130 -295.480 ;
        RECT 194.315 -295.395 196.175 -295.045 ;
        RECT 192.355 -296.255 192.525 -295.715 ;
        RECT 193.335 -296.255 193.505 -295.715 ;
        RECT 194.315 -296.255 194.485 -295.395 ;
        RECT 192.585 -298.595 193.785 -298.425 ;
        RECT 184.315 -300.930 184.485 -299.210 ;
        RECT 185.295 -300.930 185.465 -299.210 ;
        RECT 187.360 -299.745 187.530 -299.205 ;
        RECT 188.340 -299.745 188.510 -299.205 ;
        RECT 186.770 -299.980 187.135 -299.915 ;
        RECT 186.270 -300.120 187.135 -299.980 ;
        RECT 186.160 -300.185 187.135 -300.120 ;
        RECT 186.160 -300.930 186.465 -300.185 ;
        RECT 186.770 -300.215 187.135 -300.185 ;
        RECT 189.320 -300.065 189.490 -299.205 ;
        RECT 184.315 -301.080 186.465 -300.930 ;
        RECT 184.315 -301.120 186.410 -301.080 ;
        RECT 187.360 -301.140 187.530 -300.360 ;
        RECT 187.850 -300.900 188.020 -300.360 ;
        RECT 188.340 -301.140 188.510 -300.360 ;
        RECT 188.830 -300.900 189.000 -300.360 ;
        RECT 189.320 -300.415 190.710 -300.065 ;
        RECT 182.535 -301.485 183.670 -301.475 ;
        RECT 185.725 -301.485 186.095 -301.355 ;
        RECT 182.535 -301.675 186.095 -301.485 ;
        RECT 186.660 -301.570 189.735 -301.140 ;
        RECT 183.665 -301.680 186.095 -301.675 ;
        RECT 183.665 -301.685 184.020 -301.680 ;
        RECT 185.725 -301.710 186.095 -301.680 ;
        RECT 183.825 -303.435 183.995 -301.895 ;
        RECT 184.315 -303.435 184.485 -301.895 ;
        RECT 184.805 -303.435 184.975 -301.895 ;
        RECT 185.295 -303.435 185.465 -301.895 ;
        RECT 185.785 -303.435 185.955 -301.895 ;
        RECT 184.310 -303.695 184.485 -303.435 ;
        RECT 187.880 -303.605 188.185 -301.570 ;
        RECT 190.330 -302.390 190.680 -300.415 ;
        RECT 191.550 -301.685 191.720 -298.765 ;
        RECT 192.585 -298.805 192.795 -298.595 ;
        RECT 191.530 -301.980 191.740 -301.685 ;
        RECT 192.605 -301.715 192.775 -298.805 ;
        RECT 193.095 -301.705 193.265 -298.765 ;
        RECT 193.575 -298.815 193.785 -298.595 ;
        RECT 192.590 -301.980 192.800 -301.715 ;
        RECT 191.530 -302.160 192.800 -301.980 ;
        RECT 193.075 -301.975 193.285 -301.705 ;
        RECT 193.585 -301.805 193.755 -298.815 ;
        RECT 194.645 -301.735 194.815 -298.765 ;
        RECT 193.075 -302.170 193.780 -301.975 ;
        RECT 193.565 -302.230 193.780 -302.170 ;
        RECT 192.355 -302.390 193.130 -302.340 ;
        RECT 190.330 -302.570 193.130 -302.390 ;
        RECT 190.330 -302.580 190.680 -302.570 ;
        RECT 192.355 -302.615 193.130 -302.570 ;
        RECT 193.565 -302.505 194.470 -302.230 ;
        RECT 193.565 -302.855 193.780 -302.505 ;
        RECT 191.005 -302.925 191.780 -302.880 ;
        RECT 190.820 -303.095 191.780 -302.925 ;
        RECT 191.005 -303.155 191.780 -303.095 ;
        RECT 192.010 -303.055 193.780 -302.855 ;
        RECT 194.640 -302.955 194.855 -301.735 ;
        RECT 195.825 -302.080 196.175 -295.395 ;
        RECT 197.165 -301.710 197.380 -291.835 ;
        RECT 198.800 -293.950 199.180 -290.430 ;
        RECT 200.310 -290.210 209.245 -290.020 ;
        RECT 223.695 -290.025 227.325 -289.295 ;
        RECT 200.310 -292.100 200.500 -290.210 ;
        RECT 206.345 -291.705 209.670 -291.565 ;
        RECT 206.345 -291.995 211.520 -291.705 ;
        RECT 200.195 -292.370 200.560 -292.100 ;
        RECT 206.345 -292.400 206.775 -291.995 ;
        RECT 207.645 -292.180 207.820 -291.995 ;
        RECT 209.270 -292.010 211.520 -291.995 ;
        RECT 202.085 -292.830 206.775 -292.400 ;
        RECT 201.325 -293.950 201.975 -293.820 ;
        RECT 198.800 -294.280 201.975 -293.950 ;
        RECT 202.785 -294.110 202.955 -292.830 ;
        RECT 203.275 -294.110 203.445 -293.070 ;
        RECT 203.765 -294.110 203.935 -292.830 ;
        RECT 204.255 -293.940 204.425 -293.070 ;
        RECT 207.160 -293.720 207.330 -292.180 ;
        RECT 207.650 -293.720 207.820 -292.180 ;
        RECT 208.140 -293.720 208.310 -292.180 ;
        RECT 208.630 -293.720 208.800 -292.180 ;
        RECT 209.120 -293.720 209.290 -292.180 ;
        RECT 207.000 -293.935 207.355 -293.930 ;
        RECT 209.060 -293.935 209.430 -293.905 ;
        RECT 207.000 -293.940 209.430 -293.935 ;
        RECT 204.255 -294.110 209.430 -293.940 ;
        RECT 211.215 -294.045 211.520 -292.010 ;
        RECT 204.260 -294.130 209.430 -294.110 ;
        RECT 204.260 -294.140 207.005 -294.130 ;
        RECT 202.195 -294.280 202.560 -294.250 ;
        RECT 209.060 -294.260 209.430 -294.130 ;
        RECT 198.800 -294.330 202.560 -294.280 ;
        RECT 201.325 -294.485 202.560 -294.330 ;
        RECT 206.735 -294.420 207.410 -294.380 ;
        RECT 206.635 -294.430 207.410 -294.420 ;
        RECT 201.325 -294.570 201.975 -294.485 ;
        RECT 202.195 -294.550 202.560 -294.485 ;
        RECT 201.460 -294.820 201.840 -294.570 ;
        RECT 205.600 -294.610 207.410 -294.430 ;
        RECT 209.995 -294.475 213.920 -294.045 ;
        RECT 206.635 -294.620 207.410 -294.610 ;
        RECT 206.735 -294.650 207.410 -294.620 ;
        RECT 207.650 -294.535 209.745 -294.495 ;
        RECT 207.650 -294.685 209.800 -294.535 ;
        RECT 202.785 -295.760 202.955 -294.720 ;
        RECT 203.765 -295.760 203.935 -294.720 ;
        RECT 204.745 -295.760 204.915 -294.720 ;
        RECT 207.650 -296.405 207.820 -294.685 ;
        RECT 208.630 -296.405 208.800 -294.685 ;
        RECT 209.495 -295.430 209.800 -294.685 ;
        RECT 210.695 -295.255 210.865 -294.475 ;
        RECT 211.185 -295.255 211.355 -294.715 ;
        RECT 211.675 -295.255 211.845 -294.475 ;
        RECT 212.165 -295.255 212.335 -294.715 ;
        RECT 210.105 -295.430 210.470 -295.400 ;
        RECT 209.495 -295.495 210.470 -295.430 ;
        RECT 209.605 -295.635 210.470 -295.495 ;
        RECT 210.105 -295.700 210.470 -295.635 ;
        RECT 212.655 -295.550 214.515 -295.200 ;
        RECT 210.695 -296.410 210.865 -295.870 ;
        RECT 211.675 -296.410 211.845 -295.870 ;
        RECT 212.655 -296.410 212.825 -295.550 ;
        RECT 210.925 -298.750 212.125 -298.580 ;
        RECT 202.655 -301.085 202.825 -299.365 ;
        RECT 203.635 -301.085 203.805 -299.365 ;
        RECT 205.700 -299.900 205.870 -299.360 ;
        RECT 206.680 -299.900 206.850 -299.360 ;
        RECT 205.110 -300.135 205.475 -300.070 ;
        RECT 204.610 -300.275 205.475 -300.135 ;
        RECT 204.500 -300.340 205.475 -300.275 ;
        RECT 204.500 -301.085 204.805 -300.340 ;
        RECT 205.110 -300.370 205.475 -300.340 ;
        RECT 207.660 -300.220 207.830 -299.360 ;
        RECT 202.655 -301.235 204.805 -301.085 ;
        RECT 202.655 -301.275 204.750 -301.235 ;
        RECT 205.700 -301.295 205.870 -300.515 ;
        RECT 206.190 -301.055 206.360 -300.515 ;
        RECT 206.680 -301.295 206.850 -300.515 ;
        RECT 207.170 -301.055 207.340 -300.515 ;
        RECT 207.660 -300.570 209.050 -300.220 ;
        RECT 200.875 -301.640 202.010 -301.630 ;
        RECT 204.065 -301.640 204.435 -301.510 ;
        RECT 197.165 -301.925 198.590 -301.710 ;
        RECT 200.875 -301.830 204.435 -301.640 ;
        RECT 205.000 -301.725 208.075 -301.295 ;
        RECT 202.005 -301.835 204.435 -301.830 ;
        RECT 202.005 -301.840 202.360 -301.835 ;
        RECT 204.065 -301.865 204.435 -301.835 ;
        RECT 195.770 -302.440 196.295 -302.080 ;
        RECT 198.375 -302.955 198.590 -301.925 ;
        RECT 185.935 -303.695 188.185 -303.605 ;
        RECT 183.725 -303.910 188.185 -303.695 ;
        RECT 183.725 -304.000 185.970 -303.910 ;
        RECT 187.880 -305.385 188.185 -303.910 ;
        RECT 191.550 -304.795 191.720 -303.325 ;
        RECT 192.010 -303.405 192.235 -303.055 ;
        RECT 193.970 -303.155 198.590 -302.955 ;
        RECT 194.210 -303.170 198.590 -303.155 ;
        RECT 191.515 -305.385 191.750 -304.795 ;
        RECT 192.040 -304.865 192.210 -303.405 ;
        RECT 192.530 -304.790 192.700 -303.325 ;
        RECT 193.740 -304.740 193.910 -303.325 ;
        RECT 194.210 -303.370 194.430 -303.170 ;
        RECT 192.495 -305.385 192.730 -304.790 ;
        RECT 193.705 -305.385 193.940 -304.740 ;
        RECT 194.230 -304.865 194.400 -303.370 ;
        RECT 202.165 -303.590 202.335 -302.050 ;
        RECT 202.655 -303.590 202.825 -302.050 ;
        RECT 203.145 -303.590 203.315 -302.050 ;
        RECT 203.635 -303.590 203.805 -302.050 ;
        RECT 204.125 -303.590 204.295 -302.050 ;
        RECT 202.650 -303.850 202.825 -303.590 ;
        RECT 206.220 -303.760 206.525 -301.725 ;
        RECT 208.670 -302.545 209.020 -300.570 ;
        RECT 209.890 -301.840 210.060 -298.920 ;
        RECT 210.925 -298.960 211.135 -298.750 ;
        RECT 209.870 -302.135 210.080 -301.840 ;
        RECT 210.945 -301.870 211.115 -298.960 ;
        RECT 211.435 -301.860 211.605 -298.920 ;
        RECT 211.915 -298.970 212.125 -298.750 ;
        RECT 210.930 -302.135 211.140 -301.870 ;
        RECT 209.870 -302.315 211.140 -302.135 ;
        RECT 211.415 -302.130 211.625 -301.860 ;
        RECT 211.925 -301.960 212.095 -298.970 ;
        RECT 212.985 -301.890 213.155 -298.920 ;
        RECT 211.415 -302.325 212.120 -302.130 ;
        RECT 211.905 -302.385 212.120 -302.325 ;
        RECT 210.695 -302.545 211.470 -302.495 ;
        RECT 208.670 -302.725 211.470 -302.545 ;
        RECT 208.670 -302.735 209.020 -302.725 ;
        RECT 210.695 -302.770 211.470 -302.725 ;
        RECT 211.905 -302.660 212.810 -302.385 ;
        RECT 211.905 -303.010 212.120 -302.660 ;
        RECT 209.345 -303.080 210.120 -303.035 ;
        RECT 209.160 -303.250 210.120 -303.080 ;
        RECT 209.345 -303.310 210.120 -303.250 ;
        RECT 210.350 -303.210 212.120 -303.010 ;
        RECT 212.980 -303.110 213.195 -301.890 ;
        RECT 214.165 -302.235 214.515 -295.550 ;
        RECT 214.110 -302.595 214.635 -302.235 ;
        RECT 216.685 -303.110 218.370 -302.295 ;
        RECT 204.275 -303.850 206.525 -303.760 ;
        RECT 202.065 -304.065 206.525 -303.850 ;
        RECT 202.065 -304.155 204.310 -304.065 ;
        RECT 187.880 -305.950 195.265 -305.385 ;
        RECT 206.220 -305.540 206.525 -304.065 ;
        RECT 209.890 -304.950 210.060 -303.480 ;
        RECT 210.350 -303.560 210.575 -303.210 ;
        RECT 212.310 -303.310 218.370 -303.110 ;
        RECT 212.550 -303.325 218.370 -303.310 ;
        RECT 209.855 -305.540 210.090 -304.950 ;
        RECT 210.380 -305.020 210.550 -303.560 ;
        RECT 210.870 -304.945 211.040 -303.480 ;
        RECT 212.080 -304.895 212.250 -303.480 ;
        RECT 212.550 -303.525 212.770 -303.325 ;
        RECT 210.835 -305.540 211.070 -304.945 ;
        RECT 212.045 -305.540 212.280 -304.895 ;
        RECT 212.570 -305.020 212.740 -303.525 ;
        RECT 216.685 -303.950 218.370 -303.325 ;
        RECT 206.220 -306.105 213.605 -305.540 ;
        RECT 179.235 -310.040 180.250 -309.305 ;
        RECT 127.120 -310.050 136.895 -310.045 ;
        RECT 214.890 -310.210 216.475 -308.755 ;
        RECT 223.695 -310.030 224.425 -290.025 ;
        RECT 226.945 -290.245 227.325 -290.025 ;
        RECT 253.370 -290.215 253.560 -285.740 ;
        RECT 272.935 -288.790 273.315 -284.435 ;
        RECT 274.010 -284.440 276.440 -284.435 ;
        RECT 274.010 -284.445 274.365 -284.440 ;
        RECT 276.070 -284.470 276.440 -284.440 ;
        RECT 274.170 -286.195 274.340 -284.655 ;
        RECT 274.660 -286.195 274.830 -284.655 ;
        RECT 275.150 -286.195 275.320 -284.655 ;
        RECT 275.640 -286.195 275.810 -284.655 ;
        RECT 276.130 -286.195 276.300 -284.655 ;
        RECT 274.655 -286.455 274.830 -286.195 ;
        RECT 278.225 -286.365 278.530 -284.330 ;
        RECT 280.675 -285.150 281.025 -283.175 ;
        RECT 281.895 -284.445 282.065 -281.525 ;
        RECT 282.930 -281.565 283.140 -281.355 ;
        RECT 281.875 -284.740 282.085 -284.445 ;
        RECT 282.950 -284.475 283.120 -281.565 ;
        RECT 283.440 -284.465 283.610 -281.525 ;
        RECT 283.920 -281.575 284.130 -281.355 ;
        RECT 282.935 -284.740 283.145 -284.475 ;
        RECT 281.875 -284.920 283.145 -284.740 ;
        RECT 283.420 -284.735 283.630 -284.465 ;
        RECT 283.930 -284.565 284.100 -281.575 ;
        RECT 284.990 -284.495 285.160 -281.525 ;
        RECT 283.420 -284.930 284.125 -284.735 ;
        RECT 283.910 -284.990 284.125 -284.930 ;
        RECT 282.700 -285.150 283.475 -285.100 ;
        RECT 280.675 -285.330 283.475 -285.150 ;
        RECT 280.675 -285.340 281.025 -285.330 ;
        RECT 282.700 -285.375 283.475 -285.330 ;
        RECT 283.910 -285.265 284.815 -284.990 ;
        RECT 283.910 -285.615 284.125 -285.265 ;
        RECT 281.350 -285.685 282.125 -285.640 ;
        RECT 281.165 -285.855 282.125 -285.685 ;
        RECT 281.350 -285.915 282.125 -285.855 ;
        RECT 282.355 -285.815 284.125 -285.615 ;
        RECT 284.985 -285.715 285.200 -284.495 ;
        RECT 286.170 -284.840 286.520 -278.155 ;
        RECT 323.425 -278.680 323.595 -276.960 ;
        RECT 324.405 -278.680 324.575 -276.960 ;
        RECT 325.270 -277.705 325.575 -276.960 ;
        RECT 326.470 -277.530 326.640 -276.750 ;
        RECT 326.960 -277.530 327.130 -276.990 ;
        RECT 327.450 -277.530 327.620 -276.750 ;
        RECT 362.865 -276.760 363.515 -276.675 ;
        RECT 363.735 -276.740 364.100 -276.675 ;
        RECT 367.140 -276.800 368.950 -276.620 ;
        RECT 371.535 -276.665 375.460 -276.235 ;
        RECT 409.685 -276.280 410.335 -275.820 ;
        RECT 411.145 -276.110 411.315 -274.830 ;
        RECT 411.635 -276.110 411.805 -275.070 ;
        RECT 412.125 -276.110 412.295 -274.830 ;
        RECT 412.615 -275.940 412.785 -275.070 ;
        RECT 415.520 -275.720 415.690 -274.180 ;
        RECT 416.010 -275.720 416.180 -274.180 ;
        RECT 416.500 -275.720 416.670 -274.180 ;
        RECT 416.990 -275.720 417.160 -274.180 ;
        RECT 417.480 -275.720 417.650 -274.180 ;
        RECT 415.360 -275.935 415.715 -275.930 ;
        RECT 417.420 -275.935 417.790 -275.905 ;
        RECT 415.360 -275.940 417.790 -275.935 ;
        RECT 412.615 -276.110 417.790 -275.940 ;
        RECT 419.575 -276.045 419.880 -274.010 ;
        RECT 412.620 -276.130 417.790 -276.110 ;
        RECT 412.620 -276.140 415.365 -276.130 ;
        RECT 410.555 -276.280 410.920 -276.250 ;
        RECT 417.420 -276.260 417.790 -276.130 ;
        RECT 409.685 -276.485 410.920 -276.280 ;
        RECT 415.095 -276.420 415.770 -276.380 ;
        RECT 414.995 -276.430 415.770 -276.420 ;
        RECT 409.685 -276.570 410.335 -276.485 ;
        RECT 410.555 -276.550 410.920 -276.485 ;
        RECT 413.960 -276.610 415.770 -276.430 ;
        RECT 418.355 -276.475 422.280 -276.045 ;
        RECT 414.995 -276.620 415.770 -276.610 ;
        RECT 415.095 -276.650 415.770 -276.620 ;
        RECT 416.010 -276.535 418.105 -276.495 ;
        RECT 368.175 -276.810 368.950 -276.800 ;
        RECT 368.275 -276.840 368.950 -276.810 ;
        RECT 369.190 -276.725 371.285 -276.685 ;
        RECT 369.190 -276.875 371.340 -276.725 ;
        RECT 327.940 -277.530 328.110 -276.990 ;
        RECT 325.880 -277.705 326.245 -277.675 ;
        RECT 325.270 -277.770 326.245 -277.705 ;
        RECT 325.380 -277.910 326.245 -277.770 ;
        RECT 325.880 -277.975 326.245 -277.910 ;
        RECT 328.430 -277.825 330.290 -277.475 ;
        RECT 326.470 -278.685 326.640 -278.145 ;
        RECT 327.450 -278.685 327.620 -278.145 ;
        RECT 328.430 -278.685 328.600 -277.825 ;
        RECT 292.750 -280.635 294.355 -280.465 ;
        RECT 291.855 -283.315 292.025 -280.815 ;
        RECT 291.850 -283.545 292.025 -283.315 ;
        RECT 292.750 -283.545 292.950 -280.635 ;
        RECT 293.195 -280.835 293.370 -280.635 ;
        RECT 293.200 -283.355 293.370 -280.835 ;
        RECT 293.690 -283.320 293.860 -280.815 ;
        RECT 294.180 -280.830 294.355 -280.635 ;
        RECT 291.850 -283.745 292.950 -283.545 ;
        RECT 293.675 -283.920 293.865 -283.320 ;
        RECT 294.180 -283.355 294.350 -280.830 ;
        RECT 294.830 -283.735 295.000 -280.815 ;
        RECT 296.460 -283.385 296.630 -280.815 ;
        RECT 297.600 -282.265 297.770 -280.815 ;
        RECT 326.700 -281.025 327.900 -280.855 ;
        RECT 297.595 -282.730 297.780 -282.265 ;
        RECT 297.595 -282.915 298.280 -282.730 ;
        RECT 296.460 -283.555 297.255 -283.385 ;
        RECT 295.575 -283.735 296.265 -283.680 ;
        RECT 291.855 -284.110 293.865 -283.920 ;
        RECT 294.200 -283.905 296.265 -283.735 ;
        RECT 290.670 -284.165 291.360 -284.115 ;
        RECT 288.720 -284.335 291.360 -284.165 ;
        RECT 286.115 -285.200 286.640 -284.840 ;
        RECT 288.720 -285.715 288.935 -284.335 ;
        RECT 290.670 -284.385 291.360 -284.335 ;
        RECT 290.950 -284.840 291.640 -284.795 ;
        RECT 289.900 -285.010 291.640 -284.840 ;
        RECT 289.900 -285.645 290.260 -285.010 ;
        RECT 290.950 -285.065 291.640 -285.010 ;
        RECT 289.900 -285.690 290.320 -285.645 ;
        RECT 276.280 -286.455 278.530 -286.365 ;
        RECT 274.070 -286.670 278.530 -286.455 ;
        RECT 274.070 -286.760 276.315 -286.670 ;
        RECT 278.225 -288.145 278.530 -286.670 ;
        RECT 281.895 -287.555 282.065 -286.085 ;
        RECT 282.355 -286.165 282.580 -285.815 ;
        RECT 284.315 -285.915 288.935 -285.715 ;
        RECT 284.555 -285.930 288.935 -285.915 ;
        RECT 281.860 -288.145 282.095 -287.555 ;
        RECT 282.385 -287.625 282.555 -286.165 ;
        RECT 282.875 -287.550 283.045 -286.085 ;
        RECT 284.085 -287.500 284.255 -286.085 ;
        RECT 284.555 -286.130 284.775 -285.930 ;
        RECT 289.925 -286.040 290.320 -285.690 ;
        RECT 282.840 -288.145 283.075 -287.550 ;
        RECT 284.050 -288.145 284.285 -287.500 ;
        RECT 284.575 -287.625 284.745 -286.130 ;
        RECT 291.365 -287.250 291.535 -285.795 ;
        RECT 291.355 -287.805 291.540 -287.250 ;
        RECT 291.855 -287.335 292.025 -284.110 ;
        RECT 293.000 -284.460 293.190 -284.110 ;
        RECT 294.200 -284.300 294.370 -283.905 ;
        RECT 295.575 -283.950 296.265 -283.905 ;
        RECT 292.950 -285.150 293.220 -284.460 ;
        RECT 293.715 -284.470 294.370 -284.300 ;
        RECT 294.700 -284.385 295.390 -284.115 ;
        RECT 296.625 -284.460 296.895 -283.770 ;
        RECT 297.085 -283.775 297.255 -283.555 ;
        RECT 297.085 -284.045 297.915 -283.775 ;
        RECT 293.715 -287.335 293.885 -284.470 ;
        RECT 297.085 -284.620 297.255 -284.045 ;
        RECT 297.515 -284.620 297.785 -284.535 ;
        RECT 294.205 -284.815 295.000 -284.640 ;
        RECT 297.085 -284.645 297.785 -284.620 ;
        RECT 296.945 -284.790 297.785 -284.645 ;
        RECT 294.205 -287.335 294.375 -284.815 ;
        RECT 294.830 -287.335 295.000 -284.815 ;
        RECT 295.320 -287.250 295.490 -284.795 ;
        RECT 295.970 -287.245 296.140 -284.795 ;
        RECT 288.670 -287.825 291.725 -287.805 ;
        RECT 295.315 -287.825 295.500 -287.250 ;
        RECT 295.955 -287.825 296.140 -287.245 ;
        RECT 296.460 -287.335 296.630 -284.795 ;
        RECT 296.945 -284.815 297.255 -284.790 ;
        RECT 296.950 -287.335 297.120 -284.815 ;
        RECT 297.515 -284.830 297.785 -284.790 ;
        RECT 298.090 -285.380 298.280 -282.915 ;
        RECT 318.430 -283.360 318.600 -281.640 ;
        RECT 319.410 -283.360 319.580 -281.640 ;
        RECT 321.475 -282.175 321.645 -281.635 ;
        RECT 322.455 -282.175 322.625 -281.635 ;
        RECT 320.885 -282.410 321.250 -282.345 ;
        RECT 320.385 -282.550 321.250 -282.410 ;
        RECT 320.275 -282.615 321.250 -282.550 ;
        RECT 320.275 -283.360 320.580 -282.615 ;
        RECT 320.885 -282.645 321.250 -282.615 ;
        RECT 323.435 -282.495 323.605 -281.635 ;
        RECT 318.430 -283.510 320.580 -283.360 ;
        RECT 318.430 -283.550 320.525 -283.510 ;
        RECT 321.475 -283.570 321.645 -282.790 ;
        RECT 321.965 -283.330 322.135 -282.790 ;
        RECT 322.455 -283.570 322.625 -282.790 ;
        RECT 322.945 -283.330 323.115 -282.790 ;
        RECT 323.435 -282.845 324.825 -282.495 ;
        RECT 316.650 -283.915 317.785 -283.905 ;
        RECT 319.840 -283.915 320.210 -283.785 ;
        RECT 316.650 -284.105 320.210 -283.915 ;
        RECT 320.775 -284.000 323.850 -283.570 ;
        RECT 298.090 -285.570 299.550 -285.380 ;
        RECT 297.600 -287.240 297.770 -285.795 ;
        RECT 298.090 -285.820 298.280 -285.570 ;
        RECT 297.590 -287.825 297.775 -287.240 ;
        RECT 298.090 -287.335 298.260 -285.820 ;
        RECT 288.670 -288.145 298.340 -287.825 ;
        RECT 278.225 -288.370 298.340 -288.145 ;
        RECT 278.225 -288.710 289.235 -288.370 ;
        RECT 290.975 -288.630 298.340 -288.370 ;
        RECT 226.945 -290.625 243.495 -290.245 ;
        RECT 226.945 -291.535 227.325 -290.625 ;
        RECT 226.945 -291.915 227.655 -291.535 ;
        RECT 227.275 -293.860 227.655 -291.915 ;
        RECT 232.320 -291.745 235.645 -291.605 ;
        RECT 232.320 -292.035 237.495 -291.745 ;
        RECT 241.365 -292.030 241.825 -291.605 ;
        RECT 232.320 -292.440 232.750 -292.035 ;
        RECT 233.620 -292.220 233.795 -292.035 ;
        RECT 235.245 -292.050 237.495 -292.035 ;
        RECT 228.060 -292.870 232.750 -292.440 ;
        RECT 227.275 -294.320 227.950 -293.860 ;
        RECT 228.760 -294.150 228.930 -292.870 ;
        RECT 229.250 -294.150 229.420 -293.110 ;
        RECT 229.740 -294.150 229.910 -292.870 ;
        RECT 230.230 -293.980 230.400 -293.110 ;
        RECT 233.135 -293.760 233.305 -292.220 ;
        RECT 233.625 -293.760 233.795 -292.220 ;
        RECT 234.115 -293.760 234.285 -292.220 ;
        RECT 234.605 -293.760 234.775 -292.220 ;
        RECT 235.095 -293.760 235.265 -292.220 ;
        RECT 232.975 -293.975 233.330 -293.970 ;
        RECT 235.035 -293.975 235.405 -293.945 ;
        RECT 232.975 -293.980 235.405 -293.975 ;
        RECT 230.230 -294.150 235.405 -293.980 ;
        RECT 237.190 -294.085 237.495 -292.050 ;
        RECT 230.235 -294.170 235.405 -294.150 ;
        RECT 230.235 -294.180 232.980 -294.170 ;
        RECT 228.170 -294.320 228.535 -294.290 ;
        RECT 235.035 -294.300 235.405 -294.170 ;
        RECT 227.275 -294.405 228.535 -294.320 ;
        RECT 227.300 -294.525 228.535 -294.405 ;
        RECT 232.710 -294.460 233.385 -294.420 ;
        RECT 232.610 -294.470 233.385 -294.460 ;
        RECT 227.300 -294.610 227.950 -294.525 ;
        RECT 228.170 -294.590 228.535 -294.525 ;
        RECT 231.575 -294.650 233.385 -294.470 ;
        RECT 235.970 -294.515 239.895 -294.085 ;
        RECT 232.610 -294.660 233.385 -294.650 ;
        RECT 232.710 -294.690 233.385 -294.660 ;
        RECT 233.625 -294.575 235.720 -294.535 ;
        RECT 233.625 -294.725 235.775 -294.575 ;
        RECT 228.760 -295.800 228.930 -294.760 ;
        RECT 229.740 -295.800 229.910 -294.760 ;
        RECT 230.720 -295.800 230.890 -294.760 ;
        RECT 233.625 -296.445 233.795 -294.725 ;
        RECT 234.605 -296.445 234.775 -294.725 ;
        RECT 235.470 -295.470 235.775 -294.725 ;
        RECT 236.670 -295.295 236.840 -294.515 ;
        RECT 237.160 -295.295 237.330 -294.755 ;
        RECT 237.650 -295.295 237.820 -294.515 ;
        RECT 238.140 -295.295 238.310 -294.755 ;
        RECT 236.080 -295.470 236.445 -295.440 ;
        RECT 235.470 -295.535 236.445 -295.470 ;
        RECT 235.580 -295.675 236.445 -295.535 ;
        RECT 236.080 -295.740 236.445 -295.675 ;
        RECT 238.630 -295.590 240.490 -295.240 ;
        RECT 236.670 -296.450 236.840 -295.910 ;
        RECT 237.650 -296.450 237.820 -295.910 ;
        RECT 238.630 -296.450 238.800 -295.590 ;
        RECT 236.900 -298.790 238.100 -298.620 ;
        RECT 228.630 -301.125 228.800 -299.405 ;
        RECT 229.610 -301.125 229.780 -299.405 ;
        RECT 231.675 -299.940 231.845 -299.400 ;
        RECT 232.655 -299.940 232.825 -299.400 ;
        RECT 231.085 -300.175 231.450 -300.110 ;
        RECT 230.585 -300.315 231.450 -300.175 ;
        RECT 230.475 -300.380 231.450 -300.315 ;
        RECT 230.475 -301.125 230.780 -300.380 ;
        RECT 231.085 -300.410 231.450 -300.380 ;
        RECT 233.635 -300.260 233.805 -299.400 ;
        RECT 228.630 -301.275 230.780 -301.125 ;
        RECT 228.630 -301.315 230.725 -301.275 ;
        RECT 231.675 -301.335 231.845 -300.555 ;
        RECT 232.165 -301.095 232.335 -300.555 ;
        RECT 232.655 -301.335 232.825 -300.555 ;
        RECT 233.145 -301.095 233.315 -300.555 ;
        RECT 233.635 -300.610 235.025 -300.260 ;
        RECT 226.850 -301.680 227.985 -301.670 ;
        RECT 230.040 -301.680 230.410 -301.550 ;
        RECT 226.850 -301.870 230.410 -301.680 ;
        RECT 230.975 -301.765 234.050 -301.335 ;
        RECT 227.980 -301.875 230.410 -301.870 ;
        RECT 227.980 -301.880 228.335 -301.875 ;
        RECT 230.040 -301.905 230.410 -301.875 ;
        RECT 228.140 -303.630 228.310 -302.090 ;
        RECT 228.630 -303.630 228.800 -302.090 ;
        RECT 229.120 -303.630 229.290 -302.090 ;
        RECT 229.610 -303.630 229.780 -302.090 ;
        RECT 230.100 -303.630 230.270 -302.090 ;
        RECT 228.625 -303.890 228.800 -303.630 ;
        RECT 232.195 -303.800 232.500 -301.765 ;
        RECT 234.645 -302.585 234.995 -300.610 ;
        RECT 235.865 -301.880 236.035 -298.960 ;
        RECT 236.900 -299.000 237.110 -298.790 ;
        RECT 235.845 -302.175 236.055 -301.880 ;
        RECT 236.920 -301.910 237.090 -299.000 ;
        RECT 237.410 -301.900 237.580 -298.960 ;
        RECT 237.890 -299.010 238.100 -298.790 ;
        RECT 236.905 -302.175 237.115 -301.910 ;
        RECT 235.845 -302.355 237.115 -302.175 ;
        RECT 237.390 -302.170 237.600 -301.900 ;
        RECT 237.900 -302.000 238.070 -299.010 ;
        RECT 238.960 -301.930 239.130 -298.960 ;
        RECT 237.390 -302.365 238.095 -302.170 ;
        RECT 237.880 -302.425 238.095 -302.365 ;
        RECT 236.670 -302.585 237.445 -302.535 ;
        RECT 234.645 -302.765 237.445 -302.585 ;
        RECT 234.645 -302.775 234.995 -302.765 ;
        RECT 236.670 -302.810 237.445 -302.765 ;
        RECT 237.880 -302.700 238.785 -302.425 ;
        RECT 237.880 -303.050 238.095 -302.700 ;
        RECT 235.320 -303.120 236.095 -303.075 ;
        RECT 235.135 -303.290 236.095 -303.120 ;
        RECT 235.320 -303.350 236.095 -303.290 ;
        RECT 236.325 -303.250 238.095 -303.050 ;
        RECT 238.955 -303.150 239.170 -301.930 ;
        RECT 240.140 -302.275 240.490 -295.590 ;
        RECT 241.480 -301.905 241.695 -292.030 ;
        RECT 243.115 -294.145 243.495 -290.625 ;
        RECT 244.625 -290.405 253.560 -290.215 ;
        RECT 269.380 -289.595 273.315 -288.790 ;
        RECT 244.625 -292.295 244.815 -290.405 ;
        RECT 250.660 -291.900 253.985 -291.760 ;
        RECT 250.660 -292.190 255.835 -291.900 ;
        RECT 244.510 -292.565 244.875 -292.295 ;
        RECT 250.660 -292.595 251.090 -292.190 ;
        RECT 251.960 -292.375 252.135 -292.190 ;
        RECT 253.585 -292.205 255.835 -292.190 ;
        RECT 246.400 -293.025 251.090 -292.595 ;
        RECT 245.640 -294.145 246.290 -294.015 ;
        RECT 243.115 -294.475 246.290 -294.145 ;
        RECT 247.100 -294.305 247.270 -293.025 ;
        RECT 247.590 -294.305 247.760 -293.265 ;
        RECT 248.080 -294.305 248.250 -293.025 ;
        RECT 248.570 -294.135 248.740 -293.265 ;
        RECT 251.475 -293.915 251.645 -292.375 ;
        RECT 251.965 -293.915 252.135 -292.375 ;
        RECT 252.455 -293.915 252.625 -292.375 ;
        RECT 252.945 -293.915 253.115 -292.375 ;
        RECT 253.435 -293.915 253.605 -292.375 ;
        RECT 251.315 -294.130 251.670 -294.125 ;
        RECT 253.375 -294.130 253.745 -294.100 ;
        RECT 251.315 -294.135 253.745 -294.130 ;
        RECT 248.570 -294.305 253.745 -294.135 ;
        RECT 255.530 -294.240 255.835 -292.205 ;
        RECT 248.575 -294.325 253.745 -294.305 ;
        RECT 248.575 -294.335 251.320 -294.325 ;
        RECT 246.510 -294.475 246.875 -294.445 ;
        RECT 253.375 -294.455 253.745 -294.325 ;
        RECT 243.115 -294.525 246.875 -294.475 ;
        RECT 245.640 -294.680 246.875 -294.525 ;
        RECT 251.050 -294.615 251.725 -294.575 ;
        RECT 250.950 -294.625 251.725 -294.615 ;
        RECT 245.640 -294.765 246.290 -294.680 ;
        RECT 246.510 -294.745 246.875 -294.680 ;
        RECT 245.775 -295.015 246.155 -294.765 ;
        RECT 249.915 -294.805 251.725 -294.625 ;
        RECT 254.310 -294.670 258.235 -294.240 ;
        RECT 250.950 -294.815 251.725 -294.805 ;
        RECT 251.050 -294.845 251.725 -294.815 ;
        RECT 251.965 -294.730 254.060 -294.690 ;
        RECT 251.965 -294.880 254.115 -294.730 ;
        RECT 247.100 -295.955 247.270 -294.915 ;
        RECT 248.080 -295.955 248.250 -294.915 ;
        RECT 249.060 -295.955 249.230 -294.915 ;
        RECT 251.965 -296.600 252.135 -294.880 ;
        RECT 252.945 -296.600 253.115 -294.880 ;
        RECT 253.810 -295.625 254.115 -294.880 ;
        RECT 255.010 -295.450 255.180 -294.670 ;
        RECT 255.500 -295.450 255.670 -294.910 ;
        RECT 255.990 -295.450 256.160 -294.670 ;
        RECT 256.480 -295.450 256.650 -294.910 ;
        RECT 254.420 -295.625 254.785 -295.595 ;
        RECT 253.810 -295.690 254.785 -295.625 ;
        RECT 253.920 -295.830 254.785 -295.690 ;
        RECT 254.420 -295.895 254.785 -295.830 ;
        RECT 256.970 -295.745 258.830 -295.395 ;
        RECT 255.010 -296.605 255.180 -296.065 ;
        RECT 255.990 -296.605 256.160 -296.065 ;
        RECT 256.970 -296.605 257.140 -295.745 ;
        RECT 255.240 -298.945 256.440 -298.775 ;
        RECT 246.970 -301.280 247.140 -299.560 ;
        RECT 247.950 -301.280 248.120 -299.560 ;
        RECT 250.015 -300.095 250.185 -299.555 ;
        RECT 250.995 -300.095 251.165 -299.555 ;
        RECT 249.425 -300.330 249.790 -300.265 ;
        RECT 248.925 -300.470 249.790 -300.330 ;
        RECT 248.815 -300.535 249.790 -300.470 ;
        RECT 248.815 -301.280 249.120 -300.535 ;
        RECT 249.425 -300.565 249.790 -300.535 ;
        RECT 251.975 -300.415 252.145 -299.555 ;
        RECT 246.970 -301.430 249.120 -301.280 ;
        RECT 246.970 -301.470 249.065 -301.430 ;
        RECT 250.015 -301.490 250.185 -300.710 ;
        RECT 250.505 -301.250 250.675 -300.710 ;
        RECT 250.995 -301.490 251.165 -300.710 ;
        RECT 251.485 -301.250 251.655 -300.710 ;
        RECT 251.975 -300.765 253.365 -300.415 ;
        RECT 245.190 -301.835 246.325 -301.825 ;
        RECT 248.380 -301.835 248.750 -301.705 ;
        RECT 241.480 -302.120 242.905 -301.905 ;
        RECT 245.190 -302.025 248.750 -301.835 ;
        RECT 249.315 -301.920 252.390 -301.490 ;
        RECT 246.320 -302.030 248.750 -302.025 ;
        RECT 246.320 -302.035 246.675 -302.030 ;
        RECT 248.380 -302.060 248.750 -302.030 ;
        RECT 240.085 -302.635 240.610 -302.275 ;
        RECT 242.690 -303.150 242.905 -302.120 ;
        RECT 230.250 -303.890 232.500 -303.800 ;
        RECT 228.040 -304.105 232.500 -303.890 ;
        RECT 228.040 -304.195 230.285 -304.105 ;
        RECT 232.195 -305.580 232.500 -304.105 ;
        RECT 235.865 -304.990 236.035 -303.520 ;
        RECT 236.325 -303.600 236.550 -303.250 ;
        RECT 238.285 -303.350 242.905 -303.150 ;
        RECT 238.525 -303.365 242.905 -303.350 ;
        RECT 235.830 -305.580 236.065 -304.990 ;
        RECT 236.355 -305.060 236.525 -303.600 ;
        RECT 236.845 -304.985 237.015 -303.520 ;
        RECT 238.055 -304.935 238.225 -303.520 ;
        RECT 238.525 -303.565 238.745 -303.365 ;
        RECT 236.810 -305.580 237.045 -304.985 ;
        RECT 238.020 -305.580 238.255 -304.935 ;
        RECT 238.545 -305.060 238.715 -303.565 ;
        RECT 246.480 -303.785 246.650 -302.245 ;
        RECT 246.970 -303.785 247.140 -302.245 ;
        RECT 247.460 -303.785 247.630 -302.245 ;
        RECT 247.950 -303.785 248.120 -302.245 ;
        RECT 248.440 -303.785 248.610 -302.245 ;
        RECT 246.965 -304.045 247.140 -303.785 ;
        RECT 250.535 -303.955 250.840 -301.920 ;
        RECT 252.985 -302.740 253.335 -300.765 ;
        RECT 254.205 -302.035 254.375 -299.115 ;
        RECT 255.240 -299.155 255.450 -298.945 ;
        RECT 254.185 -302.330 254.395 -302.035 ;
        RECT 255.260 -302.065 255.430 -299.155 ;
        RECT 255.750 -302.055 255.920 -299.115 ;
        RECT 256.230 -299.165 256.440 -298.945 ;
        RECT 255.245 -302.330 255.455 -302.065 ;
        RECT 254.185 -302.510 255.455 -302.330 ;
        RECT 255.730 -302.325 255.940 -302.055 ;
        RECT 256.240 -302.155 256.410 -299.165 ;
        RECT 257.300 -302.085 257.470 -299.115 ;
        RECT 255.730 -302.520 256.435 -302.325 ;
        RECT 256.220 -302.580 256.435 -302.520 ;
        RECT 255.010 -302.740 255.785 -302.690 ;
        RECT 252.985 -302.920 255.785 -302.740 ;
        RECT 252.985 -302.930 253.335 -302.920 ;
        RECT 255.010 -302.965 255.785 -302.920 ;
        RECT 256.220 -302.855 257.125 -302.580 ;
        RECT 256.220 -303.205 256.435 -302.855 ;
        RECT 253.660 -303.275 254.435 -303.230 ;
        RECT 253.475 -303.445 254.435 -303.275 ;
        RECT 253.660 -303.505 254.435 -303.445 ;
        RECT 254.665 -303.405 256.435 -303.205 ;
        RECT 257.295 -303.305 257.510 -302.085 ;
        RECT 258.480 -302.430 258.830 -295.745 ;
        RECT 258.425 -302.790 258.950 -302.430 ;
        RECT 261.075 -303.305 262.145 -302.730 ;
        RECT 248.590 -304.045 250.840 -303.955 ;
        RECT 246.380 -304.260 250.840 -304.045 ;
        RECT 246.380 -304.350 248.625 -304.260 ;
        RECT 232.195 -306.145 239.580 -305.580 ;
        RECT 250.535 -305.735 250.840 -304.260 ;
        RECT 254.205 -305.145 254.375 -303.675 ;
        RECT 254.665 -303.755 254.890 -303.405 ;
        RECT 256.625 -303.505 262.635 -303.305 ;
        RECT 256.865 -303.520 262.635 -303.505 ;
        RECT 254.170 -305.735 254.405 -305.145 ;
        RECT 254.695 -305.215 254.865 -303.755 ;
        RECT 255.185 -305.140 255.355 -303.675 ;
        RECT 256.395 -305.090 256.565 -303.675 ;
        RECT 256.865 -303.720 257.085 -303.520 ;
        RECT 255.150 -305.735 255.385 -305.140 ;
        RECT 256.360 -305.735 256.595 -305.090 ;
        RECT 256.885 -305.215 257.055 -303.720 ;
        RECT 261.075 -303.830 262.145 -303.520 ;
        RECT 250.535 -306.300 257.920 -305.735 ;
        RECT 269.380 -309.200 270.185 -289.595 ;
        RECT 272.935 -290.075 273.315 -289.595 ;
        RECT 299.360 -290.045 299.550 -285.570 ;
        RECT 316.705 -288.925 317.085 -284.105 ;
        RECT 317.780 -284.110 320.210 -284.105 ;
        RECT 317.780 -284.115 318.135 -284.110 ;
        RECT 319.840 -284.140 320.210 -284.110 ;
        RECT 317.940 -285.865 318.110 -284.325 ;
        RECT 318.430 -285.865 318.600 -284.325 ;
        RECT 318.920 -285.865 319.090 -284.325 ;
        RECT 319.410 -285.865 319.580 -284.325 ;
        RECT 319.900 -285.865 320.070 -284.325 ;
        RECT 318.425 -286.125 318.600 -285.865 ;
        RECT 321.995 -286.035 322.300 -284.000 ;
        RECT 324.445 -284.820 324.795 -282.845 ;
        RECT 325.665 -284.115 325.835 -281.195 ;
        RECT 326.700 -281.235 326.910 -281.025 ;
        RECT 325.645 -284.410 325.855 -284.115 ;
        RECT 326.720 -284.145 326.890 -281.235 ;
        RECT 327.210 -284.135 327.380 -281.195 ;
        RECT 327.690 -281.245 327.900 -281.025 ;
        RECT 326.705 -284.410 326.915 -284.145 ;
        RECT 325.645 -284.590 326.915 -284.410 ;
        RECT 327.190 -284.405 327.400 -284.135 ;
        RECT 327.700 -284.235 327.870 -281.245 ;
        RECT 328.760 -284.165 328.930 -281.195 ;
        RECT 327.190 -284.600 327.895 -284.405 ;
        RECT 327.680 -284.660 327.895 -284.600 ;
        RECT 326.470 -284.820 327.245 -284.770 ;
        RECT 324.445 -285.000 327.245 -284.820 ;
        RECT 324.445 -285.010 324.795 -285.000 ;
        RECT 326.470 -285.045 327.245 -285.000 ;
        RECT 327.680 -284.935 328.585 -284.660 ;
        RECT 327.680 -285.285 327.895 -284.935 ;
        RECT 325.120 -285.355 325.895 -285.310 ;
        RECT 324.935 -285.525 325.895 -285.355 ;
        RECT 325.120 -285.585 325.895 -285.525 ;
        RECT 326.125 -285.485 327.895 -285.285 ;
        RECT 328.755 -285.385 328.970 -284.165 ;
        RECT 329.940 -284.510 330.290 -277.825 ;
        RECT 364.325 -277.950 364.495 -276.910 ;
        RECT 365.305 -277.950 365.475 -276.910 ;
        RECT 366.285 -277.950 366.455 -276.910 ;
        RECT 369.190 -278.595 369.360 -276.875 ;
        RECT 370.170 -278.595 370.340 -276.875 ;
        RECT 371.035 -277.620 371.340 -276.875 ;
        RECT 372.235 -277.445 372.405 -276.665 ;
        RECT 372.725 -277.445 372.895 -276.905 ;
        RECT 373.215 -277.445 373.385 -276.665 ;
        RECT 416.010 -276.685 418.160 -276.535 ;
        RECT 373.705 -277.445 373.875 -276.905 ;
        RECT 371.645 -277.620 372.010 -277.590 ;
        RECT 371.035 -277.685 372.010 -277.620 ;
        RECT 371.145 -277.825 372.010 -277.685 ;
        RECT 371.645 -277.890 372.010 -277.825 ;
        RECT 374.195 -277.740 376.055 -277.390 ;
        RECT 372.235 -278.600 372.405 -278.060 ;
        RECT 373.215 -278.600 373.385 -278.060 ;
        RECT 374.195 -278.600 374.365 -277.740 ;
        RECT 336.520 -280.305 338.125 -280.135 ;
        RECT 335.625 -282.985 335.795 -280.485 ;
        RECT 335.620 -283.215 335.795 -282.985 ;
        RECT 336.520 -283.215 336.720 -280.305 ;
        RECT 336.965 -280.505 337.140 -280.305 ;
        RECT 336.970 -283.025 337.140 -280.505 ;
        RECT 337.460 -282.990 337.630 -280.485 ;
        RECT 337.950 -280.500 338.125 -280.305 ;
        RECT 335.620 -283.415 336.720 -283.215 ;
        RECT 337.445 -283.590 337.635 -282.990 ;
        RECT 337.950 -283.025 338.120 -280.500 ;
        RECT 338.600 -283.405 338.770 -280.485 ;
        RECT 340.230 -283.055 340.400 -280.485 ;
        RECT 341.370 -281.935 341.540 -280.485 ;
        RECT 372.465 -280.940 373.665 -280.770 ;
        RECT 341.365 -282.400 341.550 -281.935 ;
        RECT 341.365 -282.585 342.050 -282.400 ;
        RECT 340.230 -283.225 341.025 -283.055 ;
        RECT 339.345 -283.405 340.035 -283.350 ;
        RECT 335.625 -283.780 337.635 -283.590 ;
        RECT 337.970 -283.575 340.035 -283.405 ;
        RECT 334.440 -283.835 335.130 -283.785 ;
        RECT 332.490 -284.005 335.130 -283.835 ;
        RECT 329.885 -284.870 330.410 -284.510 ;
        RECT 332.490 -285.385 332.705 -284.005 ;
        RECT 334.440 -284.055 335.130 -284.005 ;
        RECT 334.720 -284.510 335.410 -284.465 ;
        RECT 333.670 -284.680 335.410 -284.510 ;
        RECT 333.670 -285.315 334.030 -284.680 ;
        RECT 334.720 -284.735 335.410 -284.680 ;
        RECT 333.670 -285.360 334.090 -285.315 ;
        RECT 320.050 -286.125 322.300 -286.035 ;
        RECT 317.840 -286.340 322.300 -286.125 ;
        RECT 317.840 -286.430 320.085 -286.340 ;
        RECT 321.995 -287.815 322.300 -286.340 ;
        RECT 325.665 -287.225 325.835 -285.755 ;
        RECT 326.125 -285.835 326.350 -285.485 ;
        RECT 328.085 -285.585 332.705 -285.385 ;
        RECT 328.325 -285.600 332.705 -285.585 ;
        RECT 325.630 -287.815 325.865 -287.225 ;
        RECT 326.155 -287.295 326.325 -285.835 ;
        RECT 326.645 -287.220 326.815 -285.755 ;
        RECT 327.855 -287.170 328.025 -285.755 ;
        RECT 328.325 -285.800 328.545 -285.600 ;
        RECT 333.695 -285.710 334.090 -285.360 ;
        RECT 326.610 -287.815 326.845 -287.220 ;
        RECT 327.820 -287.815 328.055 -287.170 ;
        RECT 328.345 -287.295 328.515 -285.800 ;
        RECT 335.135 -286.920 335.305 -285.465 ;
        RECT 335.125 -287.475 335.310 -286.920 ;
        RECT 335.625 -287.005 335.795 -283.780 ;
        RECT 336.770 -284.130 336.960 -283.780 ;
        RECT 337.970 -283.970 338.140 -283.575 ;
        RECT 339.345 -283.620 340.035 -283.575 ;
        RECT 336.720 -284.820 336.990 -284.130 ;
        RECT 337.485 -284.140 338.140 -283.970 ;
        RECT 338.470 -284.055 339.160 -283.785 ;
        RECT 340.395 -284.130 340.665 -283.440 ;
        RECT 340.855 -283.445 341.025 -283.225 ;
        RECT 340.855 -283.715 341.685 -283.445 ;
        RECT 337.485 -287.005 337.655 -284.140 ;
        RECT 340.855 -284.290 341.025 -283.715 ;
        RECT 341.285 -284.290 341.555 -284.205 ;
        RECT 337.975 -284.485 338.770 -284.310 ;
        RECT 340.855 -284.315 341.555 -284.290 ;
        RECT 340.715 -284.460 341.555 -284.315 ;
        RECT 337.975 -287.005 338.145 -284.485 ;
        RECT 338.600 -287.005 338.770 -284.485 ;
        RECT 339.090 -286.920 339.260 -284.465 ;
        RECT 339.740 -286.915 339.910 -284.465 ;
        RECT 332.440 -287.495 335.495 -287.475 ;
        RECT 339.085 -287.495 339.270 -286.920 ;
        RECT 339.725 -287.495 339.910 -286.915 ;
        RECT 340.230 -287.005 340.400 -284.465 ;
        RECT 340.715 -284.485 341.025 -284.460 ;
        RECT 340.720 -287.005 340.890 -284.485 ;
        RECT 341.285 -284.500 341.555 -284.460 ;
        RECT 341.860 -285.050 342.050 -282.585 ;
        RECT 364.195 -283.275 364.365 -281.555 ;
        RECT 365.175 -283.275 365.345 -281.555 ;
        RECT 367.240 -282.090 367.410 -281.550 ;
        RECT 368.220 -282.090 368.390 -281.550 ;
        RECT 366.650 -282.325 367.015 -282.260 ;
        RECT 366.150 -282.465 367.015 -282.325 ;
        RECT 366.040 -282.530 367.015 -282.465 ;
        RECT 366.040 -283.275 366.345 -282.530 ;
        RECT 366.650 -282.560 367.015 -282.530 ;
        RECT 369.200 -282.410 369.370 -281.550 ;
        RECT 364.195 -283.425 366.345 -283.275 ;
        RECT 364.195 -283.465 366.290 -283.425 ;
        RECT 367.240 -283.485 367.410 -282.705 ;
        RECT 367.730 -283.245 367.900 -282.705 ;
        RECT 368.220 -283.485 368.390 -282.705 ;
        RECT 368.710 -283.245 368.880 -282.705 ;
        RECT 369.200 -282.760 370.590 -282.410 ;
        RECT 362.415 -283.830 363.550 -283.820 ;
        RECT 365.605 -283.830 365.975 -283.700 ;
        RECT 362.415 -284.020 365.975 -283.830 ;
        RECT 366.540 -283.915 369.615 -283.485 ;
        RECT 341.860 -285.240 343.320 -285.050 ;
        RECT 341.370 -286.910 341.540 -285.465 ;
        RECT 341.860 -285.490 342.050 -285.240 ;
        RECT 341.360 -287.495 341.545 -286.910 ;
        RECT 341.860 -287.005 342.030 -285.490 ;
        RECT 332.440 -287.815 342.110 -287.495 ;
        RECT 321.995 -288.040 342.110 -287.815 ;
        RECT 321.995 -288.380 333.005 -288.040 ;
        RECT 334.745 -288.300 342.110 -288.040 ;
        RECT 272.935 -290.455 289.485 -290.075 ;
        RECT 272.935 -291.365 273.315 -290.455 ;
        RECT 272.935 -291.745 273.645 -291.365 ;
        RECT 273.265 -293.690 273.645 -291.745 ;
        RECT 278.310 -291.575 281.635 -291.435 ;
        RECT 278.310 -291.865 283.485 -291.575 ;
        RECT 287.355 -291.860 287.815 -291.435 ;
        RECT 278.310 -292.270 278.740 -291.865 ;
        RECT 279.610 -292.050 279.785 -291.865 ;
        RECT 281.235 -291.880 283.485 -291.865 ;
        RECT 274.050 -292.700 278.740 -292.270 ;
        RECT 273.265 -294.150 273.940 -293.690 ;
        RECT 274.750 -293.980 274.920 -292.700 ;
        RECT 275.240 -293.980 275.410 -292.940 ;
        RECT 275.730 -293.980 275.900 -292.700 ;
        RECT 276.220 -293.810 276.390 -292.940 ;
        RECT 279.125 -293.590 279.295 -292.050 ;
        RECT 279.615 -293.590 279.785 -292.050 ;
        RECT 280.105 -293.590 280.275 -292.050 ;
        RECT 280.595 -293.590 280.765 -292.050 ;
        RECT 281.085 -293.590 281.255 -292.050 ;
        RECT 278.965 -293.805 279.320 -293.800 ;
        RECT 281.025 -293.805 281.395 -293.775 ;
        RECT 278.965 -293.810 281.395 -293.805 ;
        RECT 276.220 -293.980 281.395 -293.810 ;
        RECT 283.180 -293.915 283.485 -291.880 ;
        RECT 276.225 -294.000 281.395 -293.980 ;
        RECT 276.225 -294.010 278.970 -294.000 ;
        RECT 274.160 -294.150 274.525 -294.120 ;
        RECT 281.025 -294.130 281.395 -294.000 ;
        RECT 273.265 -294.235 274.525 -294.150 ;
        RECT 273.290 -294.355 274.525 -294.235 ;
        RECT 278.700 -294.290 279.375 -294.250 ;
        RECT 278.600 -294.300 279.375 -294.290 ;
        RECT 273.290 -294.440 273.940 -294.355 ;
        RECT 274.160 -294.420 274.525 -294.355 ;
        RECT 277.565 -294.480 279.375 -294.300 ;
        RECT 281.960 -294.345 285.885 -293.915 ;
        RECT 278.600 -294.490 279.375 -294.480 ;
        RECT 278.700 -294.520 279.375 -294.490 ;
        RECT 279.615 -294.405 281.710 -294.365 ;
        RECT 279.615 -294.555 281.765 -294.405 ;
        RECT 274.750 -295.630 274.920 -294.590 ;
        RECT 275.730 -295.630 275.900 -294.590 ;
        RECT 276.710 -295.630 276.880 -294.590 ;
        RECT 279.615 -296.275 279.785 -294.555 ;
        RECT 280.595 -296.275 280.765 -294.555 ;
        RECT 281.460 -295.300 281.765 -294.555 ;
        RECT 282.660 -295.125 282.830 -294.345 ;
        RECT 283.150 -295.125 283.320 -294.585 ;
        RECT 283.640 -295.125 283.810 -294.345 ;
        RECT 284.130 -295.125 284.300 -294.585 ;
        RECT 282.070 -295.300 282.435 -295.270 ;
        RECT 281.460 -295.365 282.435 -295.300 ;
        RECT 281.570 -295.505 282.435 -295.365 ;
        RECT 282.070 -295.570 282.435 -295.505 ;
        RECT 284.620 -295.420 286.480 -295.070 ;
        RECT 282.660 -296.280 282.830 -295.740 ;
        RECT 283.640 -296.280 283.810 -295.740 ;
        RECT 284.620 -296.280 284.790 -295.420 ;
        RECT 282.890 -298.620 284.090 -298.450 ;
        RECT 274.620 -300.955 274.790 -299.235 ;
        RECT 275.600 -300.955 275.770 -299.235 ;
        RECT 277.665 -299.770 277.835 -299.230 ;
        RECT 278.645 -299.770 278.815 -299.230 ;
        RECT 277.075 -300.005 277.440 -299.940 ;
        RECT 276.575 -300.145 277.440 -300.005 ;
        RECT 276.465 -300.210 277.440 -300.145 ;
        RECT 276.465 -300.955 276.770 -300.210 ;
        RECT 277.075 -300.240 277.440 -300.210 ;
        RECT 279.625 -300.090 279.795 -299.230 ;
        RECT 274.620 -301.105 276.770 -300.955 ;
        RECT 274.620 -301.145 276.715 -301.105 ;
        RECT 277.665 -301.165 277.835 -300.385 ;
        RECT 278.155 -300.925 278.325 -300.385 ;
        RECT 278.645 -301.165 278.815 -300.385 ;
        RECT 279.135 -300.925 279.305 -300.385 ;
        RECT 279.625 -300.440 281.015 -300.090 ;
        RECT 272.840 -301.510 273.975 -301.500 ;
        RECT 276.030 -301.510 276.400 -301.380 ;
        RECT 272.840 -301.700 276.400 -301.510 ;
        RECT 276.965 -301.595 280.040 -301.165 ;
        RECT 273.970 -301.705 276.400 -301.700 ;
        RECT 273.970 -301.710 274.325 -301.705 ;
        RECT 276.030 -301.735 276.400 -301.705 ;
        RECT 274.130 -303.460 274.300 -301.920 ;
        RECT 274.620 -303.460 274.790 -301.920 ;
        RECT 275.110 -303.460 275.280 -301.920 ;
        RECT 275.600 -303.460 275.770 -301.920 ;
        RECT 276.090 -303.460 276.260 -301.920 ;
        RECT 274.615 -303.720 274.790 -303.460 ;
        RECT 278.185 -303.630 278.490 -301.595 ;
        RECT 280.635 -302.415 280.985 -300.440 ;
        RECT 281.855 -301.710 282.025 -298.790 ;
        RECT 282.890 -298.830 283.100 -298.620 ;
        RECT 281.835 -302.005 282.045 -301.710 ;
        RECT 282.910 -301.740 283.080 -298.830 ;
        RECT 283.400 -301.730 283.570 -298.790 ;
        RECT 283.880 -298.840 284.090 -298.620 ;
        RECT 282.895 -302.005 283.105 -301.740 ;
        RECT 281.835 -302.185 283.105 -302.005 ;
        RECT 283.380 -302.000 283.590 -301.730 ;
        RECT 283.890 -301.830 284.060 -298.840 ;
        RECT 284.950 -301.760 285.120 -298.790 ;
        RECT 283.380 -302.195 284.085 -302.000 ;
        RECT 283.870 -302.255 284.085 -302.195 ;
        RECT 282.660 -302.415 283.435 -302.365 ;
        RECT 280.635 -302.595 283.435 -302.415 ;
        RECT 280.635 -302.605 280.985 -302.595 ;
        RECT 282.660 -302.640 283.435 -302.595 ;
        RECT 283.870 -302.530 284.775 -302.255 ;
        RECT 283.870 -302.880 284.085 -302.530 ;
        RECT 281.310 -302.950 282.085 -302.905 ;
        RECT 281.125 -303.120 282.085 -302.950 ;
        RECT 281.310 -303.180 282.085 -303.120 ;
        RECT 282.315 -303.080 284.085 -302.880 ;
        RECT 284.945 -302.980 285.160 -301.760 ;
        RECT 286.130 -302.105 286.480 -295.420 ;
        RECT 287.470 -301.735 287.685 -291.860 ;
        RECT 289.105 -293.975 289.485 -290.455 ;
        RECT 290.615 -290.235 299.550 -290.045 ;
        RECT 313.140 -289.745 317.085 -288.925 ;
        RECT 343.130 -289.715 343.320 -285.240 ;
        RECT 362.470 -289.130 362.850 -284.020 ;
        RECT 363.545 -284.025 365.975 -284.020 ;
        RECT 363.545 -284.030 363.900 -284.025 ;
        RECT 365.605 -284.055 365.975 -284.025 ;
        RECT 363.705 -285.780 363.875 -284.240 ;
        RECT 364.195 -285.780 364.365 -284.240 ;
        RECT 364.685 -285.780 364.855 -284.240 ;
        RECT 365.175 -285.780 365.345 -284.240 ;
        RECT 365.665 -285.780 365.835 -284.240 ;
        RECT 364.190 -286.040 364.365 -285.780 ;
        RECT 367.760 -285.950 368.065 -283.915 ;
        RECT 370.210 -284.735 370.560 -282.760 ;
        RECT 371.430 -284.030 371.600 -281.110 ;
        RECT 372.465 -281.150 372.675 -280.940 ;
        RECT 371.410 -284.325 371.620 -284.030 ;
        RECT 372.485 -284.060 372.655 -281.150 ;
        RECT 372.975 -284.050 373.145 -281.110 ;
        RECT 373.455 -281.160 373.665 -280.940 ;
        RECT 372.470 -284.325 372.680 -284.060 ;
        RECT 371.410 -284.505 372.680 -284.325 ;
        RECT 372.955 -284.320 373.165 -284.050 ;
        RECT 373.465 -284.150 373.635 -281.160 ;
        RECT 374.525 -284.080 374.695 -281.110 ;
        RECT 372.955 -284.515 373.660 -284.320 ;
        RECT 373.445 -284.575 373.660 -284.515 ;
        RECT 372.235 -284.735 373.010 -284.685 ;
        RECT 370.210 -284.915 373.010 -284.735 ;
        RECT 370.210 -284.925 370.560 -284.915 ;
        RECT 372.235 -284.960 373.010 -284.915 ;
        RECT 373.445 -284.850 374.350 -284.575 ;
        RECT 373.445 -285.200 373.660 -284.850 ;
        RECT 370.885 -285.270 371.660 -285.225 ;
        RECT 370.700 -285.440 371.660 -285.270 ;
        RECT 370.885 -285.500 371.660 -285.440 ;
        RECT 371.890 -285.400 373.660 -285.200 ;
        RECT 374.520 -285.300 374.735 -284.080 ;
        RECT 375.705 -284.425 376.055 -277.740 ;
        RECT 411.145 -277.760 411.315 -276.720 ;
        RECT 412.125 -277.760 412.295 -276.720 ;
        RECT 413.105 -277.760 413.275 -276.720 ;
        RECT 416.010 -278.405 416.180 -276.685 ;
        RECT 416.990 -278.405 417.160 -276.685 ;
        RECT 417.855 -277.430 418.160 -276.685 ;
        RECT 419.055 -277.255 419.225 -276.475 ;
        RECT 419.545 -277.255 419.715 -276.715 ;
        RECT 420.035 -277.255 420.205 -276.475 ;
        RECT 420.525 -277.255 420.695 -276.715 ;
        RECT 418.465 -277.430 418.830 -277.400 ;
        RECT 417.855 -277.495 418.830 -277.430 ;
        RECT 417.965 -277.635 418.830 -277.495 ;
        RECT 418.465 -277.700 418.830 -277.635 ;
        RECT 421.015 -277.550 422.875 -277.200 ;
        RECT 419.055 -278.410 419.225 -277.870 ;
        RECT 420.035 -278.410 420.205 -277.870 ;
        RECT 421.015 -278.410 421.185 -277.550 ;
        RECT 382.285 -280.220 383.890 -280.050 ;
        RECT 381.390 -282.900 381.560 -280.400 ;
        RECT 381.385 -283.130 381.560 -282.900 ;
        RECT 382.285 -283.130 382.485 -280.220 ;
        RECT 382.730 -280.420 382.905 -280.220 ;
        RECT 382.735 -282.940 382.905 -280.420 ;
        RECT 383.225 -282.905 383.395 -280.400 ;
        RECT 383.715 -280.415 383.890 -280.220 ;
        RECT 381.385 -283.330 382.485 -283.130 ;
        RECT 383.210 -283.505 383.400 -282.905 ;
        RECT 383.715 -282.940 383.885 -280.415 ;
        RECT 384.365 -283.320 384.535 -280.400 ;
        RECT 385.995 -282.970 386.165 -280.400 ;
        RECT 387.135 -281.850 387.305 -280.400 ;
        RECT 419.285 -280.750 420.485 -280.580 ;
        RECT 387.130 -282.315 387.315 -281.850 ;
        RECT 387.130 -282.500 387.815 -282.315 ;
        RECT 385.995 -283.140 386.790 -282.970 ;
        RECT 385.110 -283.320 385.800 -283.265 ;
        RECT 381.390 -283.695 383.400 -283.505 ;
        RECT 383.735 -283.490 385.800 -283.320 ;
        RECT 380.205 -283.750 380.895 -283.700 ;
        RECT 378.255 -283.920 380.895 -283.750 ;
        RECT 375.650 -284.785 376.175 -284.425 ;
        RECT 378.255 -285.300 378.470 -283.920 ;
        RECT 380.205 -283.970 380.895 -283.920 ;
        RECT 380.485 -284.425 381.175 -284.380 ;
        RECT 379.435 -284.595 381.175 -284.425 ;
        RECT 379.435 -285.230 379.795 -284.595 ;
        RECT 380.485 -284.650 381.175 -284.595 ;
        RECT 379.435 -285.275 379.855 -285.230 ;
        RECT 365.815 -286.040 368.065 -285.950 ;
        RECT 363.605 -286.255 368.065 -286.040 ;
        RECT 363.605 -286.345 365.850 -286.255 ;
        RECT 367.760 -287.730 368.065 -286.255 ;
        RECT 371.430 -287.140 371.600 -285.670 ;
        RECT 371.890 -285.750 372.115 -285.400 ;
        RECT 373.850 -285.500 378.470 -285.300 ;
        RECT 374.090 -285.515 378.470 -285.500 ;
        RECT 371.395 -287.730 371.630 -287.140 ;
        RECT 371.920 -287.210 372.090 -285.750 ;
        RECT 372.410 -287.135 372.580 -285.670 ;
        RECT 373.620 -287.085 373.790 -285.670 ;
        RECT 374.090 -285.715 374.310 -285.515 ;
        RECT 379.460 -285.625 379.855 -285.275 ;
        RECT 372.375 -287.730 372.610 -287.135 ;
        RECT 373.585 -287.730 373.820 -287.085 ;
        RECT 374.110 -287.210 374.280 -285.715 ;
        RECT 380.900 -286.835 381.070 -285.380 ;
        RECT 380.890 -287.390 381.075 -286.835 ;
        RECT 381.390 -286.920 381.560 -283.695 ;
        RECT 382.535 -284.045 382.725 -283.695 ;
        RECT 383.735 -283.885 383.905 -283.490 ;
        RECT 385.110 -283.535 385.800 -283.490 ;
        RECT 382.485 -284.735 382.755 -284.045 ;
        RECT 383.250 -284.055 383.905 -283.885 ;
        RECT 384.235 -283.970 384.925 -283.700 ;
        RECT 386.160 -284.045 386.430 -283.355 ;
        RECT 386.620 -283.360 386.790 -283.140 ;
        RECT 386.620 -283.630 387.450 -283.360 ;
        RECT 383.250 -286.920 383.420 -284.055 ;
        RECT 386.620 -284.205 386.790 -283.630 ;
        RECT 387.050 -284.205 387.320 -284.120 ;
        RECT 383.740 -284.400 384.535 -284.225 ;
        RECT 386.620 -284.230 387.320 -284.205 ;
        RECT 386.480 -284.375 387.320 -284.230 ;
        RECT 383.740 -286.920 383.910 -284.400 ;
        RECT 384.365 -286.920 384.535 -284.400 ;
        RECT 384.855 -286.835 385.025 -284.380 ;
        RECT 385.505 -286.830 385.675 -284.380 ;
        RECT 378.205 -287.410 381.260 -287.390 ;
        RECT 384.850 -287.410 385.035 -286.835 ;
        RECT 385.490 -287.410 385.675 -286.830 ;
        RECT 385.995 -286.920 386.165 -284.380 ;
        RECT 386.480 -284.400 386.790 -284.375 ;
        RECT 386.485 -286.920 386.655 -284.400 ;
        RECT 387.050 -284.415 387.320 -284.375 ;
        RECT 387.625 -284.965 387.815 -282.500 ;
        RECT 411.015 -283.085 411.185 -281.365 ;
        RECT 411.995 -283.085 412.165 -281.365 ;
        RECT 414.060 -281.900 414.230 -281.360 ;
        RECT 415.040 -281.900 415.210 -281.360 ;
        RECT 413.470 -282.135 413.835 -282.070 ;
        RECT 412.970 -282.275 413.835 -282.135 ;
        RECT 412.860 -282.340 413.835 -282.275 ;
        RECT 412.860 -283.085 413.165 -282.340 ;
        RECT 413.470 -282.370 413.835 -282.340 ;
        RECT 416.020 -282.220 416.190 -281.360 ;
        RECT 411.015 -283.235 413.165 -283.085 ;
        RECT 411.015 -283.275 413.110 -283.235 ;
        RECT 414.060 -283.295 414.230 -282.515 ;
        RECT 414.550 -283.055 414.720 -282.515 ;
        RECT 415.040 -283.295 415.210 -282.515 ;
        RECT 415.530 -283.055 415.700 -282.515 ;
        RECT 416.020 -282.570 417.410 -282.220 ;
        RECT 409.235 -283.640 410.370 -283.630 ;
        RECT 412.425 -283.640 412.795 -283.510 ;
        RECT 409.235 -283.830 412.795 -283.640 ;
        RECT 413.360 -283.725 416.435 -283.295 ;
        RECT 387.625 -285.155 389.085 -284.965 ;
        RECT 387.135 -286.825 387.305 -285.380 ;
        RECT 387.625 -285.405 387.815 -285.155 ;
        RECT 387.125 -287.410 387.310 -286.825 ;
        RECT 387.625 -286.920 387.795 -285.405 ;
        RECT 378.205 -287.730 387.875 -287.410 ;
        RECT 367.760 -287.955 387.875 -287.730 ;
        RECT 367.760 -288.295 378.770 -287.955 ;
        RECT 380.510 -288.215 387.875 -287.955 ;
        RECT 313.140 -290.010 333.255 -289.745 ;
        RECT 290.615 -292.125 290.805 -290.235 ;
        RECT 296.650 -291.730 299.975 -291.590 ;
        RECT 296.650 -292.020 301.825 -291.730 ;
        RECT 290.500 -292.395 290.865 -292.125 ;
        RECT 296.650 -292.425 297.080 -292.020 ;
        RECT 297.950 -292.205 298.125 -292.020 ;
        RECT 299.575 -292.035 301.825 -292.020 ;
        RECT 292.390 -292.855 297.080 -292.425 ;
        RECT 291.630 -293.975 292.280 -293.845 ;
        RECT 289.105 -294.305 292.280 -293.975 ;
        RECT 293.090 -294.135 293.260 -292.855 ;
        RECT 293.580 -294.135 293.750 -293.095 ;
        RECT 294.070 -294.135 294.240 -292.855 ;
        RECT 294.560 -293.965 294.730 -293.095 ;
        RECT 297.465 -293.745 297.635 -292.205 ;
        RECT 297.955 -293.745 298.125 -292.205 ;
        RECT 298.445 -293.745 298.615 -292.205 ;
        RECT 298.935 -293.745 299.105 -292.205 ;
        RECT 299.425 -293.745 299.595 -292.205 ;
        RECT 297.305 -293.960 297.660 -293.955 ;
        RECT 299.365 -293.960 299.735 -293.930 ;
        RECT 297.305 -293.965 299.735 -293.960 ;
        RECT 294.560 -294.135 299.735 -293.965 ;
        RECT 301.520 -294.070 301.825 -292.035 ;
        RECT 294.565 -294.155 299.735 -294.135 ;
        RECT 294.565 -294.165 297.310 -294.155 ;
        RECT 292.500 -294.305 292.865 -294.275 ;
        RECT 299.365 -294.285 299.735 -294.155 ;
        RECT 289.105 -294.355 292.865 -294.305 ;
        RECT 291.630 -294.510 292.865 -294.355 ;
        RECT 297.040 -294.445 297.715 -294.405 ;
        RECT 296.940 -294.455 297.715 -294.445 ;
        RECT 291.630 -294.595 292.280 -294.510 ;
        RECT 292.500 -294.575 292.865 -294.510 ;
        RECT 291.765 -294.845 292.145 -294.595 ;
        RECT 295.905 -294.635 297.715 -294.455 ;
        RECT 300.300 -294.500 304.225 -294.070 ;
        RECT 296.940 -294.645 297.715 -294.635 ;
        RECT 297.040 -294.675 297.715 -294.645 ;
        RECT 297.955 -294.560 300.050 -294.520 ;
        RECT 297.955 -294.710 300.105 -294.560 ;
        RECT 293.090 -295.785 293.260 -294.745 ;
        RECT 294.070 -295.785 294.240 -294.745 ;
        RECT 295.050 -295.785 295.220 -294.745 ;
        RECT 297.955 -296.430 298.125 -294.710 ;
        RECT 298.935 -296.430 299.105 -294.710 ;
        RECT 299.800 -295.455 300.105 -294.710 ;
        RECT 301.000 -295.280 301.170 -294.500 ;
        RECT 301.490 -295.280 301.660 -294.740 ;
        RECT 301.980 -295.280 302.150 -294.500 ;
        RECT 302.470 -295.280 302.640 -294.740 ;
        RECT 300.410 -295.455 300.775 -295.425 ;
        RECT 299.800 -295.520 300.775 -295.455 ;
        RECT 299.910 -295.660 300.775 -295.520 ;
        RECT 300.410 -295.725 300.775 -295.660 ;
        RECT 302.960 -295.575 304.820 -295.225 ;
        RECT 301.000 -296.435 301.170 -295.895 ;
        RECT 301.980 -296.435 302.150 -295.895 ;
        RECT 302.960 -296.435 303.130 -295.575 ;
        RECT 301.230 -298.775 302.430 -298.605 ;
        RECT 292.960 -301.110 293.130 -299.390 ;
        RECT 293.940 -301.110 294.110 -299.390 ;
        RECT 296.005 -299.925 296.175 -299.385 ;
        RECT 296.985 -299.925 297.155 -299.385 ;
        RECT 295.415 -300.160 295.780 -300.095 ;
        RECT 294.915 -300.300 295.780 -300.160 ;
        RECT 294.805 -300.365 295.780 -300.300 ;
        RECT 294.805 -301.110 295.110 -300.365 ;
        RECT 295.415 -300.395 295.780 -300.365 ;
        RECT 297.965 -300.245 298.135 -299.385 ;
        RECT 292.960 -301.260 295.110 -301.110 ;
        RECT 292.960 -301.300 295.055 -301.260 ;
        RECT 296.005 -301.320 296.175 -300.540 ;
        RECT 296.495 -301.080 296.665 -300.540 ;
        RECT 296.985 -301.320 297.155 -300.540 ;
        RECT 297.475 -301.080 297.645 -300.540 ;
        RECT 297.965 -300.595 299.355 -300.245 ;
        RECT 291.180 -301.665 292.315 -301.655 ;
        RECT 294.370 -301.665 294.740 -301.535 ;
        RECT 287.470 -301.950 288.895 -301.735 ;
        RECT 291.180 -301.855 294.740 -301.665 ;
        RECT 295.305 -301.750 298.380 -301.320 ;
        RECT 292.310 -301.860 294.740 -301.855 ;
        RECT 292.310 -301.865 292.665 -301.860 ;
        RECT 294.370 -301.890 294.740 -301.860 ;
        RECT 286.075 -302.465 286.600 -302.105 ;
        RECT 288.680 -302.980 288.895 -301.950 ;
        RECT 276.240 -303.720 278.490 -303.630 ;
        RECT 274.030 -303.935 278.490 -303.720 ;
        RECT 274.030 -304.025 276.275 -303.935 ;
        RECT 278.185 -305.410 278.490 -303.935 ;
        RECT 281.855 -304.820 282.025 -303.350 ;
        RECT 282.315 -303.430 282.540 -303.080 ;
        RECT 284.275 -303.180 288.895 -302.980 ;
        RECT 284.515 -303.195 288.895 -303.180 ;
        RECT 281.820 -305.410 282.055 -304.820 ;
        RECT 282.345 -304.890 282.515 -303.430 ;
        RECT 282.835 -304.815 283.005 -303.350 ;
        RECT 284.045 -304.765 284.215 -303.350 ;
        RECT 284.515 -303.395 284.735 -303.195 ;
        RECT 282.800 -305.410 283.035 -304.815 ;
        RECT 284.010 -305.410 284.245 -304.765 ;
        RECT 284.535 -304.890 284.705 -303.395 ;
        RECT 292.470 -303.615 292.640 -302.075 ;
        RECT 292.960 -303.615 293.130 -302.075 ;
        RECT 293.450 -303.615 293.620 -302.075 ;
        RECT 293.940 -303.615 294.110 -302.075 ;
        RECT 294.430 -303.615 294.600 -302.075 ;
        RECT 292.955 -303.875 293.130 -303.615 ;
        RECT 296.525 -303.785 296.830 -301.750 ;
        RECT 298.975 -302.570 299.325 -300.595 ;
        RECT 300.195 -301.865 300.365 -298.945 ;
        RECT 301.230 -298.985 301.440 -298.775 ;
        RECT 300.175 -302.160 300.385 -301.865 ;
        RECT 301.250 -301.895 301.420 -298.985 ;
        RECT 301.740 -301.885 301.910 -298.945 ;
        RECT 302.220 -298.995 302.430 -298.775 ;
        RECT 301.235 -302.160 301.445 -301.895 ;
        RECT 300.175 -302.340 301.445 -302.160 ;
        RECT 301.720 -302.155 301.930 -301.885 ;
        RECT 302.230 -301.985 302.400 -298.995 ;
        RECT 303.290 -301.915 303.460 -298.945 ;
        RECT 301.720 -302.350 302.425 -302.155 ;
        RECT 302.210 -302.410 302.425 -302.350 ;
        RECT 301.000 -302.570 301.775 -302.520 ;
        RECT 298.975 -302.750 301.775 -302.570 ;
        RECT 298.975 -302.760 299.325 -302.750 ;
        RECT 301.000 -302.795 301.775 -302.750 ;
        RECT 302.210 -302.685 303.115 -302.410 ;
        RECT 302.210 -303.035 302.425 -302.685 ;
        RECT 299.650 -303.105 300.425 -303.060 ;
        RECT 299.465 -303.275 300.425 -303.105 ;
        RECT 299.650 -303.335 300.425 -303.275 ;
        RECT 300.655 -303.235 302.425 -303.035 ;
        RECT 303.285 -303.135 303.500 -301.915 ;
        RECT 304.470 -302.260 304.820 -295.575 ;
        RECT 304.415 -302.620 304.940 -302.260 ;
        RECT 306.705 -303.135 308.165 -302.290 ;
        RECT 294.580 -303.875 296.830 -303.785 ;
        RECT 292.370 -304.090 296.830 -303.875 ;
        RECT 292.370 -304.180 294.615 -304.090 ;
        RECT 278.185 -305.975 285.570 -305.410 ;
        RECT 296.525 -305.565 296.830 -304.090 ;
        RECT 300.195 -304.975 300.365 -303.505 ;
        RECT 300.655 -303.585 300.880 -303.235 ;
        RECT 302.615 -303.335 308.625 -303.135 ;
        RECT 302.855 -303.350 308.625 -303.335 ;
        RECT 300.160 -305.565 300.395 -304.975 ;
        RECT 300.685 -305.045 300.855 -303.585 ;
        RECT 301.175 -304.970 301.345 -303.505 ;
        RECT 302.385 -304.920 302.555 -303.505 ;
        RECT 302.855 -303.550 303.075 -303.350 ;
        RECT 301.140 -305.565 301.375 -304.970 ;
        RECT 302.350 -305.565 302.585 -304.920 ;
        RECT 302.875 -305.045 303.045 -303.550 ;
        RECT 306.705 -303.785 308.165 -303.350 ;
        RECT 296.525 -306.130 303.910 -305.565 ;
        RECT 269.290 -310.035 270.260 -309.200 ;
        RECT 49.650 -311.510 50.410 -311.240 ;
        RECT 49.650 -311.715 49.920 -311.510 ;
        RECT -91.515 -311.940 -90.825 -311.935 ;
        RECT -117.245 -312.290 -114.550 -312.240 ;
        RECT -107.545 -312.165 -106.755 -312.000 ;
        RECT -33.040 -312.030 -32.225 -311.935 ;
        RECT -92.205 -312.165 -91.520 -312.140 ;
        RECT -107.545 -312.425 -91.520 -312.165 ;
        RECT -107.545 -312.580 -106.755 -312.425 ;
        RECT -92.205 -312.430 -91.520 -312.425 ;
        RECT 214.975 -314.110 216.305 -310.210 ;
        RECT 313.140 -312.860 314.225 -290.010 ;
        RECT 316.705 -290.125 333.255 -290.010 ;
        RECT 316.705 -291.035 317.085 -290.125 ;
        RECT 316.705 -291.415 317.415 -291.035 ;
        RECT 317.035 -293.360 317.415 -291.415 ;
        RECT 322.080 -291.245 325.405 -291.105 ;
        RECT 322.080 -291.535 327.255 -291.245 ;
        RECT 331.125 -291.530 331.585 -291.105 ;
        RECT 322.080 -291.940 322.510 -291.535 ;
        RECT 323.380 -291.720 323.555 -291.535 ;
        RECT 325.005 -291.550 327.255 -291.535 ;
        RECT 317.820 -292.370 322.510 -291.940 ;
        RECT 317.035 -293.820 317.710 -293.360 ;
        RECT 318.520 -293.650 318.690 -292.370 ;
        RECT 319.010 -293.650 319.180 -292.610 ;
        RECT 319.500 -293.650 319.670 -292.370 ;
        RECT 319.990 -293.480 320.160 -292.610 ;
        RECT 322.895 -293.260 323.065 -291.720 ;
        RECT 323.385 -293.260 323.555 -291.720 ;
        RECT 323.875 -293.260 324.045 -291.720 ;
        RECT 324.365 -293.260 324.535 -291.720 ;
        RECT 324.855 -293.260 325.025 -291.720 ;
        RECT 322.735 -293.475 323.090 -293.470 ;
        RECT 324.795 -293.475 325.165 -293.445 ;
        RECT 322.735 -293.480 325.165 -293.475 ;
        RECT 319.990 -293.650 325.165 -293.480 ;
        RECT 326.950 -293.585 327.255 -291.550 ;
        RECT 319.995 -293.670 325.165 -293.650 ;
        RECT 319.995 -293.680 322.740 -293.670 ;
        RECT 317.930 -293.820 318.295 -293.790 ;
        RECT 324.795 -293.800 325.165 -293.670 ;
        RECT 317.035 -293.905 318.295 -293.820 ;
        RECT 317.060 -294.025 318.295 -293.905 ;
        RECT 322.470 -293.960 323.145 -293.920 ;
        RECT 322.370 -293.970 323.145 -293.960 ;
        RECT 317.060 -294.110 317.710 -294.025 ;
        RECT 317.930 -294.090 318.295 -294.025 ;
        RECT 321.335 -294.150 323.145 -293.970 ;
        RECT 325.730 -294.015 329.655 -293.585 ;
        RECT 322.370 -294.160 323.145 -294.150 ;
        RECT 322.470 -294.190 323.145 -294.160 ;
        RECT 323.385 -294.075 325.480 -294.035 ;
        RECT 323.385 -294.225 325.535 -294.075 ;
        RECT 318.520 -295.300 318.690 -294.260 ;
        RECT 319.500 -295.300 319.670 -294.260 ;
        RECT 320.480 -295.300 320.650 -294.260 ;
        RECT 323.385 -295.945 323.555 -294.225 ;
        RECT 324.365 -295.945 324.535 -294.225 ;
        RECT 325.230 -294.970 325.535 -294.225 ;
        RECT 326.430 -294.795 326.600 -294.015 ;
        RECT 326.920 -294.795 327.090 -294.255 ;
        RECT 327.410 -294.795 327.580 -294.015 ;
        RECT 327.900 -294.795 328.070 -294.255 ;
        RECT 325.840 -294.970 326.205 -294.940 ;
        RECT 325.230 -295.035 326.205 -294.970 ;
        RECT 325.340 -295.175 326.205 -295.035 ;
        RECT 325.840 -295.240 326.205 -295.175 ;
        RECT 328.390 -295.090 330.250 -294.740 ;
        RECT 326.430 -295.950 326.600 -295.410 ;
        RECT 327.410 -295.950 327.580 -295.410 ;
        RECT 328.390 -295.950 328.560 -295.090 ;
        RECT 326.660 -298.290 327.860 -298.120 ;
        RECT 318.390 -300.625 318.560 -298.905 ;
        RECT 319.370 -300.625 319.540 -298.905 ;
        RECT 321.435 -299.440 321.605 -298.900 ;
        RECT 322.415 -299.440 322.585 -298.900 ;
        RECT 320.845 -299.675 321.210 -299.610 ;
        RECT 320.345 -299.815 321.210 -299.675 ;
        RECT 320.235 -299.880 321.210 -299.815 ;
        RECT 320.235 -300.625 320.540 -299.880 ;
        RECT 320.845 -299.910 321.210 -299.880 ;
        RECT 323.395 -299.760 323.565 -298.900 ;
        RECT 317.475 -300.690 318.150 -300.660 ;
        RECT 317.375 -300.700 318.150 -300.690 ;
        RECT 314.735 -300.880 318.150 -300.700 ;
        RECT 318.390 -300.775 320.540 -300.625 ;
        RECT 318.390 -300.815 320.485 -300.775 ;
        RECT 321.435 -300.835 321.605 -300.055 ;
        RECT 321.925 -300.595 322.095 -300.055 ;
        RECT 322.415 -300.835 322.585 -300.055 ;
        RECT 322.905 -300.595 323.075 -300.055 ;
        RECT 323.395 -300.110 324.785 -299.760 ;
        RECT 315.650 -306.015 316.330 -300.880 ;
        RECT 317.375 -300.890 318.150 -300.880 ;
        RECT 317.475 -300.930 318.150 -300.890 ;
        RECT 316.610 -301.180 317.745 -301.170 ;
        RECT 319.800 -301.180 320.170 -301.050 ;
        RECT 316.610 -301.370 320.170 -301.180 ;
        RECT 320.735 -301.265 323.810 -300.835 ;
        RECT 317.740 -301.375 320.170 -301.370 ;
        RECT 317.740 -301.380 318.095 -301.375 ;
        RECT 319.800 -301.405 320.170 -301.375 ;
        RECT 317.900 -303.130 318.070 -301.590 ;
        RECT 318.390 -303.130 318.560 -301.590 ;
        RECT 318.880 -303.130 319.050 -301.590 ;
        RECT 319.370 -303.130 319.540 -301.590 ;
        RECT 319.860 -303.130 320.030 -301.590 ;
        RECT 318.385 -303.390 318.560 -303.130 ;
        RECT 321.955 -303.300 322.260 -301.265 ;
        RECT 324.405 -302.085 324.755 -300.110 ;
        RECT 325.625 -301.380 325.795 -298.460 ;
        RECT 326.660 -298.500 326.870 -298.290 ;
        RECT 325.605 -301.675 325.815 -301.380 ;
        RECT 326.680 -301.410 326.850 -298.500 ;
        RECT 327.170 -301.400 327.340 -298.460 ;
        RECT 327.650 -298.510 327.860 -298.290 ;
        RECT 326.665 -301.675 326.875 -301.410 ;
        RECT 325.605 -301.855 326.875 -301.675 ;
        RECT 327.150 -301.670 327.360 -301.400 ;
        RECT 327.660 -301.500 327.830 -298.510 ;
        RECT 328.720 -301.430 328.890 -298.460 ;
        RECT 327.150 -301.865 327.855 -301.670 ;
        RECT 327.640 -301.925 327.855 -301.865 ;
        RECT 326.430 -302.085 327.205 -302.035 ;
        RECT 324.405 -302.265 327.205 -302.085 ;
        RECT 324.405 -302.275 324.755 -302.265 ;
        RECT 326.430 -302.310 327.205 -302.265 ;
        RECT 327.640 -302.200 328.545 -301.925 ;
        RECT 327.640 -302.550 327.855 -302.200 ;
        RECT 325.080 -302.620 325.855 -302.575 ;
        RECT 324.895 -302.790 325.855 -302.620 ;
        RECT 325.080 -302.850 325.855 -302.790 ;
        RECT 326.085 -302.750 327.855 -302.550 ;
        RECT 328.715 -302.650 328.930 -301.430 ;
        RECT 329.900 -301.775 330.250 -295.090 ;
        RECT 331.240 -301.405 331.455 -291.530 ;
        RECT 332.875 -293.645 333.255 -290.125 ;
        RECT 334.385 -289.905 343.320 -289.715 ;
        RECT 359.095 -289.660 362.850 -289.130 ;
        RECT 388.895 -289.630 389.085 -285.155 ;
        RECT 409.290 -288.735 409.670 -283.830 ;
        RECT 410.365 -283.835 412.795 -283.830 ;
        RECT 410.365 -283.840 410.720 -283.835 ;
        RECT 412.425 -283.865 412.795 -283.835 ;
        RECT 410.525 -285.590 410.695 -284.050 ;
        RECT 411.015 -285.590 411.185 -284.050 ;
        RECT 411.505 -285.590 411.675 -284.050 ;
        RECT 411.995 -285.590 412.165 -284.050 ;
        RECT 412.485 -285.590 412.655 -284.050 ;
        RECT 411.010 -285.850 411.185 -285.590 ;
        RECT 414.580 -285.760 414.885 -283.725 ;
        RECT 417.030 -284.545 417.380 -282.570 ;
        RECT 418.250 -283.840 418.420 -280.920 ;
        RECT 419.285 -280.960 419.495 -280.750 ;
        RECT 418.230 -284.135 418.440 -283.840 ;
        RECT 419.305 -283.870 419.475 -280.960 ;
        RECT 419.795 -283.860 419.965 -280.920 ;
        RECT 420.275 -280.970 420.485 -280.750 ;
        RECT 419.290 -284.135 419.500 -283.870 ;
        RECT 418.230 -284.315 419.500 -284.135 ;
        RECT 419.775 -284.130 419.985 -283.860 ;
        RECT 420.285 -283.960 420.455 -280.970 ;
        RECT 421.345 -283.890 421.515 -280.920 ;
        RECT 419.775 -284.325 420.480 -284.130 ;
        RECT 420.265 -284.385 420.480 -284.325 ;
        RECT 419.055 -284.545 419.830 -284.495 ;
        RECT 417.030 -284.725 419.830 -284.545 ;
        RECT 417.030 -284.735 417.380 -284.725 ;
        RECT 419.055 -284.770 419.830 -284.725 ;
        RECT 420.265 -284.660 421.170 -284.385 ;
        RECT 420.265 -285.010 420.480 -284.660 ;
        RECT 417.705 -285.080 418.480 -285.035 ;
        RECT 417.520 -285.250 418.480 -285.080 ;
        RECT 417.705 -285.310 418.480 -285.250 ;
        RECT 418.710 -285.210 420.480 -285.010 ;
        RECT 421.340 -285.110 421.555 -283.890 ;
        RECT 422.525 -284.235 422.875 -277.550 ;
        RECT 429.105 -280.030 430.710 -279.860 ;
        RECT 428.210 -282.710 428.380 -280.210 ;
        RECT 428.205 -282.940 428.380 -282.710 ;
        RECT 429.105 -282.940 429.305 -280.030 ;
        RECT 429.550 -280.230 429.725 -280.030 ;
        RECT 429.555 -282.750 429.725 -280.230 ;
        RECT 430.045 -282.715 430.215 -280.210 ;
        RECT 430.535 -280.225 430.710 -280.030 ;
        RECT 428.205 -283.140 429.305 -282.940 ;
        RECT 430.030 -283.315 430.220 -282.715 ;
        RECT 430.535 -282.750 430.705 -280.225 ;
        RECT 431.185 -283.130 431.355 -280.210 ;
        RECT 432.815 -282.780 432.985 -280.210 ;
        RECT 433.955 -281.660 434.125 -280.210 ;
        RECT 433.950 -282.125 434.135 -281.660 ;
        RECT 433.950 -282.310 434.635 -282.125 ;
        RECT 432.815 -282.950 433.610 -282.780 ;
        RECT 431.930 -283.130 432.620 -283.075 ;
        RECT 428.210 -283.505 430.220 -283.315 ;
        RECT 430.555 -283.300 432.620 -283.130 ;
        RECT 427.025 -283.560 427.715 -283.510 ;
        RECT 425.075 -283.730 427.715 -283.560 ;
        RECT 422.470 -284.595 422.995 -284.235 ;
        RECT 425.075 -285.110 425.290 -283.730 ;
        RECT 427.025 -283.780 427.715 -283.730 ;
        RECT 427.305 -284.235 427.995 -284.190 ;
        RECT 426.255 -284.405 427.995 -284.235 ;
        RECT 426.255 -285.040 426.615 -284.405 ;
        RECT 427.305 -284.460 427.995 -284.405 ;
        RECT 426.255 -285.085 426.675 -285.040 ;
        RECT 412.635 -285.850 414.885 -285.760 ;
        RECT 410.425 -286.065 414.885 -285.850 ;
        RECT 410.425 -286.155 412.670 -286.065 ;
        RECT 414.580 -287.540 414.885 -286.065 ;
        RECT 418.250 -286.950 418.420 -285.480 ;
        RECT 418.710 -285.560 418.935 -285.210 ;
        RECT 420.670 -285.310 425.290 -285.110 ;
        RECT 420.910 -285.325 425.290 -285.310 ;
        RECT 418.215 -287.540 418.450 -286.950 ;
        RECT 418.740 -287.020 418.910 -285.560 ;
        RECT 419.230 -286.945 419.400 -285.480 ;
        RECT 420.440 -286.895 420.610 -285.480 ;
        RECT 420.910 -285.525 421.130 -285.325 ;
        RECT 426.280 -285.435 426.675 -285.085 ;
        RECT 419.195 -287.540 419.430 -286.945 ;
        RECT 420.405 -287.540 420.640 -286.895 ;
        RECT 420.930 -287.020 421.100 -285.525 ;
        RECT 427.720 -286.645 427.890 -285.190 ;
        RECT 427.710 -287.200 427.895 -286.645 ;
        RECT 428.210 -286.730 428.380 -283.505 ;
        RECT 429.355 -283.855 429.545 -283.505 ;
        RECT 430.555 -283.695 430.725 -283.300 ;
        RECT 431.930 -283.345 432.620 -283.300 ;
        RECT 429.305 -284.545 429.575 -283.855 ;
        RECT 430.070 -283.865 430.725 -283.695 ;
        RECT 431.055 -283.780 431.745 -283.510 ;
        RECT 432.980 -283.855 433.250 -283.165 ;
        RECT 433.440 -283.170 433.610 -282.950 ;
        RECT 433.440 -283.440 434.270 -283.170 ;
        RECT 430.070 -286.730 430.240 -283.865 ;
        RECT 433.440 -284.015 433.610 -283.440 ;
        RECT 433.870 -284.015 434.140 -283.930 ;
        RECT 430.560 -284.210 431.355 -284.035 ;
        RECT 433.440 -284.040 434.140 -284.015 ;
        RECT 433.300 -284.185 434.140 -284.040 ;
        RECT 430.560 -286.730 430.730 -284.210 ;
        RECT 431.185 -286.730 431.355 -284.210 ;
        RECT 431.675 -286.645 431.845 -284.190 ;
        RECT 432.325 -286.640 432.495 -284.190 ;
        RECT 425.025 -287.220 428.080 -287.200 ;
        RECT 431.670 -287.220 431.855 -286.645 ;
        RECT 432.310 -287.220 432.495 -286.640 ;
        RECT 432.815 -286.730 432.985 -284.190 ;
        RECT 433.300 -284.210 433.610 -284.185 ;
        RECT 433.305 -286.730 433.475 -284.210 ;
        RECT 433.870 -284.225 434.140 -284.185 ;
        RECT 434.445 -284.775 434.635 -282.310 ;
        RECT 434.445 -284.965 435.905 -284.775 ;
        RECT 433.955 -286.635 434.125 -285.190 ;
        RECT 434.445 -285.215 434.635 -284.965 ;
        RECT 433.945 -287.220 434.130 -286.635 ;
        RECT 434.445 -286.730 434.615 -285.215 ;
        RECT 425.025 -287.540 434.695 -287.220 ;
        RECT 414.580 -287.765 434.695 -287.540 ;
        RECT 414.580 -288.105 425.590 -287.765 ;
        RECT 427.330 -288.025 434.695 -287.765 ;
        RECT 334.385 -291.795 334.575 -289.905 ;
        RECT 359.095 -289.980 379.020 -289.660 ;
        RECT 340.420 -291.400 343.745 -291.260 ;
        RECT 340.420 -291.690 345.595 -291.400 ;
        RECT 334.270 -292.065 334.635 -291.795 ;
        RECT 340.420 -292.095 340.850 -291.690 ;
        RECT 341.720 -291.875 341.895 -291.690 ;
        RECT 343.345 -291.705 345.595 -291.690 ;
        RECT 336.160 -292.525 340.850 -292.095 ;
        RECT 335.400 -293.645 336.050 -293.515 ;
        RECT 332.875 -293.975 336.050 -293.645 ;
        RECT 336.860 -293.805 337.030 -292.525 ;
        RECT 337.350 -293.805 337.520 -292.765 ;
        RECT 337.840 -293.805 338.010 -292.525 ;
        RECT 338.330 -293.635 338.500 -292.765 ;
        RECT 341.235 -293.415 341.405 -291.875 ;
        RECT 341.725 -293.415 341.895 -291.875 ;
        RECT 342.215 -293.415 342.385 -291.875 ;
        RECT 342.705 -293.415 342.875 -291.875 ;
        RECT 343.195 -293.415 343.365 -291.875 ;
        RECT 341.075 -293.630 341.430 -293.625 ;
        RECT 343.135 -293.630 343.505 -293.600 ;
        RECT 341.075 -293.635 343.505 -293.630 ;
        RECT 338.330 -293.805 343.505 -293.635 ;
        RECT 345.290 -293.740 345.595 -291.705 ;
        RECT 338.335 -293.825 343.505 -293.805 ;
        RECT 338.335 -293.835 341.080 -293.825 ;
        RECT 336.270 -293.975 336.635 -293.945 ;
        RECT 343.135 -293.955 343.505 -293.825 ;
        RECT 332.875 -294.025 336.635 -293.975 ;
        RECT 335.400 -294.180 336.635 -294.025 ;
        RECT 340.810 -294.115 341.485 -294.075 ;
        RECT 340.710 -294.125 341.485 -294.115 ;
        RECT 335.400 -294.265 336.050 -294.180 ;
        RECT 336.270 -294.245 336.635 -294.180 ;
        RECT 335.535 -294.515 335.915 -294.265 ;
        RECT 339.675 -294.305 341.485 -294.125 ;
        RECT 344.070 -294.170 347.995 -293.740 ;
        RECT 340.710 -294.315 341.485 -294.305 ;
        RECT 340.810 -294.345 341.485 -294.315 ;
        RECT 341.725 -294.230 343.820 -294.190 ;
        RECT 341.725 -294.380 343.875 -294.230 ;
        RECT 336.860 -295.455 337.030 -294.415 ;
        RECT 337.840 -295.455 338.010 -294.415 ;
        RECT 338.820 -295.455 338.990 -294.415 ;
        RECT 341.725 -296.100 341.895 -294.380 ;
        RECT 342.705 -296.100 342.875 -294.380 ;
        RECT 343.570 -295.125 343.875 -294.380 ;
        RECT 344.770 -294.950 344.940 -294.170 ;
        RECT 345.260 -294.950 345.430 -294.410 ;
        RECT 345.750 -294.950 345.920 -294.170 ;
        RECT 346.240 -294.950 346.410 -294.410 ;
        RECT 344.180 -295.125 344.545 -295.095 ;
        RECT 343.570 -295.190 344.545 -295.125 ;
        RECT 343.680 -295.330 344.545 -295.190 ;
        RECT 344.180 -295.395 344.545 -295.330 ;
        RECT 346.730 -295.245 348.590 -294.895 ;
        RECT 344.770 -296.105 344.940 -295.565 ;
        RECT 345.750 -296.105 345.920 -295.565 ;
        RECT 346.730 -296.105 346.900 -295.245 ;
        RECT 345.000 -298.445 346.200 -298.275 ;
        RECT 336.730 -300.780 336.900 -299.060 ;
        RECT 337.710 -300.780 337.880 -299.060 ;
        RECT 339.775 -299.595 339.945 -299.055 ;
        RECT 340.755 -299.595 340.925 -299.055 ;
        RECT 339.185 -299.830 339.550 -299.765 ;
        RECT 338.685 -299.970 339.550 -299.830 ;
        RECT 338.575 -300.035 339.550 -299.970 ;
        RECT 338.575 -300.780 338.880 -300.035 ;
        RECT 339.185 -300.065 339.550 -300.035 ;
        RECT 341.735 -299.915 341.905 -299.055 ;
        RECT 335.815 -300.845 336.490 -300.815 ;
        RECT 335.715 -300.855 336.490 -300.845 ;
        RECT 333.645 -301.035 336.490 -300.855 ;
        RECT 336.730 -300.930 338.880 -300.780 ;
        RECT 336.730 -300.970 338.825 -300.930 ;
        RECT 339.775 -300.990 339.945 -300.210 ;
        RECT 340.265 -300.750 340.435 -300.210 ;
        RECT 340.755 -300.990 340.925 -300.210 ;
        RECT 341.245 -300.750 341.415 -300.210 ;
        RECT 341.735 -300.265 343.125 -299.915 ;
        RECT 331.240 -301.620 332.665 -301.405 ;
        RECT 329.845 -302.135 330.370 -301.775 ;
        RECT 332.450 -302.650 332.665 -301.620 ;
        RECT 320.010 -303.390 322.260 -303.300 ;
        RECT 317.800 -303.605 322.260 -303.390 ;
        RECT 317.800 -303.695 320.045 -303.605 ;
        RECT 321.955 -305.080 322.260 -303.605 ;
        RECT 325.625 -304.490 325.795 -303.020 ;
        RECT 326.085 -303.100 326.310 -302.750 ;
        RECT 328.045 -302.850 332.665 -302.650 ;
        RECT 328.285 -302.865 332.665 -302.850 ;
        RECT 325.590 -305.080 325.825 -304.490 ;
        RECT 326.115 -304.560 326.285 -303.100 ;
        RECT 326.605 -304.485 326.775 -303.020 ;
        RECT 327.815 -304.435 327.985 -303.020 ;
        RECT 328.285 -303.065 328.505 -302.865 ;
        RECT 326.570 -305.080 326.805 -304.485 ;
        RECT 327.780 -305.080 328.015 -304.435 ;
        RECT 328.305 -304.560 328.475 -303.065 ;
        RECT 321.955 -305.645 329.340 -305.080 ;
        RECT 333.645 -306.015 334.325 -301.035 ;
        RECT 335.715 -301.045 336.490 -301.035 ;
        RECT 335.815 -301.085 336.490 -301.045 ;
        RECT 334.950 -301.335 336.085 -301.325 ;
        RECT 338.140 -301.335 338.510 -301.205 ;
        RECT 334.950 -301.525 338.510 -301.335 ;
        RECT 339.075 -301.420 342.150 -300.990 ;
        RECT 336.080 -301.530 338.510 -301.525 ;
        RECT 336.080 -301.535 336.435 -301.530 ;
        RECT 338.140 -301.560 338.510 -301.530 ;
        RECT 336.240 -303.285 336.410 -301.745 ;
        RECT 336.730 -303.285 336.900 -301.745 ;
        RECT 337.220 -303.285 337.390 -301.745 ;
        RECT 337.710 -303.285 337.880 -301.745 ;
        RECT 338.200 -303.285 338.370 -301.745 ;
        RECT 336.725 -303.545 336.900 -303.285 ;
        RECT 340.295 -303.455 340.600 -301.420 ;
        RECT 342.745 -302.240 343.095 -300.265 ;
        RECT 343.965 -301.535 344.135 -298.615 ;
        RECT 345.000 -298.655 345.210 -298.445 ;
        RECT 343.945 -301.830 344.155 -301.535 ;
        RECT 345.020 -301.565 345.190 -298.655 ;
        RECT 345.510 -301.555 345.680 -298.615 ;
        RECT 345.990 -298.665 346.200 -298.445 ;
        RECT 345.005 -301.830 345.215 -301.565 ;
        RECT 343.945 -302.010 345.215 -301.830 ;
        RECT 345.490 -301.825 345.700 -301.555 ;
        RECT 346.000 -301.655 346.170 -298.665 ;
        RECT 347.060 -301.585 347.230 -298.615 ;
        RECT 345.490 -302.020 346.195 -301.825 ;
        RECT 345.980 -302.080 346.195 -302.020 ;
        RECT 344.770 -302.240 345.545 -302.190 ;
        RECT 342.745 -302.420 345.545 -302.240 ;
        RECT 342.745 -302.430 343.095 -302.420 ;
        RECT 344.770 -302.465 345.545 -302.420 ;
        RECT 345.980 -302.355 346.885 -302.080 ;
        RECT 345.980 -302.705 346.195 -302.355 ;
        RECT 343.420 -302.775 344.195 -302.730 ;
        RECT 343.235 -302.945 344.195 -302.775 ;
        RECT 343.420 -303.005 344.195 -302.945 ;
        RECT 344.425 -302.905 346.195 -302.705 ;
        RECT 347.055 -302.805 347.270 -301.585 ;
        RECT 348.240 -301.930 348.590 -295.245 ;
        RECT 348.185 -302.290 348.710 -301.930 ;
        RECT 350.530 -302.805 351.835 -302.000 ;
        RECT 338.350 -303.545 340.600 -303.455 ;
        RECT 336.140 -303.760 340.600 -303.545 ;
        RECT 336.140 -303.850 338.385 -303.760 ;
        RECT 340.295 -305.235 340.600 -303.760 ;
        RECT 343.965 -304.645 344.135 -303.175 ;
        RECT 344.425 -303.255 344.650 -302.905 ;
        RECT 346.385 -303.005 352.395 -302.805 ;
        RECT 346.625 -303.020 352.395 -303.005 ;
        RECT 343.930 -305.235 344.165 -304.645 ;
        RECT 344.455 -304.715 344.625 -303.255 ;
        RECT 344.945 -304.640 345.115 -303.175 ;
        RECT 346.155 -304.590 346.325 -303.175 ;
        RECT 346.625 -303.220 346.845 -303.020 ;
        RECT 344.910 -305.235 345.145 -304.640 ;
        RECT 346.120 -305.235 346.355 -304.590 ;
        RECT 346.645 -304.715 346.815 -303.220 ;
        RECT 350.530 -303.520 351.835 -303.020 ;
        RECT 340.295 -305.800 347.680 -305.235 ;
        RECT 315.650 -306.695 334.325 -306.015 ;
        RECT 215.060 -314.155 216.260 -314.110 ;
        RECT 312.855 -314.275 314.575 -312.860 ;
        RECT 48.450 -317.940 49.130 -317.930 ;
        RECT 315.650 -317.940 316.330 -306.695 ;
        RECT 359.095 -309.160 359.945 -289.980 ;
        RECT 362.470 -290.040 379.020 -289.980 ;
        RECT 362.470 -290.950 362.850 -290.040 ;
        RECT 362.470 -291.330 363.180 -290.950 ;
        RECT 362.800 -293.275 363.180 -291.330 ;
        RECT 367.845 -291.160 371.170 -291.020 ;
        RECT 367.845 -291.450 373.020 -291.160 ;
        RECT 376.890 -291.445 377.350 -291.020 ;
        RECT 367.845 -291.855 368.275 -291.450 ;
        RECT 369.145 -291.635 369.320 -291.450 ;
        RECT 370.770 -291.465 373.020 -291.450 ;
        RECT 363.585 -292.285 368.275 -291.855 ;
        RECT 362.800 -293.735 363.475 -293.275 ;
        RECT 364.285 -293.565 364.455 -292.285 ;
        RECT 364.775 -293.565 364.945 -292.525 ;
        RECT 365.265 -293.565 365.435 -292.285 ;
        RECT 365.755 -293.395 365.925 -292.525 ;
        RECT 368.660 -293.175 368.830 -291.635 ;
        RECT 369.150 -293.175 369.320 -291.635 ;
        RECT 369.640 -293.175 369.810 -291.635 ;
        RECT 370.130 -293.175 370.300 -291.635 ;
        RECT 370.620 -293.175 370.790 -291.635 ;
        RECT 368.500 -293.390 368.855 -293.385 ;
        RECT 370.560 -293.390 370.930 -293.360 ;
        RECT 368.500 -293.395 370.930 -293.390 ;
        RECT 365.755 -293.565 370.930 -293.395 ;
        RECT 372.715 -293.500 373.020 -291.465 ;
        RECT 365.760 -293.585 370.930 -293.565 ;
        RECT 365.760 -293.595 368.505 -293.585 ;
        RECT 363.695 -293.735 364.060 -293.705 ;
        RECT 370.560 -293.715 370.930 -293.585 ;
        RECT 362.800 -293.820 364.060 -293.735 ;
        RECT 362.825 -293.940 364.060 -293.820 ;
        RECT 368.235 -293.875 368.910 -293.835 ;
        RECT 368.135 -293.885 368.910 -293.875 ;
        RECT 362.825 -294.025 363.475 -293.940 ;
        RECT 363.695 -294.005 364.060 -293.940 ;
        RECT 367.100 -294.065 368.910 -293.885 ;
        RECT 371.495 -293.930 375.420 -293.500 ;
        RECT 368.135 -294.075 368.910 -294.065 ;
        RECT 368.235 -294.105 368.910 -294.075 ;
        RECT 369.150 -293.990 371.245 -293.950 ;
        RECT 369.150 -294.140 371.300 -293.990 ;
        RECT 364.285 -295.215 364.455 -294.175 ;
        RECT 365.265 -295.215 365.435 -294.175 ;
        RECT 366.245 -295.215 366.415 -294.175 ;
        RECT 369.150 -295.860 369.320 -294.140 ;
        RECT 370.130 -295.860 370.300 -294.140 ;
        RECT 370.995 -294.885 371.300 -294.140 ;
        RECT 372.195 -294.710 372.365 -293.930 ;
        RECT 372.685 -294.710 372.855 -294.170 ;
        RECT 373.175 -294.710 373.345 -293.930 ;
        RECT 373.665 -294.710 373.835 -294.170 ;
        RECT 371.605 -294.885 371.970 -294.855 ;
        RECT 370.995 -294.950 371.970 -294.885 ;
        RECT 371.105 -295.090 371.970 -294.950 ;
        RECT 371.605 -295.155 371.970 -295.090 ;
        RECT 374.155 -295.005 376.015 -294.655 ;
        RECT 372.195 -295.865 372.365 -295.325 ;
        RECT 373.175 -295.865 373.345 -295.325 ;
        RECT 374.155 -295.865 374.325 -295.005 ;
        RECT 372.425 -298.205 373.625 -298.035 ;
        RECT 364.155 -300.540 364.325 -298.820 ;
        RECT 365.135 -300.540 365.305 -298.820 ;
        RECT 367.200 -299.355 367.370 -298.815 ;
        RECT 368.180 -299.355 368.350 -298.815 ;
        RECT 366.610 -299.590 366.975 -299.525 ;
        RECT 366.110 -299.730 366.975 -299.590 ;
        RECT 366.000 -299.795 366.975 -299.730 ;
        RECT 366.000 -300.540 366.305 -299.795 ;
        RECT 366.610 -299.825 366.975 -299.795 ;
        RECT 369.160 -299.675 369.330 -298.815 ;
        RECT 363.240 -300.605 363.915 -300.575 ;
        RECT 363.140 -300.615 363.915 -300.605 ;
        RECT 360.500 -300.795 363.915 -300.615 ;
        RECT 364.155 -300.690 366.305 -300.540 ;
        RECT 364.155 -300.730 366.250 -300.690 ;
        RECT 367.200 -300.750 367.370 -299.970 ;
        RECT 367.690 -300.510 367.860 -299.970 ;
        RECT 368.180 -300.750 368.350 -299.970 ;
        RECT 368.670 -300.510 368.840 -299.970 ;
        RECT 369.160 -300.025 370.550 -299.675 ;
        RECT 361.415 -305.930 362.095 -300.795 ;
        RECT 363.140 -300.805 363.915 -300.795 ;
        RECT 363.240 -300.845 363.915 -300.805 ;
        RECT 362.375 -301.095 363.510 -301.085 ;
        RECT 365.565 -301.095 365.935 -300.965 ;
        RECT 362.375 -301.285 365.935 -301.095 ;
        RECT 366.500 -301.180 369.575 -300.750 ;
        RECT 363.505 -301.290 365.935 -301.285 ;
        RECT 363.505 -301.295 363.860 -301.290 ;
        RECT 365.565 -301.320 365.935 -301.290 ;
        RECT 363.665 -303.045 363.835 -301.505 ;
        RECT 364.155 -303.045 364.325 -301.505 ;
        RECT 364.645 -303.045 364.815 -301.505 ;
        RECT 365.135 -303.045 365.305 -301.505 ;
        RECT 365.625 -303.045 365.795 -301.505 ;
        RECT 364.150 -303.305 364.325 -303.045 ;
        RECT 367.720 -303.215 368.025 -301.180 ;
        RECT 370.170 -302.000 370.520 -300.025 ;
        RECT 371.390 -301.295 371.560 -298.375 ;
        RECT 372.425 -298.415 372.635 -298.205 ;
        RECT 371.370 -301.590 371.580 -301.295 ;
        RECT 372.445 -301.325 372.615 -298.415 ;
        RECT 372.935 -301.315 373.105 -298.375 ;
        RECT 373.415 -298.425 373.625 -298.205 ;
        RECT 372.430 -301.590 372.640 -301.325 ;
        RECT 371.370 -301.770 372.640 -301.590 ;
        RECT 372.915 -301.585 373.125 -301.315 ;
        RECT 373.425 -301.415 373.595 -298.425 ;
        RECT 374.485 -301.345 374.655 -298.375 ;
        RECT 372.915 -301.780 373.620 -301.585 ;
        RECT 373.405 -301.840 373.620 -301.780 ;
        RECT 372.195 -302.000 372.970 -301.950 ;
        RECT 370.170 -302.180 372.970 -302.000 ;
        RECT 370.170 -302.190 370.520 -302.180 ;
        RECT 372.195 -302.225 372.970 -302.180 ;
        RECT 373.405 -302.115 374.310 -301.840 ;
        RECT 373.405 -302.465 373.620 -302.115 ;
        RECT 370.845 -302.535 371.620 -302.490 ;
        RECT 370.660 -302.705 371.620 -302.535 ;
        RECT 370.845 -302.765 371.620 -302.705 ;
        RECT 371.850 -302.665 373.620 -302.465 ;
        RECT 374.480 -302.565 374.695 -301.345 ;
        RECT 375.665 -301.690 376.015 -295.005 ;
        RECT 377.005 -301.320 377.220 -291.445 ;
        RECT 378.640 -293.560 379.020 -290.040 ;
        RECT 380.150 -289.820 389.085 -289.630 ;
        RECT 405.475 -289.470 409.880 -288.735 ;
        RECT 435.715 -289.440 435.905 -284.965 ;
        RECT 380.150 -291.710 380.340 -289.820 ;
        RECT 405.475 -289.850 425.840 -289.470 ;
        RECT 405.475 -289.865 409.880 -289.850 ;
        RECT 386.185 -291.315 389.510 -291.175 ;
        RECT 386.185 -291.605 391.360 -291.315 ;
        RECT 380.035 -291.980 380.400 -291.710 ;
        RECT 386.185 -292.010 386.615 -291.605 ;
        RECT 387.485 -291.790 387.660 -291.605 ;
        RECT 389.110 -291.620 391.360 -291.605 ;
        RECT 381.925 -292.440 386.615 -292.010 ;
        RECT 381.165 -293.560 381.815 -293.430 ;
        RECT 378.640 -293.890 381.815 -293.560 ;
        RECT 382.625 -293.720 382.795 -292.440 ;
        RECT 383.115 -293.720 383.285 -292.680 ;
        RECT 383.605 -293.720 383.775 -292.440 ;
        RECT 384.095 -293.550 384.265 -292.680 ;
        RECT 387.000 -293.330 387.170 -291.790 ;
        RECT 387.490 -293.330 387.660 -291.790 ;
        RECT 387.980 -293.330 388.150 -291.790 ;
        RECT 388.470 -293.330 388.640 -291.790 ;
        RECT 388.960 -293.330 389.130 -291.790 ;
        RECT 386.840 -293.545 387.195 -293.540 ;
        RECT 388.900 -293.545 389.270 -293.515 ;
        RECT 386.840 -293.550 389.270 -293.545 ;
        RECT 384.095 -293.720 389.270 -293.550 ;
        RECT 391.055 -293.655 391.360 -291.620 ;
        RECT 384.100 -293.740 389.270 -293.720 ;
        RECT 384.100 -293.750 386.845 -293.740 ;
        RECT 382.035 -293.890 382.400 -293.860 ;
        RECT 388.900 -293.870 389.270 -293.740 ;
        RECT 378.640 -293.940 382.400 -293.890 ;
        RECT 381.165 -294.095 382.400 -293.940 ;
        RECT 386.575 -294.030 387.250 -293.990 ;
        RECT 386.475 -294.040 387.250 -294.030 ;
        RECT 381.165 -294.180 381.815 -294.095 ;
        RECT 382.035 -294.160 382.400 -294.095 ;
        RECT 381.300 -294.430 381.680 -294.180 ;
        RECT 385.440 -294.220 387.250 -294.040 ;
        RECT 389.835 -294.085 393.760 -293.655 ;
        RECT 386.475 -294.230 387.250 -294.220 ;
        RECT 386.575 -294.260 387.250 -294.230 ;
        RECT 387.490 -294.145 389.585 -294.105 ;
        RECT 387.490 -294.295 389.640 -294.145 ;
        RECT 382.625 -295.370 382.795 -294.330 ;
        RECT 383.605 -295.370 383.775 -294.330 ;
        RECT 384.585 -295.370 384.755 -294.330 ;
        RECT 387.490 -296.015 387.660 -294.295 ;
        RECT 388.470 -296.015 388.640 -294.295 ;
        RECT 389.335 -295.040 389.640 -294.295 ;
        RECT 390.535 -294.865 390.705 -294.085 ;
        RECT 391.025 -294.865 391.195 -294.325 ;
        RECT 391.515 -294.865 391.685 -294.085 ;
        RECT 392.005 -294.865 392.175 -294.325 ;
        RECT 389.945 -295.040 390.310 -295.010 ;
        RECT 389.335 -295.105 390.310 -295.040 ;
        RECT 389.445 -295.245 390.310 -295.105 ;
        RECT 389.945 -295.310 390.310 -295.245 ;
        RECT 392.495 -295.160 394.355 -294.810 ;
        RECT 390.535 -296.020 390.705 -295.480 ;
        RECT 391.515 -296.020 391.685 -295.480 ;
        RECT 392.495 -296.020 392.665 -295.160 ;
        RECT 390.765 -298.360 391.965 -298.190 ;
        RECT 382.495 -300.695 382.665 -298.975 ;
        RECT 383.475 -300.695 383.645 -298.975 ;
        RECT 385.540 -299.510 385.710 -298.970 ;
        RECT 386.520 -299.510 386.690 -298.970 ;
        RECT 384.950 -299.745 385.315 -299.680 ;
        RECT 384.450 -299.885 385.315 -299.745 ;
        RECT 384.340 -299.950 385.315 -299.885 ;
        RECT 384.340 -300.695 384.645 -299.950 ;
        RECT 384.950 -299.980 385.315 -299.950 ;
        RECT 387.500 -299.830 387.670 -298.970 ;
        RECT 381.580 -300.760 382.255 -300.730 ;
        RECT 381.480 -300.770 382.255 -300.760 ;
        RECT 379.410 -300.950 382.255 -300.770 ;
        RECT 382.495 -300.845 384.645 -300.695 ;
        RECT 382.495 -300.885 384.590 -300.845 ;
        RECT 385.540 -300.905 385.710 -300.125 ;
        RECT 386.030 -300.665 386.200 -300.125 ;
        RECT 386.520 -300.905 386.690 -300.125 ;
        RECT 387.010 -300.665 387.180 -300.125 ;
        RECT 387.500 -300.180 388.890 -299.830 ;
        RECT 377.005 -301.535 378.430 -301.320 ;
        RECT 375.610 -302.050 376.135 -301.690 ;
        RECT 378.215 -302.565 378.430 -301.535 ;
        RECT 365.775 -303.305 368.025 -303.215 ;
        RECT 363.565 -303.520 368.025 -303.305 ;
        RECT 363.565 -303.610 365.810 -303.520 ;
        RECT 367.720 -304.995 368.025 -303.520 ;
        RECT 371.390 -304.405 371.560 -302.935 ;
        RECT 371.850 -303.015 372.075 -302.665 ;
        RECT 373.810 -302.765 378.430 -302.565 ;
        RECT 374.050 -302.780 378.430 -302.765 ;
        RECT 371.355 -304.995 371.590 -304.405 ;
        RECT 371.880 -304.475 372.050 -303.015 ;
        RECT 372.370 -304.400 372.540 -302.935 ;
        RECT 373.580 -304.350 373.750 -302.935 ;
        RECT 374.050 -302.980 374.270 -302.780 ;
        RECT 372.335 -304.995 372.570 -304.400 ;
        RECT 373.545 -304.995 373.780 -304.350 ;
        RECT 374.070 -304.475 374.240 -302.980 ;
        RECT 367.720 -305.560 375.105 -304.995 ;
        RECT 379.410 -305.930 380.090 -300.950 ;
        RECT 381.480 -300.960 382.255 -300.950 ;
        RECT 381.580 -301.000 382.255 -300.960 ;
        RECT 380.715 -301.250 381.850 -301.240 ;
        RECT 383.905 -301.250 384.275 -301.120 ;
        RECT 380.715 -301.440 384.275 -301.250 ;
        RECT 384.840 -301.335 387.915 -300.905 ;
        RECT 381.845 -301.445 384.275 -301.440 ;
        RECT 381.845 -301.450 382.200 -301.445 ;
        RECT 383.905 -301.475 384.275 -301.445 ;
        RECT 382.005 -303.200 382.175 -301.660 ;
        RECT 382.495 -303.200 382.665 -301.660 ;
        RECT 382.985 -303.200 383.155 -301.660 ;
        RECT 383.475 -303.200 383.645 -301.660 ;
        RECT 383.965 -303.200 384.135 -301.660 ;
        RECT 382.490 -303.460 382.665 -303.200 ;
        RECT 386.060 -303.370 386.365 -301.335 ;
        RECT 388.510 -302.155 388.860 -300.180 ;
        RECT 389.730 -301.450 389.900 -298.530 ;
        RECT 390.765 -298.570 390.975 -298.360 ;
        RECT 389.710 -301.745 389.920 -301.450 ;
        RECT 390.785 -301.480 390.955 -298.570 ;
        RECT 391.275 -301.470 391.445 -298.530 ;
        RECT 391.755 -298.580 391.965 -298.360 ;
        RECT 390.770 -301.745 390.980 -301.480 ;
        RECT 389.710 -301.925 390.980 -301.745 ;
        RECT 391.255 -301.740 391.465 -301.470 ;
        RECT 391.765 -301.570 391.935 -298.580 ;
        RECT 392.825 -301.500 392.995 -298.530 ;
        RECT 391.255 -301.935 391.960 -301.740 ;
        RECT 391.745 -301.995 391.960 -301.935 ;
        RECT 390.535 -302.155 391.310 -302.105 ;
        RECT 388.510 -302.335 391.310 -302.155 ;
        RECT 388.510 -302.345 388.860 -302.335 ;
        RECT 390.535 -302.380 391.310 -302.335 ;
        RECT 391.745 -302.270 392.650 -301.995 ;
        RECT 391.745 -302.620 391.960 -302.270 ;
        RECT 389.185 -302.690 389.960 -302.645 ;
        RECT 389.000 -302.860 389.960 -302.690 ;
        RECT 389.185 -302.920 389.960 -302.860 ;
        RECT 390.190 -302.820 391.960 -302.620 ;
        RECT 392.820 -302.720 393.035 -301.500 ;
        RECT 394.005 -301.845 394.355 -295.160 ;
        RECT 393.950 -302.205 394.475 -301.845 ;
        RECT 396.960 -302.720 397.470 -302.530 ;
        RECT 384.115 -303.460 386.365 -303.370 ;
        RECT 381.905 -303.675 386.365 -303.460 ;
        RECT 381.905 -303.765 384.150 -303.675 ;
        RECT 386.060 -305.150 386.365 -303.675 ;
        RECT 389.730 -304.560 389.900 -303.090 ;
        RECT 390.190 -303.170 390.415 -302.820 ;
        RECT 392.150 -302.920 398.160 -302.720 ;
        RECT 392.390 -302.935 398.160 -302.920 ;
        RECT 389.695 -305.150 389.930 -304.560 ;
        RECT 390.220 -304.630 390.390 -303.170 ;
        RECT 390.710 -304.555 390.880 -303.090 ;
        RECT 391.920 -304.505 392.090 -303.090 ;
        RECT 392.390 -303.135 392.610 -302.935 ;
        RECT 396.960 -303.085 397.470 -302.935 ;
        RECT 390.675 -305.150 390.910 -304.555 ;
        RECT 391.885 -305.150 392.120 -304.505 ;
        RECT 392.410 -304.630 392.580 -303.135 ;
        RECT 386.060 -305.715 393.445 -305.150 ;
        RECT 361.415 -306.610 380.090 -305.930 ;
        RECT 358.900 -310.060 360.130 -309.160 ;
        RECT -119.230 -318.620 316.330 -317.940 ;
        RECT -119.230 -318.645 -107.700 -318.620 ;
        RECT -119.230 -319.435 -118.550 -318.645 ;
        RECT 361.415 -319.435 362.095 -306.610 ;
        RECT 405.475 -312.875 406.605 -289.865 ;
        RECT 409.290 -290.760 409.670 -289.865 ;
        RECT 409.290 -291.140 410.000 -290.760 ;
        RECT 409.620 -293.085 410.000 -291.140 ;
        RECT 414.665 -290.970 417.990 -290.830 ;
        RECT 414.665 -291.260 419.840 -290.970 ;
        RECT 423.710 -291.255 424.170 -290.830 ;
        RECT 414.665 -291.665 415.095 -291.260 ;
        RECT 415.965 -291.445 416.140 -291.260 ;
        RECT 417.590 -291.275 419.840 -291.260 ;
        RECT 410.405 -292.095 415.095 -291.665 ;
        RECT 409.620 -293.545 410.295 -293.085 ;
        RECT 411.105 -293.375 411.275 -292.095 ;
        RECT 411.595 -293.375 411.765 -292.335 ;
        RECT 412.085 -293.375 412.255 -292.095 ;
        RECT 412.575 -293.205 412.745 -292.335 ;
        RECT 415.480 -292.985 415.650 -291.445 ;
        RECT 415.970 -292.985 416.140 -291.445 ;
        RECT 416.460 -292.985 416.630 -291.445 ;
        RECT 416.950 -292.985 417.120 -291.445 ;
        RECT 417.440 -292.985 417.610 -291.445 ;
        RECT 415.320 -293.200 415.675 -293.195 ;
        RECT 417.380 -293.200 417.750 -293.170 ;
        RECT 415.320 -293.205 417.750 -293.200 ;
        RECT 412.575 -293.375 417.750 -293.205 ;
        RECT 419.535 -293.310 419.840 -291.275 ;
        RECT 412.580 -293.395 417.750 -293.375 ;
        RECT 412.580 -293.405 415.325 -293.395 ;
        RECT 410.515 -293.545 410.880 -293.515 ;
        RECT 417.380 -293.525 417.750 -293.395 ;
        RECT 409.620 -293.630 410.880 -293.545 ;
        RECT 409.645 -293.750 410.880 -293.630 ;
        RECT 415.055 -293.685 415.730 -293.645 ;
        RECT 414.955 -293.695 415.730 -293.685 ;
        RECT 409.645 -293.835 410.295 -293.750 ;
        RECT 410.515 -293.815 410.880 -293.750 ;
        RECT 413.920 -293.875 415.730 -293.695 ;
        RECT 418.315 -293.740 422.240 -293.310 ;
        RECT 414.955 -293.885 415.730 -293.875 ;
        RECT 415.055 -293.915 415.730 -293.885 ;
        RECT 415.970 -293.800 418.065 -293.760 ;
        RECT 415.970 -293.950 418.120 -293.800 ;
        RECT 411.105 -295.025 411.275 -293.985 ;
        RECT 412.085 -295.025 412.255 -293.985 ;
        RECT 413.065 -295.025 413.235 -293.985 ;
        RECT 415.970 -295.670 416.140 -293.950 ;
        RECT 416.950 -295.670 417.120 -293.950 ;
        RECT 417.815 -294.695 418.120 -293.950 ;
        RECT 419.015 -294.520 419.185 -293.740 ;
        RECT 419.505 -294.520 419.675 -293.980 ;
        RECT 419.995 -294.520 420.165 -293.740 ;
        RECT 420.485 -294.520 420.655 -293.980 ;
        RECT 418.425 -294.695 418.790 -294.665 ;
        RECT 417.815 -294.760 418.790 -294.695 ;
        RECT 417.925 -294.900 418.790 -294.760 ;
        RECT 418.425 -294.965 418.790 -294.900 ;
        RECT 420.975 -294.815 422.835 -294.465 ;
        RECT 419.015 -295.675 419.185 -295.135 ;
        RECT 419.995 -295.675 420.165 -295.135 ;
        RECT 420.975 -295.675 421.145 -294.815 ;
        RECT 419.245 -298.015 420.445 -297.845 ;
        RECT 410.975 -300.350 411.145 -298.630 ;
        RECT 411.955 -300.350 412.125 -298.630 ;
        RECT 414.020 -299.165 414.190 -298.625 ;
        RECT 415.000 -299.165 415.170 -298.625 ;
        RECT 413.430 -299.400 413.795 -299.335 ;
        RECT 412.930 -299.540 413.795 -299.400 ;
        RECT 412.820 -299.605 413.795 -299.540 ;
        RECT 412.820 -300.350 413.125 -299.605 ;
        RECT 413.430 -299.635 413.795 -299.605 ;
        RECT 415.980 -299.485 416.150 -298.625 ;
        RECT 410.060 -300.415 410.735 -300.385 ;
        RECT 409.960 -300.425 410.735 -300.415 ;
        RECT 407.320 -300.605 410.735 -300.425 ;
        RECT 410.975 -300.500 413.125 -300.350 ;
        RECT 410.975 -300.540 413.070 -300.500 ;
        RECT 414.020 -300.560 414.190 -299.780 ;
        RECT 414.510 -300.320 414.680 -299.780 ;
        RECT 415.000 -300.560 415.170 -299.780 ;
        RECT 415.490 -300.320 415.660 -299.780 ;
        RECT 415.980 -299.835 417.370 -299.485 ;
        RECT 408.235 -305.740 408.915 -300.605 ;
        RECT 409.960 -300.615 410.735 -300.605 ;
        RECT 410.060 -300.655 410.735 -300.615 ;
        RECT 409.195 -300.905 410.330 -300.895 ;
        RECT 412.385 -300.905 412.755 -300.775 ;
        RECT 409.195 -301.095 412.755 -300.905 ;
        RECT 413.320 -300.990 416.395 -300.560 ;
        RECT 410.325 -301.100 412.755 -301.095 ;
        RECT 410.325 -301.105 410.680 -301.100 ;
        RECT 412.385 -301.130 412.755 -301.100 ;
        RECT 410.485 -302.855 410.655 -301.315 ;
        RECT 410.975 -302.855 411.145 -301.315 ;
        RECT 411.465 -302.855 411.635 -301.315 ;
        RECT 411.955 -302.855 412.125 -301.315 ;
        RECT 412.445 -302.855 412.615 -301.315 ;
        RECT 410.970 -303.115 411.145 -302.855 ;
        RECT 414.540 -303.025 414.845 -300.990 ;
        RECT 416.990 -301.810 417.340 -299.835 ;
        RECT 418.210 -301.105 418.380 -298.185 ;
        RECT 419.245 -298.225 419.455 -298.015 ;
        RECT 418.190 -301.400 418.400 -301.105 ;
        RECT 419.265 -301.135 419.435 -298.225 ;
        RECT 419.755 -301.125 419.925 -298.185 ;
        RECT 420.235 -298.235 420.445 -298.015 ;
        RECT 419.250 -301.400 419.460 -301.135 ;
        RECT 418.190 -301.580 419.460 -301.400 ;
        RECT 419.735 -301.395 419.945 -301.125 ;
        RECT 420.245 -301.225 420.415 -298.235 ;
        RECT 421.305 -301.155 421.475 -298.185 ;
        RECT 419.735 -301.590 420.440 -301.395 ;
        RECT 420.225 -301.650 420.440 -301.590 ;
        RECT 419.015 -301.810 419.790 -301.760 ;
        RECT 416.990 -301.990 419.790 -301.810 ;
        RECT 416.990 -302.000 417.340 -301.990 ;
        RECT 419.015 -302.035 419.790 -301.990 ;
        RECT 420.225 -301.925 421.130 -301.650 ;
        RECT 420.225 -302.275 420.440 -301.925 ;
        RECT 417.665 -302.345 418.440 -302.300 ;
        RECT 417.480 -302.515 418.440 -302.345 ;
        RECT 417.665 -302.575 418.440 -302.515 ;
        RECT 418.670 -302.475 420.440 -302.275 ;
        RECT 421.300 -302.375 421.515 -301.155 ;
        RECT 422.485 -301.500 422.835 -294.815 ;
        RECT 423.825 -301.130 424.040 -291.255 ;
        RECT 425.460 -293.370 425.840 -289.850 ;
        RECT 426.970 -289.630 435.905 -289.440 ;
        RECT 426.970 -291.520 427.160 -289.630 ;
        RECT 433.005 -291.125 436.330 -290.985 ;
        RECT 433.005 -291.415 438.180 -291.125 ;
        RECT 426.855 -291.790 427.220 -291.520 ;
        RECT 433.005 -291.820 433.435 -291.415 ;
        RECT 434.305 -291.600 434.480 -291.415 ;
        RECT 435.930 -291.430 438.180 -291.415 ;
        RECT 428.745 -292.250 433.435 -291.820 ;
        RECT 427.985 -293.370 428.635 -293.240 ;
        RECT 425.460 -293.700 428.635 -293.370 ;
        RECT 429.445 -293.530 429.615 -292.250 ;
        RECT 429.935 -293.530 430.105 -292.490 ;
        RECT 430.425 -293.530 430.595 -292.250 ;
        RECT 430.915 -293.360 431.085 -292.490 ;
        RECT 433.820 -293.140 433.990 -291.600 ;
        RECT 434.310 -293.140 434.480 -291.600 ;
        RECT 434.800 -293.140 434.970 -291.600 ;
        RECT 435.290 -293.140 435.460 -291.600 ;
        RECT 435.780 -293.140 435.950 -291.600 ;
        RECT 433.660 -293.355 434.015 -293.350 ;
        RECT 435.720 -293.355 436.090 -293.325 ;
        RECT 433.660 -293.360 436.090 -293.355 ;
        RECT 430.915 -293.530 436.090 -293.360 ;
        RECT 437.875 -293.465 438.180 -291.430 ;
        RECT 430.920 -293.550 436.090 -293.530 ;
        RECT 430.920 -293.560 433.665 -293.550 ;
        RECT 428.855 -293.700 429.220 -293.670 ;
        RECT 435.720 -293.680 436.090 -293.550 ;
        RECT 425.460 -293.750 429.220 -293.700 ;
        RECT 427.985 -293.905 429.220 -293.750 ;
        RECT 433.395 -293.840 434.070 -293.800 ;
        RECT 433.295 -293.850 434.070 -293.840 ;
        RECT 427.985 -293.990 428.635 -293.905 ;
        RECT 428.855 -293.970 429.220 -293.905 ;
        RECT 428.120 -294.240 428.500 -293.990 ;
        RECT 432.260 -294.030 434.070 -293.850 ;
        RECT 436.655 -293.895 440.580 -293.465 ;
        RECT 433.295 -294.040 434.070 -294.030 ;
        RECT 433.395 -294.070 434.070 -294.040 ;
        RECT 434.310 -293.955 436.405 -293.915 ;
        RECT 434.310 -294.105 436.460 -293.955 ;
        RECT 429.445 -295.180 429.615 -294.140 ;
        RECT 430.425 -295.180 430.595 -294.140 ;
        RECT 431.405 -295.180 431.575 -294.140 ;
        RECT 434.310 -295.825 434.480 -294.105 ;
        RECT 435.290 -295.825 435.460 -294.105 ;
        RECT 436.155 -294.850 436.460 -294.105 ;
        RECT 437.355 -294.675 437.525 -293.895 ;
        RECT 437.845 -294.675 438.015 -294.135 ;
        RECT 438.335 -294.675 438.505 -293.895 ;
        RECT 438.825 -294.675 438.995 -294.135 ;
        RECT 436.765 -294.850 437.130 -294.820 ;
        RECT 436.155 -294.915 437.130 -294.850 ;
        RECT 436.265 -295.055 437.130 -294.915 ;
        RECT 436.765 -295.120 437.130 -295.055 ;
        RECT 439.315 -294.970 441.175 -294.620 ;
        RECT 437.355 -295.830 437.525 -295.290 ;
        RECT 438.335 -295.830 438.505 -295.290 ;
        RECT 439.315 -295.830 439.485 -294.970 ;
        RECT 437.585 -298.170 438.785 -298.000 ;
        RECT 429.315 -300.505 429.485 -298.785 ;
        RECT 430.295 -300.505 430.465 -298.785 ;
        RECT 432.360 -299.320 432.530 -298.780 ;
        RECT 433.340 -299.320 433.510 -298.780 ;
        RECT 431.770 -299.555 432.135 -299.490 ;
        RECT 431.270 -299.695 432.135 -299.555 ;
        RECT 431.160 -299.760 432.135 -299.695 ;
        RECT 431.160 -300.505 431.465 -299.760 ;
        RECT 431.770 -299.790 432.135 -299.760 ;
        RECT 434.320 -299.640 434.490 -298.780 ;
        RECT 428.400 -300.570 429.075 -300.540 ;
        RECT 428.300 -300.580 429.075 -300.570 ;
        RECT 426.230 -300.760 429.075 -300.580 ;
        RECT 429.315 -300.655 431.465 -300.505 ;
        RECT 429.315 -300.695 431.410 -300.655 ;
        RECT 432.360 -300.715 432.530 -299.935 ;
        RECT 432.850 -300.475 433.020 -299.935 ;
        RECT 433.340 -300.715 433.510 -299.935 ;
        RECT 433.830 -300.475 434.000 -299.935 ;
        RECT 434.320 -299.990 435.710 -299.640 ;
        RECT 423.825 -301.345 425.250 -301.130 ;
        RECT 422.430 -301.860 422.955 -301.500 ;
        RECT 425.035 -302.375 425.250 -301.345 ;
        RECT 412.595 -303.115 414.845 -303.025 ;
        RECT 410.385 -303.330 414.845 -303.115 ;
        RECT 410.385 -303.420 412.630 -303.330 ;
        RECT 414.540 -304.805 414.845 -303.330 ;
        RECT 418.210 -304.215 418.380 -302.745 ;
        RECT 418.670 -302.825 418.895 -302.475 ;
        RECT 420.630 -302.575 425.250 -302.375 ;
        RECT 420.870 -302.590 425.250 -302.575 ;
        RECT 418.175 -304.805 418.410 -304.215 ;
        RECT 418.700 -304.285 418.870 -302.825 ;
        RECT 419.190 -304.210 419.360 -302.745 ;
        RECT 420.400 -304.160 420.570 -302.745 ;
        RECT 420.870 -302.790 421.090 -302.590 ;
        RECT 419.155 -304.805 419.390 -304.210 ;
        RECT 420.365 -304.805 420.600 -304.160 ;
        RECT 420.890 -304.285 421.060 -302.790 ;
        RECT 414.540 -305.370 421.925 -304.805 ;
        RECT 426.230 -305.740 426.910 -300.760 ;
        RECT 428.300 -300.770 429.075 -300.760 ;
        RECT 428.400 -300.810 429.075 -300.770 ;
        RECT 427.535 -301.060 428.670 -301.050 ;
        RECT 430.725 -301.060 431.095 -300.930 ;
        RECT 427.535 -301.250 431.095 -301.060 ;
        RECT 431.660 -301.145 434.735 -300.715 ;
        RECT 428.665 -301.255 431.095 -301.250 ;
        RECT 428.665 -301.260 429.020 -301.255 ;
        RECT 430.725 -301.285 431.095 -301.255 ;
        RECT 428.825 -303.010 428.995 -301.470 ;
        RECT 429.315 -303.010 429.485 -301.470 ;
        RECT 429.805 -303.010 429.975 -301.470 ;
        RECT 430.295 -303.010 430.465 -301.470 ;
        RECT 430.785 -303.010 430.955 -301.470 ;
        RECT 429.310 -303.270 429.485 -303.010 ;
        RECT 432.880 -303.180 433.185 -301.145 ;
        RECT 435.330 -301.965 435.680 -299.990 ;
        RECT 436.550 -301.260 436.720 -298.340 ;
        RECT 437.585 -298.380 437.795 -298.170 ;
        RECT 436.530 -301.555 436.740 -301.260 ;
        RECT 437.605 -301.290 437.775 -298.380 ;
        RECT 438.095 -301.280 438.265 -298.340 ;
        RECT 438.575 -298.390 438.785 -298.170 ;
        RECT 437.590 -301.555 437.800 -301.290 ;
        RECT 436.530 -301.735 437.800 -301.555 ;
        RECT 438.075 -301.550 438.285 -301.280 ;
        RECT 438.585 -301.380 438.755 -298.390 ;
        RECT 439.645 -301.310 439.815 -298.340 ;
        RECT 438.075 -301.745 438.780 -301.550 ;
        RECT 438.565 -301.805 438.780 -301.745 ;
        RECT 437.355 -301.965 438.130 -301.915 ;
        RECT 435.330 -302.145 438.130 -301.965 ;
        RECT 435.330 -302.155 435.680 -302.145 ;
        RECT 437.355 -302.190 438.130 -302.145 ;
        RECT 438.565 -302.080 439.470 -301.805 ;
        RECT 438.565 -302.430 438.780 -302.080 ;
        RECT 436.005 -302.500 436.780 -302.455 ;
        RECT 435.820 -302.670 436.780 -302.500 ;
        RECT 436.005 -302.730 436.780 -302.670 ;
        RECT 437.010 -302.630 438.780 -302.430 ;
        RECT 439.640 -302.530 439.855 -301.310 ;
        RECT 440.825 -301.655 441.175 -294.970 ;
        RECT 440.770 -302.015 441.295 -301.655 ;
        RECT 443.915 -302.530 445.710 -301.780 ;
        RECT 430.935 -303.270 433.185 -303.180 ;
        RECT 428.725 -303.485 433.185 -303.270 ;
        RECT 428.725 -303.575 430.970 -303.485 ;
        RECT 432.880 -304.960 433.185 -303.485 ;
        RECT 436.550 -304.370 436.720 -302.900 ;
        RECT 437.010 -302.980 437.235 -302.630 ;
        RECT 438.970 -302.730 445.710 -302.530 ;
        RECT 439.210 -302.745 445.710 -302.730 ;
        RECT 436.515 -304.960 436.750 -304.370 ;
        RECT 437.040 -304.440 437.210 -302.980 ;
        RECT 437.530 -304.365 437.700 -302.900 ;
        RECT 438.740 -304.315 438.910 -302.900 ;
        RECT 439.210 -302.945 439.430 -302.745 ;
        RECT 437.495 -304.960 437.730 -304.365 ;
        RECT 438.705 -304.960 438.940 -304.315 ;
        RECT 439.230 -304.440 439.400 -302.945 ;
        RECT 443.915 -303.495 445.710 -302.745 ;
        RECT 432.880 -305.525 440.265 -304.960 ;
        RECT 408.235 -306.420 426.910 -305.740 ;
        RECT 405.030 -314.255 406.965 -312.875 ;
        RECT -119.230 -320.115 362.095 -319.435 ;
        RECT -119.230 -321.285 -118.550 -320.115 ;
        RECT 408.355 -321.285 409.035 -306.420 ;
        RECT -119.230 -321.965 409.035 -321.285 ;
        RECT -33.030 -324.485 91.690 -323.805 ;
        RECT -116.780 -325.670 59.060 -324.995 ;
      LAYER met1 ;
        RECT -62.330 605.045 -60.615 605.270 ;
        RECT -62.330 603.625 -8.150 605.045 ;
        RECT -62.330 603.475 -60.615 603.625 ;
        RECT -43.075 601.445 -42.765 601.510 ;
        RECT -60.850 600.685 -60.490 600.855 ;
        RECT -61.590 600.360 -60.490 600.685 ;
        RECT -63.255 598.760 -61.755 598.990 ;
        RECT -63.255 596.570 -61.755 596.800 ;
        RECT -61.590 595.585 -61.265 600.360 ;
        RECT -60.850 600.330 -60.490 600.360 ;
        RECT -43.075 600.350 -30.720 601.445 ;
        RECT -60.195 599.175 -57.195 599.405 ;
        RECT -53.865 599.075 -53.635 600.070 ;
        RECT -54.645 598.845 -53.635 599.075 ;
        RECT -53.865 598.585 -53.635 598.845 ;
        RECT -53.875 598.355 -52.990 598.585 ;
        RECT -60.195 598.115 -57.195 598.345 ;
        RECT -53.875 598.095 -53.635 598.355 ;
        RECT -54.645 597.865 -53.635 598.095 ;
        RECT -60.195 597.625 -57.195 597.855 ;
        RECT -53.875 597.605 -53.635 597.865 ;
        RECT -53.875 597.375 -52.990 597.605 ;
        RECT -60.195 597.135 -57.195 597.365 ;
        RECT -53.865 597.115 -53.635 597.375 ;
        RECT -54.645 596.885 -53.635 597.115 ;
        RECT -60.195 596.080 -57.195 596.310 ;
        RECT -51.955 595.310 -50.040 595.540 ;
        RECT -58.645 594.080 -58.415 595.075 ;
        RECT -54.640 594.820 -50.455 595.050 ;
        RECT -50.275 594.560 -50.040 595.310 ;
        RECT -51.955 594.330 -50.040 594.560 ;
        RECT -58.645 593.850 -57.635 594.080 ;
        RECT -58.645 593.590 -58.415 593.850 ;
        RECT -54.640 593.840 -53.140 594.070 ;
        RECT -59.290 593.360 -58.405 593.590 ;
        RECT -58.645 593.100 -58.405 593.360 ;
        RECT -52.910 593.270 -52.620 593.665 ;
        RECT -50.275 593.580 -50.040 594.330 ;
        RECT -45.545 593.975 -44.045 594.205 ;
        RECT -43.075 593.730 -42.765 600.350 ;
        RECT -51.955 593.350 -50.040 593.580 ;
        RECT -43.120 593.400 -42.705 593.730 ;
        RECT -40.565 593.485 -39.065 593.715 ;
        RECT -50.460 593.345 -50.040 593.350 ;
        RECT -58.645 592.870 -57.635 593.100 ;
        RECT -52.910 593.000 -52.075 593.270 ;
        RECT -52.910 592.870 -52.620 593.000 ;
        RECT -58.645 592.610 -58.405 592.870 ;
        RECT -59.290 592.380 -58.405 592.610 ;
        RECT -58.645 592.120 -58.415 592.380 ;
        RECT -58.645 591.890 -57.635 592.120 ;
        RECT -52.715 591.165 -52.485 592.160 ;
        RECT -52.345 591.900 -52.075 593.000 ;
        RECT -45.545 592.835 -43.045 593.065 ;
        RECT -45.545 592.345 -43.045 592.575 ;
        RECT -42.690 592.540 -42.000 592.810 ;
        RECT -52.345 591.630 -50.355 591.900 ;
        RECT -53.995 590.935 -52.485 591.165 ;
        RECT -52.715 590.675 -52.485 590.935 ;
        RECT -62.240 590.315 -60.325 590.545 ;
        RECT -52.725 590.445 -51.345 590.675 ;
        RECT -62.240 589.565 -62.005 590.315 ;
        RECT -52.725 590.185 -52.485 590.445 ;
        RECT -61.825 589.825 -57.640 590.055 ;
        RECT -53.995 589.955 -52.485 590.185 ;
        RECT -52.725 589.695 -52.485 589.955 ;
        RECT -62.240 589.335 -60.325 589.565 ;
        RECT -52.725 589.465 -51.345 589.695 ;
        RECT -62.240 588.585 -62.005 589.335 ;
        RECT -52.715 589.205 -52.485 589.465 ;
        RECT -59.140 588.845 -57.640 589.075 ;
        RECT -53.995 588.975 -52.485 589.205 ;
        RECT -62.240 588.355 -60.325 588.585 ;
        RECT -62.240 588.350 -61.820 588.355 ;
        RECT -52.825 588.065 -52.075 588.195 ;
        RECT -60.115 587.795 -52.075 588.065 ;
        RECT -60.115 587.080 -59.845 587.795 ;
        RECT -52.825 587.545 -52.075 587.795 ;
        RECT -50.625 586.840 -50.355 591.630 ;
        RECT -42.585 591.305 -42.365 592.540 ;
        RECT -41.565 592.345 -39.065 592.575 ;
        RECT -45.545 590.715 -43.045 590.945 ;
        RECT -42.615 590.615 -42.345 591.305 ;
        RECT -41.565 590.715 -39.065 590.945 ;
        RECT -45.545 590.090 -43.045 590.320 ;
        RECT -45.545 589.600 -43.045 589.830 ;
        RECT -45.545 587.740 -44.045 587.970 ;
        RECT -42.585 587.275 -42.365 590.615 ;
        RECT -41.565 590.065 -39.065 590.295 ;
        RECT -41.565 589.575 -39.065 589.805 ;
        RECT -41.565 589.085 -39.065 589.315 ;
        RECT -41.565 587.740 -39.065 587.970 ;
        RECT -50.655 586.355 -50.325 586.840 ;
        RECT -42.615 586.585 -42.345 587.275 ;
        RECT -44.300 586.235 -43.845 586.295 ;
        RECT -47.860 585.840 -43.845 586.235 ;
        RECT -50.120 583.735 -49.635 583.790 ;
        RECT -47.860 583.735 -47.465 585.840 ;
        RECT -44.300 585.780 -43.845 585.840 ;
        RECT -50.120 583.340 -47.465 583.735 ;
        RECT -50.120 583.210 -49.635 583.340 ;
        RECT -60.695 582.345 -60.335 582.515 ;
        RECT -43.430 582.385 -43.070 582.555 ;
        RECT -61.435 582.020 -60.335 582.345 ;
        RECT -63.100 580.420 -61.600 580.650 ;
        RECT -63.100 578.230 -61.600 578.460 ;
        RECT -61.435 577.245 -61.110 582.020 ;
        RECT -60.695 581.990 -60.335 582.020 ;
        RECT -44.170 582.060 -43.070 582.385 ;
        RECT -60.040 580.835 -57.040 581.065 ;
        RECT -53.710 580.735 -53.480 581.730 ;
        RECT -54.490 580.505 -53.480 580.735 ;
        RECT -53.710 580.245 -53.480 580.505 ;
        RECT -45.835 580.460 -44.335 580.690 ;
        RECT -53.720 580.015 -52.835 580.245 ;
        RECT -60.040 579.775 -57.040 580.005 ;
        RECT -53.720 579.755 -53.480 580.015 ;
        RECT -54.490 579.525 -53.480 579.755 ;
        RECT -60.040 579.285 -57.040 579.515 ;
        RECT -53.720 579.265 -53.480 579.525 ;
        RECT -53.720 579.035 -52.835 579.265 ;
        RECT -60.040 578.795 -57.040 579.025 ;
        RECT -53.710 578.775 -53.480 579.035 ;
        RECT -54.490 578.545 -53.480 578.775 ;
        RECT -45.835 578.270 -44.335 578.500 ;
        RECT -60.040 577.740 -57.040 577.970 ;
        RECT -44.170 577.285 -43.845 582.060 ;
        RECT -43.430 582.030 -43.070 582.060 ;
        RECT -42.775 580.875 -39.775 581.105 ;
        RECT -36.445 580.775 -36.215 581.770 ;
        RECT -37.225 580.545 -36.215 580.775 ;
        RECT -36.445 580.285 -36.215 580.545 ;
        RECT -36.455 580.055 -35.570 580.285 ;
        RECT -42.775 579.815 -39.775 580.045 ;
        RECT -36.455 579.795 -36.215 580.055 ;
        RECT -37.225 579.565 -36.215 579.795 ;
        RECT -42.775 579.325 -39.775 579.555 ;
        RECT -36.455 579.305 -36.215 579.565 ;
        RECT -36.455 579.075 -35.570 579.305 ;
        RECT -42.775 578.835 -39.775 579.065 ;
        RECT -36.445 578.815 -36.215 579.075 ;
        RECT -37.225 578.585 -36.215 578.815 ;
        RECT -42.775 577.780 -39.775 578.010 ;
        RECT -51.800 576.970 -49.885 577.200 ;
        RECT -34.535 577.010 -32.620 577.240 ;
        RECT -58.490 575.740 -58.260 576.735 ;
        RECT -54.485 576.480 -50.300 576.710 ;
        RECT -50.120 576.220 -49.885 576.970 ;
        RECT -51.800 575.990 -49.885 576.220 ;
        RECT -58.490 575.510 -57.480 575.740 ;
        RECT -58.490 575.250 -58.260 575.510 ;
        RECT -54.485 575.500 -52.985 575.730 ;
        RECT -59.135 575.020 -58.250 575.250 ;
        RECT -58.490 574.760 -58.250 575.020 ;
        RECT -52.755 574.930 -52.465 575.325 ;
        RECT -50.120 575.240 -49.885 575.990 ;
        RECT -41.225 575.780 -40.995 576.775 ;
        RECT -37.220 576.520 -33.035 576.750 ;
        RECT -32.855 576.260 -32.620 577.010 ;
        RECT -34.535 576.030 -32.620 576.260 ;
        RECT -41.225 575.550 -40.215 575.780 ;
        RECT -41.225 575.290 -40.995 575.550 ;
        RECT -37.220 575.540 -35.720 575.770 ;
        RECT -51.800 575.010 -49.885 575.240 ;
        RECT -41.870 575.060 -40.985 575.290 ;
        RECT -50.305 575.005 -49.885 575.010 ;
        RECT -58.490 574.530 -57.480 574.760 ;
        RECT -52.755 574.660 -51.920 574.930 ;
        RECT -52.755 574.530 -52.465 574.660 ;
        RECT -58.490 574.270 -58.250 574.530 ;
        RECT -59.135 574.040 -58.250 574.270 ;
        RECT -58.490 573.780 -58.260 574.040 ;
        RECT -58.490 573.550 -57.480 573.780 ;
        RECT -73.110 382.260 -71.685 573.200 ;
        RECT -86.585 380.835 -71.685 382.260 ;
        RECT -86.585 285.865 -85.160 380.835 ;
        RECT -73.505 375.780 -71.620 376.080 ;
        RECT -68.910 376.035 -68.005 573.200 ;
        RECT -52.560 572.825 -52.330 573.820 ;
        RECT -52.190 573.560 -51.920 574.660 ;
        RECT -41.225 574.800 -40.985 575.060 ;
        RECT -35.490 574.970 -35.200 575.365 ;
        RECT -32.855 575.280 -32.620 576.030 ;
        RECT -34.535 575.050 -32.620 575.280 ;
        RECT -33.040 575.045 -32.620 575.050 ;
        RECT -41.225 574.570 -40.215 574.800 ;
        RECT -35.490 574.700 -34.655 574.970 ;
        RECT -35.490 574.570 -35.200 574.700 ;
        RECT -41.225 574.310 -40.985 574.570 ;
        RECT -41.870 574.080 -40.985 574.310 ;
        RECT -41.225 573.820 -40.995 574.080 ;
        RECT -41.225 573.590 -40.215 573.820 ;
        RECT -52.190 573.290 -50.200 573.560 ;
        RECT -53.840 572.595 -52.330 572.825 ;
        RECT -52.560 572.335 -52.330 572.595 ;
        RECT -62.085 571.975 -60.170 572.205 ;
        RECT -52.570 572.105 -51.190 572.335 ;
        RECT -62.085 571.225 -61.850 571.975 ;
        RECT -52.570 571.845 -52.330 572.105 ;
        RECT -61.670 571.485 -57.485 571.715 ;
        RECT -53.840 571.615 -52.330 571.845 ;
        RECT -52.570 571.355 -52.330 571.615 ;
        RECT -62.085 570.995 -60.170 571.225 ;
        RECT -52.570 571.125 -51.190 571.355 ;
        RECT -62.085 570.245 -61.850 570.995 ;
        RECT -52.560 570.865 -52.330 571.125 ;
        RECT -58.985 570.505 -57.485 570.735 ;
        RECT -53.840 570.635 -52.330 570.865 ;
        RECT -62.085 570.015 -60.170 570.245 ;
        RECT -62.085 570.010 -61.665 570.015 ;
        RECT -52.670 569.725 -51.920 569.855 ;
        RECT -59.960 569.455 -51.920 569.725 ;
        RECT -59.960 568.740 -59.690 569.455 ;
        RECT -52.670 569.205 -51.920 569.455 ;
        RECT -50.470 567.745 -50.200 573.290 ;
        RECT -35.295 572.865 -35.065 573.860 ;
        RECT -34.925 573.600 -34.655 574.700 ;
        RECT -34.925 573.330 -32.935 573.600 ;
        RECT -36.575 572.635 -35.065 572.865 ;
        RECT -35.295 572.375 -35.065 572.635 ;
        RECT -44.820 572.015 -42.905 572.245 ;
        RECT -35.305 572.145 -33.925 572.375 ;
        RECT -44.820 571.265 -44.585 572.015 ;
        RECT -35.305 571.885 -35.065 572.145 ;
        RECT -44.405 571.525 -40.220 571.755 ;
        RECT -36.575 571.655 -35.065 571.885 ;
        RECT -35.305 571.395 -35.065 571.655 ;
        RECT -44.820 571.035 -42.905 571.265 ;
        RECT -35.305 571.165 -33.925 571.395 ;
        RECT -44.820 570.285 -44.585 571.035 ;
        RECT -35.295 570.905 -35.065 571.165 ;
        RECT -41.720 570.545 -40.220 570.775 ;
        RECT -36.575 570.675 -35.065 570.905 ;
        RECT -44.820 570.055 -42.905 570.285 ;
        RECT -44.820 570.050 -44.400 570.055 ;
        RECT -35.405 569.765 -34.655 569.895 ;
        RECT -42.695 569.495 -34.655 569.765 ;
        RECT -42.695 568.780 -42.425 569.495 ;
        RECT -35.405 569.245 -34.655 569.495 ;
        RECT -51.100 559.945 -50.005 567.745 ;
        RECT -33.205 567.590 -32.935 573.330 ;
        RECT -33.725 566.115 -32.360 567.590 ;
        RECT -31.815 559.945 -30.720 600.350 ;
        RECT -51.100 558.850 -30.720 559.945 ;
        RECT -62.455 555.970 -12.680 557.525 ;
        RECT -43.265 554.665 -42.955 554.690 ;
        RECT -61.040 553.865 -60.680 554.035 ;
        RECT -61.780 553.540 -60.680 553.865 ;
        RECT -63.445 551.940 -61.945 552.170 ;
        RECT -63.445 549.750 -61.945 549.980 ;
        RECT -61.780 548.765 -61.455 553.540 ;
        RECT -61.040 553.510 -60.680 553.540 ;
        RECT -60.385 552.355 -57.385 552.585 ;
        RECT -54.055 552.255 -53.825 553.250 ;
        RECT -54.835 552.025 -53.825 552.255 ;
        RECT -54.055 551.765 -53.825 552.025 ;
        RECT -43.265 553.130 -30.725 554.665 ;
        RECT -54.065 551.535 -53.180 551.765 ;
        RECT -60.385 551.295 -57.385 551.525 ;
        RECT -54.065 551.275 -53.825 551.535 ;
        RECT -54.835 551.045 -53.825 551.275 ;
        RECT -60.385 550.805 -57.385 551.035 ;
        RECT -54.065 550.785 -53.825 551.045 ;
        RECT -54.065 550.555 -53.180 550.785 ;
        RECT -60.385 550.315 -57.385 550.545 ;
        RECT -54.055 550.295 -53.825 550.555 ;
        RECT -54.835 550.065 -53.825 550.295 ;
        RECT -60.385 549.260 -57.385 549.490 ;
        RECT -52.145 548.490 -50.230 548.720 ;
        RECT -58.835 547.260 -58.605 548.255 ;
        RECT -54.830 548.000 -50.645 548.230 ;
        RECT -50.465 547.740 -50.230 548.490 ;
        RECT -52.145 547.510 -50.230 547.740 ;
        RECT -58.835 547.030 -57.825 547.260 ;
        RECT -58.835 546.770 -58.605 547.030 ;
        RECT -54.830 547.020 -53.330 547.250 ;
        RECT -59.480 546.540 -58.595 546.770 ;
        RECT -58.835 546.280 -58.595 546.540 ;
        RECT -53.100 546.450 -52.810 546.845 ;
        RECT -50.465 546.760 -50.230 547.510 ;
        RECT -45.735 547.155 -44.235 547.385 ;
        RECT -43.265 546.910 -42.955 553.130 ;
        RECT -52.145 546.530 -50.230 546.760 ;
        RECT -43.310 546.580 -42.895 546.910 ;
        RECT -40.755 546.665 -39.255 546.895 ;
        RECT -50.650 546.525 -50.230 546.530 ;
        RECT -58.835 546.050 -57.825 546.280 ;
        RECT -53.100 546.180 -52.265 546.450 ;
        RECT -53.100 546.050 -52.810 546.180 ;
        RECT -58.835 545.790 -58.595 546.050 ;
        RECT -59.480 545.560 -58.595 545.790 ;
        RECT -58.835 545.300 -58.605 545.560 ;
        RECT -58.835 545.070 -57.825 545.300 ;
        RECT -52.905 544.345 -52.675 545.340 ;
        RECT -52.535 545.080 -52.265 546.180 ;
        RECT -45.735 546.015 -43.235 546.245 ;
        RECT -45.735 545.525 -43.235 545.755 ;
        RECT -42.880 545.720 -42.190 545.990 ;
        RECT -52.535 544.810 -50.545 545.080 ;
        RECT -54.185 544.115 -52.675 544.345 ;
        RECT -52.905 543.855 -52.675 544.115 ;
        RECT -62.430 543.495 -60.515 543.725 ;
        RECT -52.915 543.625 -51.535 543.855 ;
        RECT -62.430 542.745 -62.195 543.495 ;
        RECT -52.915 543.365 -52.675 543.625 ;
        RECT -62.015 543.005 -57.830 543.235 ;
        RECT -54.185 543.135 -52.675 543.365 ;
        RECT -52.915 542.875 -52.675 543.135 ;
        RECT -62.430 542.515 -60.515 542.745 ;
        RECT -52.915 542.645 -51.535 542.875 ;
        RECT -62.430 541.765 -62.195 542.515 ;
        RECT -52.905 542.385 -52.675 542.645 ;
        RECT -59.330 542.025 -57.830 542.255 ;
        RECT -54.185 542.155 -52.675 542.385 ;
        RECT -62.430 541.535 -60.515 541.765 ;
        RECT -62.430 541.530 -62.010 541.535 ;
        RECT -53.015 541.245 -52.265 541.375 ;
        RECT -60.305 540.975 -52.265 541.245 ;
        RECT -60.305 540.260 -60.035 540.975 ;
        RECT -53.015 540.725 -52.265 540.975 ;
        RECT -50.815 540.020 -50.545 544.810 ;
        RECT -42.775 544.485 -42.555 545.720 ;
        RECT -41.755 545.525 -39.255 545.755 ;
        RECT -45.735 543.895 -43.235 544.125 ;
        RECT -42.805 543.795 -42.535 544.485 ;
        RECT -41.755 543.895 -39.255 544.125 ;
        RECT -45.735 543.270 -43.235 543.500 ;
        RECT -45.735 542.780 -43.235 543.010 ;
        RECT -45.735 540.920 -44.235 541.150 ;
        RECT -42.775 540.455 -42.555 543.795 ;
        RECT -41.755 543.245 -39.255 543.475 ;
        RECT -41.755 542.755 -39.255 542.985 ;
        RECT -41.755 542.265 -39.255 542.495 ;
        RECT -41.755 540.920 -39.255 541.150 ;
        RECT -50.845 539.535 -50.515 540.020 ;
        RECT -42.805 539.765 -42.535 540.455 ;
        RECT -44.490 539.415 -44.035 539.475 ;
        RECT -48.050 539.020 -44.035 539.415 ;
        RECT -50.310 536.915 -49.825 536.970 ;
        RECT -48.050 536.915 -47.655 539.020 ;
        RECT -44.490 538.960 -44.035 539.020 ;
        RECT -50.310 536.520 -47.655 536.915 ;
        RECT -50.310 536.390 -49.825 536.520 ;
        RECT -60.885 535.525 -60.525 535.695 ;
        RECT -43.620 535.565 -43.260 535.735 ;
        RECT -61.625 535.200 -60.525 535.525 ;
        RECT -63.290 533.600 -61.790 533.830 ;
        RECT -63.290 531.410 -61.790 531.640 ;
        RECT -61.625 530.425 -61.300 535.200 ;
        RECT -60.885 535.170 -60.525 535.200 ;
        RECT -44.360 535.240 -43.260 535.565 ;
        RECT -60.230 534.015 -57.230 534.245 ;
        RECT -53.900 533.915 -53.670 534.910 ;
        RECT -54.680 533.685 -53.670 533.915 ;
        RECT -53.900 533.425 -53.670 533.685 ;
        RECT -46.025 533.640 -44.525 533.870 ;
        RECT -53.910 533.195 -53.025 533.425 ;
        RECT -60.230 532.955 -57.230 533.185 ;
        RECT -53.910 532.935 -53.670 533.195 ;
        RECT -54.680 532.705 -53.670 532.935 ;
        RECT -60.230 532.465 -57.230 532.695 ;
        RECT -53.910 532.445 -53.670 532.705 ;
        RECT -53.910 532.215 -53.025 532.445 ;
        RECT -60.230 531.975 -57.230 532.205 ;
        RECT -53.900 531.955 -53.670 532.215 ;
        RECT -54.680 531.725 -53.670 531.955 ;
        RECT -46.025 531.450 -44.525 531.680 ;
        RECT -60.230 530.920 -57.230 531.150 ;
        RECT -44.360 530.465 -44.035 535.240 ;
        RECT -43.620 535.210 -43.260 535.240 ;
        RECT -42.965 534.055 -39.965 534.285 ;
        RECT -36.635 533.955 -36.405 534.950 ;
        RECT -37.415 533.725 -36.405 533.955 ;
        RECT -36.635 533.465 -36.405 533.725 ;
        RECT -36.645 533.235 -35.760 533.465 ;
        RECT -42.965 532.995 -39.965 533.225 ;
        RECT -36.645 532.975 -36.405 533.235 ;
        RECT -37.415 532.745 -36.405 532.975 ;
        RECT -42.965 532.505 -39.965 532.735 ;
        RECT -36.645 532.485 -36.405 532.745 ;
        RECT -36.645 532.255 -35.760 532.485 ;
        RECT -42.965 532.015 -39.965 532.245 ;
        RECT -36.635 531.995 -36.405 532.255 ;
        RECT -37.415 531.765 -36.405 531.995 ;
        RECT -42.965 530.960 -39.965 531.190 ;
        RECT -51.990 530.150 -50.075 530.380 ;
        RECT -34.725 530.190 -32.810 530.420 ;
        RECT -58.680 528.920 -58.450 529.915 ;
        RECT -54.675 529.660 -50.490 529.890 ;
        RECT -50.310 529.400 -50.075 530.150 ;
        RECT -51.990 529.170 -50.075 529.400 ;
        RECT -58.680 528.690 -57.670 528.920 ;
        RECT -58.680 528.430 -58.450 528.690 ;
        RECT -54.675 528.680 -53.175 528.910 ;
        RECT -59.325 528.200 -58.440 528.430 ;
        RECT -58.680 527.940 -58.440 528.200 ;
        RECT -52.945 528.110 -52.655 528.505 ;
        RECT -50.310 528.420 -50.075 529.170 ;
        RECT -41.415 528.960 -41.185 529.955 ;
        RECT -37.410 529.700 -33.225 529.930 ;
        RECT -33.045 529.440 -32.810 530.190 ;
        RECT -34.725 529.210 -32.810 529.440 ;
        RECT -41.415 528.730 -40.405 528.960 ;
        RECT -41.415 528.470 -41.185 528.730 ;
        RECT -37.410 528.720 -35.910 528.950 ;
        RECT -51.990 528.190 -50.075 528.420 ;
        RECT -42.060 528.240 -41.175 528.470 ;
        RECT -50.495 528.185 -50.075 528.190 ;
        RECT -58.680 527.710 -57.670 527.940 ;
        RECT -52.945 527.840 -52.110 528.110 ;
        RECT -52.945 527.710 -52.655 527.840 ;
        RECT -58.680 527.450 -58.440 527.710 ;
        RECT -59.325 527.220 -58.440 527.450 ;
        RECT -58.680 526.960 -58.450 527.220 ;
        RECT -58.680 526.730 -57.670 526.960 ;
        RECT -52.750 526.005 -52.520 527.000 ;
        RECT -52.380 526.740 -52.110 527.840 ;
        RECT -41.415 527.980 -41.175 528.240 ;
        RECT -35.680 528.150 -35.390 528.545 ;
        RECT -33.045 528.460 -32.810 529.210 ;
        RECT -34.725 528.230 -32.810 528.460 ;
        RECT -33.230 528.225 -32.810 528.230 ;
        RECT -41.415 527.750 -40.405 527.980 ;
        RECT -35.680 527.880 -34.845 528.150 ;
        RECT -35.680 527.750 -35.390 527.880 ;
        RECT -41.415 527.490 -41.175 527.750 ;
        RECT -42.060 527.260 -41.175 527.490 ;
        RECT -41.415 527.000 -41.185 527.260 ;
        RECT -41.415 526.770 -40.405 527.000 ;
        RECT -52.380 526.470 -50.390 526.740 ;
        RECT -54.030 525.775 -52.520 526.005 ;
        RECT -52.750 525.515 -52.520 525.775 ;
        RECT -62.275 525.155 -60.360 525.385 ;
        RECT -52.760 525.285 -51.380 525.515 ;
        RECT -62.275 524.405 -62.040 525.155 ;
        RECT -52.760 525.025 -52.520 525.285 ;
        RECT -61.860 524.665 -57.675 524.895 ;
        RECT -54.030 524.795 -52.520 525.025 ;
        RECT -52.760 524.535 -52.520 524.795 ;
        RECT -62.275 524.175 -60.360 524.405 ;
        RECT -52.760 524.305 -51.380 524.535 ;
        RECT -62.275 523.425 -62.040 524.175 ;
        RECT -52.750 524.045 -52.520 524.305 ;
        RECT -59.175 523.685 -57.675 523.915 ;
        RECT -54.030 523.815 -52.520 524.045 ;
        RECT -62.275 523.195 -60.360 523.425 ;
        RECT -62.275 523.190 -61.855 523.195 ;
        RECT -52.860 522.905 -52.110 523.035 ;
        RECT -60.150 522.635 -52.110 522.905 ;
        RECT -60.150 521.920 -59.880 522.635 ;
        RECT -52.860 522.385 -52.110 522.635 ;
        RECT -50.660 520.175 -50.390 526.470 ;
        RECT -35.485 526.045 -35.255 527.040 ;
        RECT -35.115 526.780 -34.845 527.880 ;
        RECT -35.115 526.510 -33.125 526.780 ;
        RECT -36.765 525.815 -35.255 526.045 ;
        RECT -35.485 525.555 -35.255 525.815 ;
        RECT -45.010 525.195 -43.095 525.425 ;
        RECT -35.495 525.325 -34.115 525.555 ;
        RECT -45.010 524.445 -44.775 525.195 ;
        RECT -35.495 525.065 -35.255 525.325 ;
        RECT -44.595 524.705 -40.410 524.935 ;
        RECT -36.765 524.835 -35.255 525.065 ;
        RECT -35.495 524.575 -35.255 524.835 ;
        RECT -45.010 524.215 -43.095 524.445 ;
        RECT -35.495 524.345 -34.115 524.575 ;
        RECT -45.010 523.465 -44.775 524.215 ;
        RECT -35.485 524.085 -35.255 524.345 ;
        RECT -41.910 523.725 -40.410 523.955 ;
        RECT -36.765 523.855 -35.255 524.085 ;
        RECT -45.010 523.235 -43.095 523.465 ;
        RECT -45.010 523.230 -44.590 523.235 ;
        RECT -35.595 522.945 -34.845 523.075 ;
        RECT -42.885 522.675 -34.845 522.945 ;
        RECT -42.885 521.960 -42.615 522.675 ;
        RECT -35.595 522.425 -34.845 522.675 ;
        RECT -33.395 521.180 -33.125 526.510 ;
        RECT -50.975 514.225 -49.475 520.175 ;
        RECT -33.870 519.840 -32.670 521.180 ;
        RECT -32.225 514.225 -30.725 553.130 ;
        RECT -50.975 512.725 -30.725 514.225 ;
        RECT -62.355 511.185 -60.835 511.395 ;
        RECT -33.850 511.185 -32.395 511.590 ;
        RECT -62.355 510.300 -15.600 511.185 ;
        RECT -62.355 510.090 -60.835 510.300 ;
        RECT -33.850 509.900 -32.395 510.300 ;
        RECT -43.350 508.715 -43.040 508.925 ;
        RECT -61.125 508.100 -60.765 508.270 ;
        RECT -61.865 507.775 -60.765 508.100 ;
        RECT -63.530 506.175 -62.030 506.405 ;
        RECT -63.530 503.985 -62.030 504.215 ;
        RECT -61.865 503.000 -61.540 507.775 ;
        RECT -61.125 507.745 -60.765 507.775 ;
        RECT -43.350 507.525 -30.995 508.715 ;
        RECT -60.470 506.590 -57.470 506.820 ;
        RECT -54.140 506.490 -53.910 507.485 ;
        RECT -54.920 506.260 -53.910 506.490 ;
        RECT -54.140 506.000 -53.910 506.260 ;
        RECT -54.150 505.770 -53.265 506.000 ;
        RECT -60.470 505.530 -57.470 505.760 ;
        RECT -54.150 505.510 -53.910 505.770 ;
        RECT -54.920 505.280 -53.910 505.510 ;
        RECT -60.470 505.040 -57.470 505.270 ;
        RECT -54.150 505.020 -53.910 505.280 ;
        RECT -54.150 504.790 -53.265 505.020 ;
        RECT -60.470 504.550 -57.470 504.780 ;
        RECT -54.140 504.530 -53.910 504.790 ;
        RECT -54.920 504.300 -53.910 504.530 ;
        RECT -60.470 503.495 -57.470 503.725 ;
        RECT -52.230 502.725 -50.315 502.955 ;
        RECT -58.920 501.495 -58.690 502.490 ;
        RECT -54.915 502.235 -50.730 502.465 ;
        RECT -50.550 501.975 -50.315 502.725 ;
        RECT -52.230 501.745 -50.315 501.975 ;
        RECT -58.920 501.265 -57.910 501.495 ;
        RECT -58.920 501.005 -58.690 501.265 ;
        RECT -54.915 501.255 -53.415 501.485 ;
        RECT -59.565 500.775 -58.680 501.005 ;
        RECT -58.920 500.515 -58.680 500.775 ;
        RECT -53.185 500.685 -52.895 501.080 ;
        RECT -50.550 500.995 -50.315 501.745 ;
        RECT -45.820 501.390 -44.320 501.620 ;
        RECT -43.350 501.145 -43.040 507.525 ;
        RECT -52.230 500.765 -50.315 500.995 ;
        RECT -43.395 500.815 -42.980 501.145 ;
        RECT -40.840 500.900 -39.340 501.130 ;
        RECT -50.735 500.760 -50.315 500.765 ;
        RECT -58.920 500.285 -57.910 500.515 ;
        RECT -53.185 500.415 -52.350 500.685 ;
        RECT -53.185 500.285 -52.895 500.415 ;
        RECT -58.920 500.025 -58.680 500.285 ;
        RECT -59.565 499.795 -58.680 500.025 ;
        RECT -58.920 499.535 -58.690 499.795 ;
        RECT -58.920 499.305 -57.910 499.535 ;
        RECT -52.990 498.580 -52.760 499.575 ;
        RECT -52.620 499.315 -52.350 500.415 ;
        RECT -45.820 500.250 -43.320 500.480 ;
        RECT -45.820 499.760 -43.320 499.990 ;
        RECT -42.965 499.955 -42.275 500.225 ;
        RECT -52.620 499.045 -50.630 499.315 ;
        RECT -54.270 498.350 -52.760 498.580 ;
        RECT -52.990 498.090 -52.760 498.350 ;
        RECT -62.515 497.730 -60.600 497.960 ;
        RECT -53.000 497.860 -51.620 498.090 ;
        RECT -62.515 496.980 -62.280 497.730 ;
        RECT -53.000 497.600 -52.760 497.860 ;
        RECT -62.100 497.240 -57.915 497.470 ;
        RECT -54.270 497.370 -52.760 497.600 ;
        RECT -53.000 497.110 -52.760 497.370 ;
        RECT -62.515 496.750 -60.600 496.980 ;
        RECT -53.000 496.880 -51.620 497.110 ;
        RECT -62.515 496.000 -62.280 496.750 ;
        RECT -52.990 496.620 -52.760 496.880 ;
        RECT -59.415 496.260 -57.915 496.490 ;
        RECT -54.270 496.390 -52.760 496.620 ;
        RECT -62.515 495.770 -60.600 496.000 ;
        RECT -62.515 495.765 -62.095 495.770 ;
        RECT -53.100 495.480 -52.350 495.610 ;
        RECT -60.390 495.210 -52.350 495.480 ;
        RECT -60.390 494.495 -60.120 495.210 ;
        RECT -53.100 494.960 -52.350 495.210 ;
        RECT -50.900 494.255 -50.630 499.045 ;
        RECT -42.860 498.720 -42.640 499.955 ;
        RECT -41.840 499.760 -39.340 499.990 ;
        RECT -45.820 498.130 -43.320 498.360 ;
        RECT -42.890 498.030 -42.620 498.720 ;
        RECT -41.840 498.130 -39.340 498.360 ;
        RECT -45.820 497.505 -43.320 497.735 ;
        RECT -45.820 497.015 -43.320 497.245 ;
        RECT -45.820 495.155 -44.320 495.385 ;
        RECT -42.860 494.690 -42.640 498.030 ;
        RECT -41.840 497.480 -39.340 497.710 ;
        RECT -41.840 496.990 -39.340 497.220 ;
        RECT -41.840 496.500 -39.340 496.730 ;
        RECT -41.840 495.155 -39.340 495.385 ;
        RECT -50.930 493.770 -50.600 494.255 ;
        RECT -42.890 494.000 -42.620 494.690 ;
        RECT -44.575 493.650 -44.120 493.710 ;
        RECT -48.135 493.255 -44.120 493.650 ;
        RECT -50.395 491.150 -49.910 491.205 ;
        RECT -48.135 491.150 -47.740 493.255 ;
        RECT -44.575 493.195 -44.120 493.255 ;
        RECT -50.395 490.755 -47.740 491.150 ;
        RECT -50.395 490.625 -49.910 490.755 ;
        RECT -60.970 489.760 -60.610 489.930 ;
        RECT -43.705 489.800 -43.345 489.970 ;
        RECT -61.710 489.435 -60.610 489.760 ;
        RECT -63.375 487.835 -61.875 488.065 ;
        RECT -63.375 485.645 -61.875 485.875 ;
        RECT -61.710 484.660 -61.385 489.435 ;
        RECT -60.970 489.405 -60.610 489.435 ;
        RECT -44.445 489.475 -43.345 489.800 ;
        RECT -60.315 488.250 -57.315 488.480 ;
        RECT -53.985 488.150 -53.755 489.145 ;
        RECT -54.765 487.920 -53.755 488.150 ;
        RECT -53.985 487.660 -53.755 487.920 ;
        RECT -46.110 487.875 -44.610 488.105 ;
        RECT -53.995 487.430 -53.110 487.660 ;
        RECT -60.315 487.190 -57.315 487.420 ;
        RECT -53.995 487.170 -53.755 487.430 ;
        RECT -54.765 486.940 -53.755 487.170 ;
        RECT -60.315 486.700 -57.315 486.930 ;
        RECT -53.995 486.680 -53.755 486.940 ;
        RECT -53.995 486.450 -53.110 486.680 ;
        RECT -60.315 486.210 -57.315 486.440 ;
        RECT -53.985 486.190 -53.755 486.450 ;
        RECT -54.765 485.960 -53.755 486.190 ;
        RECT -46.110 485.685 -44.610 485.915 ;
        RECT -60.315 485.155 -57.315 485.385 ;
        RECT -44.445 484.700 -44.120 489.475 ;
        RECT -43.705 489.445 -43.345 489.475 ;
        RECT -43.050 488.290 -40.050 488.520 ;
        RECT -36.720 488.190 -36.490 489.185 ;
        RECT -37.500 487.960 -36.490 488.190 ;
        RECT -36.720 487.700 -36.490 487.960 ;
        RECT -36.730 487.470 -35.845 487.700 ;
        RECT -43.050 487.230 -40.050 487.460 ;
        RECT -36.730 487.210 -36.490 487.470 ;
        RECT -37.500 486.980 -36.490 487.210 ;
        RECT -43.050 486.740 -40.050 486.970 ;
        RECT -36.730 486.720 -36.490 486.980 ;
        RECT -36.730 486.490 -35.845 486.720 ;
        RECT -43.050 486.250 -40.050 486.480 ;
        RECT -36.720 486.230 -36.490 486.490 ;
        RECT -37.500 486.000 -36.490 486.230 ;
        RECT -43.050 485.195 -40.050 485.425 ;
        RECT -52.075 484.385 -50.160 484.615 ;
        RECT -34.810 484.425 -32.895 484.655 ;
        RECT -58.765 483.155 -58.535 484.150 ;
        RECT -54.760 483.895 -50.575 484.125 ;
        RECT -50.395 483.635 -50.160 484.385 ;
        RECT -52.075 483.405 -50.160 483.635 ;
        RECT -58.765 482.925 -57.755 483.155 ;
        RECT -58.765 482.665 -58.535 482.925 ;
        RECT -54.760 482.915 -53.260 483.145 ;
        RECT -59.410 482.435 -58.525 482.665 ;
        RECT -58.765 482.175 -58.525 482.435 ;
        RECT -53.030 482.345 -52.740 482.740 ;
        RECT -50.395 482.655 -50.160 483.405 ;
        RECT -41.500 483.195 -41.270 484.190 ;
        RECT -37.495 483.935 -33.310 484.165 ;
        RECT -33.130 483.675 -32.895 484.425 ;
        RECT -34.810 483.445 -32.895 483.675 ;
        RECT -41.500 482.965 -40.490 483.195 ;
        RECT -41.500 482.705 -41.270 482.965 ;
        RECT -37.495 482.955 -35.995 483.185 ;
        RECT -52.075 482.425 -50.160 482.655 ;
        RECT -42.145 482.475 -41.260 482.705 ;
        RECT -50.580 482.420 -50.160 482.425 ;
        RECT -58.765 481.945 -57.755 482.175 ;
        RECT -53.030 482.075 -52.195 482.345 ;
        RECT -53.030 481.945 -52.740 482.075 ;
        RECT -58.765 481.685 -58.525 481.945 ;
        RECT -59.410 481.455 -58.525 481.685 ;
        RECT -58.765 481.195 -58.535 481.455 ;
        RECT -58.765 480.965 -57.755 481.195 ;
        RECT -52.835 480.240 -52.605 481.235 ;
        RECT -52.465 480.975 -52.195 482.075 ;
        RECT -41.500 482.215 -41.260 482.475 ;
        RECT -35.765 482.385 -35.475 482.780 ;
        RECT -33.130 482.695 -32.895 483.445 ;
        RECT -34.810 482.465 -32.895 482.695 ;
        RECT -33.315 482.460 -32.895 482.465 ;
        RECT -41.500 481.985 -40.490 482.215 ;
        RECT -35.765 482.115 -34.930 482.385 ;
        RECT -35.765 481.985 -35.475 482.115 ;
        RECT -41.500 481.725 -41.260 481.985 ;
        RECT -42.145 481.495 -41.260 481.725 ;
        RECT -41.500 481.235 -41.270 481.495 ;
        RECT -41.500 481.005 -40.490 481.235 ;
        RECT -52.465 480.705 -50.475 480.975 ;
        RECT -54.115 480.010 -52.605 480.240 ;
        RECT -52.835 479.750 -52.605 480.010 ;
        RECT -62.360 479.390 -60.445 479.620 ;
        RECT -52.845 479.520 -51.465 479.750 ;
        RECT -62.360 478.640 -62.125 479.390 ;
        RECT -52.845 479.260 -52.605 479.520 ;
        RECT -61.945 478.900 -57.760 479.130 ;
        RECT -54.115 479.030 -52.605 479.260 ;
        RECT -52.845 478.770 -52.605 479.030 ;
        RECT -62.360 478.410 -60.445 478.640 ;
        RECT -52.845 478.540 -51.465 478.770 ;
        RECT -62.360 477.660 -62.125 478.410 ;
        RECT -52.835 478.280 -52.605 478.540 ;
        RECT -59.260 477.920 -57.760 478.150 ;
        RECT -54.115 478.050 -52.605 478.280 ;
        RECT -62.360 477.430 -60.445 477.660 ;
        RECT -62.360 477.425 -61.940 477.430 ;
        RECT -52.945 477.140 -52.195 477.270 ;
        RECT -60.235 476.870 -52.195 477.140 ;
        RECT -60.235 476.155 -59.965 476.870 ;
        RECT -52.945 476.620 -52.195 476.870 ;
        RECT -50.745 474.475 -50.475 480.705 ;
        RECT -35.570 480.280 -35.340 481.275 ;
        RECT -35.200 481.015 -34.930 482.115 ;
        RECT -35.200 480.745 -33.210 481.015 ;
        RECT -36.850 480.050 -35.340 480.280 ;
        RECT -35.570 479.790 -35.340 480.050 ;
        RECT -45.095 479.430 -43.180 479.660 ;
        RECT -35.580 479.560 -34.200 479.790 ;
        RECT -45.095 478.680 -44.860 479.430 ;
        RECT -35.580 479.300 -35.340 479.560 ;
        RECT -44.680 478.940 -40.495 479.170 ;
        RECT -36.850 479.070 -35.340 479.300 ;
        RECT -35.580 478.810 -35.340 479.070 ;
        RECT -45.095 478.450 -43.180 478.680 ;
        RECT -35.580 478.580 -34.200 478.810 ;
        RECT -45.095 477.700 -44.860 478.450 ;
        RECT -35.570 478.320 -35.340 478.580 ;
        RECT -41.995 477.960 -40.495 478.190 ;
        RECT -36.850 478.090 -35.340 478.320 ;
        RECT -45.095 477.470 -43.180 477.700 ;
        RECT -45.095 477.465 -44.675 477.470 ;
        RECT -35.680 477.180 -34.930 477.310 ;
        RECT -42.970 476.910 -34.930 477.180 ;
        RECT -42.970 476.195 -42.700 476.910 ;
        RECT -35.680 476.660 -34.930 476.910 ;
        RECT -33.480 475.275 -33.210 480.745 ;
        RECT -50.995 469.985 -49.805 474.475 ;
        RECT -33.855 474.025 -32.710 475.275 ;
        RECT -32.185 469.985 -30.995 507.525 ;
        RECT -50.995 468.795 -30.995 469.985 ;
        RECT -62.620 467.640 -61.125 467.725 ;
        RECT -33.940 467.640 -32.370 467.900 ;
        RECT -62.620 466.535 -18.175 467.640 ;
        RECT -62.620 466.265 -61.125 466.535 ;
        RECT -33.940 466.020 -32.370 466.535 ;
        RECT -43.680 464.780 -43.370 465.155 ;
        RECT -61.455 464.330 -61.095 464.500 ;
        RECT -62.195 464.005 -61.095 464.330 ;
        RECT -63.860 462.405 -62.360 462.635 ;
        RECT -63.860 460.215 -62.360 460.445 ;
        RECT -62.195 459.230 -61.870 464.005 ;
        RECT -61.455 463.975 -61.095 464.005 ;
        RECT -60.800 462.820 -57.800 463.050 ;
        RECT -54.470 462.720 -54.240 463.715 ;
        RECT -55.250 462.490 -54.240 462.720 ;
        RECT -54.470 462.230 -54.240 462.490 ;
        RECT -43.680 463.485 -30.790 464.780 ;
        RECT -54.480 462.000 -53.595 462.230 ;
        RECT -60.800 461.760 -57.800 461.990 ;
        RECT -54.480 461.740 -54.240 462.000 ;
        RECT -55.250 461.510 -54.240 461.740 ;
        RECT -60.800 461.270 -57.800 461.500 ;
        RECT -54.480 461.250 -54.240 461.510 ;
        RECT -54.480 461.020 -53.595 461.250 ;
        RECT -60.800 460.780 -57.800 461.010 ;
        RECT -54.470 460.760 -54.240 461.020 ;
        RECT -55.250 460.530 -54.240 460.760 ;
        RECT -60.800 459.725 -57.800 459.955 ;
        RECT -52.560 458.955 -50.645 459.185 ;
        RECT -59.250 457.725 -59.020 458.720 ;
        RECT -55.245 458.465 -51.060 458.695 ;
        RECT -50.880 458.205 -50.645 458.955 ;
        RECT -52.560 457.975 -50.645 458.205 ;
        RECT -59.250 457.495 -58.240 457.725 ;
        RECT -59.250 457.235 -59.020 457.495 ;
        RECT -55.245 457.485 -53.745 457.715 ;
        RECT -59.895 457.005 -59.010 457.235 ;
        RECT -59.250 456.745 -59.010 457.005 ;
        RECT -53.515 456.915 -53.225 457.310 ;
        RECT -50.880 457.225 -50.645 457.975 ;
        RECT -46.150 457.620 -44.650 457.850 ;
        RECT -43.680 457.375 -43.370 463.485 ;
        RECT -52.560 456.995 -50.645 457.225 ;
        RECT -43.725 457.045 -43.310 457.375 ;
        RECT -41.170 457.130 -39.670 457.360 ;
        RECT -51.065 456.990 -50.645 456.995 ;
        RECT -59.250 456.515 -58.240 456.745 ;
        RECT -53.515 456.645 -52.680 456.915 ;
        RECT -53.515 456.515 -53.225 456.645 ;
        RECT -59.250 456.255 -59.010 456.515 ;
        RECT -59.895 456.025 -59.010 456.255 ;
        RECT -59.250 455.765 -59.020 456.025 ;
        RECT -59.250 455.535 -58.240 455.765 ;
        RECT -53.320 454.810 -53.090 455.805 ;
        RECT -52.950 455.545 -52.680 456.645 ;
        RECT -46.150 456.480 -43.650 456.710 ;
        RECT -46.150 455.990 -43.650 456.220 ;
        RECT -43.295 456.185 -42.605 456.455 ;
        RECT -52.950 455.275 -50.960 455.545 ;
        RECT -54.600 454.580 -53.090 454.810 ;
        RECT -53.320 454.320 -53.090 454.580 ;
        RECT -62.845 453.960 -60.930 454.190 ;
        RECT -53.330 454.090 -51.950 454.320 ;
        RECT -62.845 453.210 -62.610 453.960 ;
        RECT -53.330 453.830 -53.090 454.090 ;
        RECT -62.430 453.470 -58.245 453.700 ;
        RECT -54.600 453.600 -53.090 453.830 ;
        RECT -53.330 453.340 -53.090 453.600 ;
        RECT -62.845 452.980 -60.930 453.210 ;
        RECT -53.330 453.110 -51.950 453.340 ;
        RECT -62.845 452.230 -62.610 452.980 ;
        RECT -53.320 452.850 -53.090 453.110 ;
        RECT -59.745 452.490 -58.245 452.720 ;
        RECT -54.600 452.620 -53.090 452.850 ;
        RECT -62.845 452.000 -60.930 452.230 ;
        RECT -62.845 451.995 -62.425 452.000 ;
        RECT -53.430 451.710 -52.680 451.840 ;
        RECT -60.720 451.440 -52.680 451.710 ;
        RECT -60.720 450.725 -60.450 451.440 ;
        RECT -53.430 451.190 -52.680 451.440 ;
        RECT -51.230 450.485 -50.960 455.275 ;
        RECT -43.190 454.950 -42.970 456.185 ;
        RECT -42.170 455.990 -39.670 456.220 ;
        RECT -46.150 454.360 -43.650 454.590 ;
        RECT -43.220 454.260 -42.950 454.950 ;
        RECT -42.170 454.360 -39.670 454.590 ;
        RECT -46.150 453.735 -43.650 453.965 ;
        RECT -46.150 453.245 -43.650 453.475 ;
        RECT -46.150 451.385 -44.650 451.615 ;
        RECT -43.190 450.920 -42.970 454.260 ;
        RECT -42.170 453.710 -39.670 453.940 ;
        RECT -42.170 453.220 -39.670 453.450 ;
        RECT -42.170 452.730 -39.670 452.960 ;
        RECT -42.170 451.385 -39.670 451.615 ;
        RECT -51.260 450.000 -50.930 450.485 ;
        RECT -43.220 450.230 -42.950 450.920 ;
        RECT -44.905 449.880 -44.450 449.940 ;
        RECT -48.465 449.485 -44.450 449.880 ;
        RECT -50.725 447.380 -50.240 447.435 ;
        RECT -48.465 447.380 -48.070 449.485 ;
        RECT -44.905 449.425 -44.450 449.485 ;
        RECT -50.725 446.985 -48.070 447.380 ;
        RECT -50.725 446.855 -50.240 446.985 ;
        RECT -61.300 445.990 -60.940 446.160 ;
        RECT -44.035 446.030 -43.675 446.200 ;
        RECT -62.040 445.665 -60.940 445.990 ;
        RECT -63.705 444.065 -62.205 444.295 ;
        RECT -63.705 441.875 -62.205 442.105 ;
        RECT -62.040 440.890 -61.715 445.665 ;
        RECT -61.300 445.635 -60.940 445.665 ;
        RECT -44.775 445.705 -43.675 446.030 ;
        RECT -60.645 444.480 -57.645 444.710 ;
        RECT -54.315 444.380 -54.085 445.375 ;
        RECT -55.095 444.150 -54.085 444.380 ;
        RECT -54.315 443.890 -54.085 444.150 ;
        RECT -46.440 444.105 -44.940 444.335 ;
        RECT -54.325 443.660 -53.440 443.890 ;
        RECT -60.645 443.420 -57.645 443.650 ;
        RECT -54.325 443.400 -54.085 443.660 ;
        RECT -55.095 443.170 -54.085 443.400 ;
        RECT -60.645 442.930 -57.645 443.160 ;
        RECT -54.325 442.910 -54.085 443.170 ;
        RECT -54.325 442.680 -53.440 442.910 ;
        RECT -60.645 442.440 -57.645 442.670 ;
        RECT -54.315 442.420 -54.085 442.680 ;
        RECT -55.095 442.190 -54.085 442.420 ;
        RECT -46.440 441.915 -44.940 442.145 ;
        RECT -60.645 441.385 -57.645 441.615 ;
        RECT -44.775 440.930 -44.450 445.705 ;
        RECT -44.035 445.675 -43.675 445.705 ;
        RECT -43.380 444.520 -40.380 444.750 ;
        RECT -37.050 444.420 -36.820 445.415 ;
        RECT -37.830 444.190 -36.820 444.420 ;
        RECT -37.050 443.930 -36.820 444.190 ;
        RECT -37.060 443.700 -36.175 443.930 ;
        RECT -43.380 443.460 -40.380 443.690 ;
        RECT -37.060 443.440 -36.820 443.700 ;
        RECT -37.830 443.210 -36.820 443.440 ;
        RECT -43.380 442.970 -40.380 443.200 ;
        RECT -37.060 442.950 -36.820 443.210 ;
        RECT -37.060 442.720 -36.175 442.950 ;
        RECT -43.380 442.480 -40.380 442.710 ;
        RECT -37.050 442.460 -36.820 442.720 ;
        RECT -37.830 442.230 -36.820 442.460 ;
        RECT -43.380 441.425 -40.380 441.655 ;
        RECT -52.405 440.615 -50.490 440.845 ;
        RECT -35.140 440.655 -33.225 440.885 ;
        RECT -59.095 439.385 -58.865 440.380 ;
        RECT -55.090 440.125 -50.905 440.355 ;
        RECT -50.725 439.865 -50.490 440.615 ;
        RECT -52.405 439.635 -50.490 439.865 ;
        RECT -59.095 439.155 -58.085 439.385 ;
        RECT -59.095 438.895 -58.865 439.155 ;
        RECT -55.090 439.145 -53.590 439.375 ;
        RECT -59.740 438.665 -58.855 438.895 ;
        RECT -59.095 438.405 -58.855 438.665 ;
        RECT -53.360 438.575 -53.070 438.970 ;
        RECT -50.725 438.885 -50.490 439.635 ;
        RECT -41.830 439.425 -41.600 440.420 ;
        RECT -37.825 440.165 -33.640 440.395 ;
        RECT -33.460 439.905 -33.225 440.655 ;
        RECT -35.140 439.675 -33.225 439.905 ;
        RECT -41.830 439.195 -40.820 439.425 ;
        RECT -41.830 438.935 -41.600 439.195 ;
        RECT -37.825 439.185 -36.325 439.415 ;
        RECT -52.405 438.655 -50.490 438.885 ;
        RECT -42.475 438.705 -41.590 438.935 ;
        RECT -50.910 438.650 -50.490 438.655 ;
        RECT -59.095 438.175 -58.085 438.405 ;
        RECT -53.360 438.305 -52.525 438.575 ;
        RECT -53.360 438.175 -53.070 438.305 ;
        RECT -59.095 437.915 -58.855 438.175 ;
        RECT -59.740 437.685 -58.855 437.915 ;
        RECT -59.095 437.425 -58.865 437.685 ;
        RECT -59.095 437.195 -58.085 437.425 ;
        RECT -53.165 436.470 -52.935 437.465 ;
        RECT -52.795 437.205 -52.525 438.305 ;
        RECT -41.830 438.445 -41.590 438.705 ;
        RECT -36.095 438.615 -35.805 439.010 ;
        RECT -33.460 438.925 -33.225 439.675 ;
        RECT -35.140 438.695 -33.225 438.925 ;
        RECT -33.645 438.690 -33.225 438.695 ;
        RECT -41.830 438.215 -40.820 438.445 ;
        RECT -36.095 438.345 -35.260 438.615 ;
        RECT -36.095 438.215 -35.805 438.345 ;
        RECT -41.830 437.955 -41.590 438.215 ;
        RECT -42.475 437.725 -41.590 437.955 ;
        RECT -41.830 437.465 -41.600 437.725 ;
        RECT -41.830 437.235 -40.820 437.465 ;
        RECT -52.795 436.935 -50.805 437.205 ;
        RECT -54.445 436.240 -52.935 436.470 ;
        RECT -53.165 435.980 -52.935 436.240 ;
        RECT -62.690 435.620 -60.775 435.850 ;
        RECT -53.175 435.750 -51.795 435.980 ;
        RECT -62.690 434.870 -62.455 435.620 ;
        RECT -53.175 435.490 -52.935 435.750 ;
        RECT -62.275 435.130 -58.090 435.360 ;
        RECT -54.445 435.260 -52.935 435.490 ;
        RECT -53.175 435.000 -52.935 435.260 ;
        RECT -62.690 434.640 -60.775 434.870 ;
        RECT -53.175 434.770 -51.795 435.000 ;
        RECT -62.690 433.890 -62.455 434.640 ;
        RECT -53.165 434.510 -52.935 434.770 ;
        RECT -59.590 434.150 -58.090 434.380 ;
        RECT -54.445 434.280 -52.935 434.510 ;
        RECT -62.690 433.660 -60.775 433.890 ;
        RECT -62.690 433.655 -62.270 433.660 ;
        RECT -53.275 433.370 -52.525 433.500 ;
        RECT -60.565 433.100 -52.525 433.370 ;
        RECT -60.565 432.385 -60.295 433.100 ;
        RECT -53.275 432.850 -52.525 433.100 ;
        RECT -51.075 430.890 -50.805 436.935 ;
        RECT -35.900 436.510 -35.670 437.505 ;
        RECT -35.530 437.245 -35.260 438.345 ;
        RECT -35.530 436.975 -33.540 437.245 ;
        RECT -37.180 436.280 -35.670 436.510 ;
        RECT -35.900 436.020 -35.670 436.280 ;
        RECT -45.425 435.660 -43.510 435.890 ;
        RECT -35.910 435.790 -34.530 436.020 ;
        RECT -45.425 434.910 -45.190 435.660 ;
        RECT -35.910 435.530 -35.670 435.790 ;
        RECT -45.010 435.170 -40.825 435.400 ;
        RECT -37.180 435.300 -35.670 435.530 ;
        RECT -35.910 435.040 -35.670 435.300 ;
        RECT -45.425 434.680 -43.510 434.910 ;
        RECT -35.910 434.810 -34.530 435.040 ;
        RECT -45.425 433.930 -45.190 434.680 ;
        RECT -35.900 434.550 -35.670 434.810 ;
        RECT -42.325 434.190 -40.825 434.420 ;
        RECT -37.180 434.320 -35.670 434.550 ;
        RECT -45.425 433.700 -43.510 433.930 ;
        RECT -45.425 433.695 -45.005 433.700 ;
        RECT -36.010 433.410 -35.260 433.540 ;
        RECT -43.300 433.140 -35.260 433.410 ;
        RECT -43.300 432.425 -43.030 433.140 ;
        RECT -36.010 432.890 -35.260 433.140 ;
        RECT -51.400 426.145 -50.105 430.890 ;
        RECT -33.810 430.060 -33.540 436.975 ;
        RECT -34.160 428.830 -33.060 430.060 ;
        RECT -32.085 426.145 -30.790 463.485 ;
        RECT -51.400 424.850 -30.790 426.145 ;
        RECT -62.935 421.695 -60.435 421.945 ;
        RECT -62.935 420.565 -20.935 421.695 ;
        RECT -62.935 420.455 -60.435 420.565 ;
        RECT -61.625 418.340 -61.265 418.510 ;
        RECT -62.365 418.015 -61.265 418.340 ;
        RECT -64.030 416.415 -62.530 416.645 ;
        RECT -64.030 414.225 -62.530 414.455 ;
        RECT -62.365 413.240 -62.040 418.015 ;
        RECT -61.625 417.985 -61.265 418.015 ;
        RECT -43.850 418.260 -43.540 419.165 ;
        RECT -60.970 416.830 -57.970 417.060 ;
        RECT -54.640 416.730 -54.410 417.725 ;
        RECT -55.420 416.500 -54.410 416.730 ;
        RECT -54.640 416.240 -54.410 416.500 ;
        RECT -43.850 417.250 -30.750 418.260 ;
        RECT -54.650 416.010 -53.765 416.240 ;
        RECT -60.970 415.770 -57.970 416.000 ;
        RECT -54.650 415.750 -54.410 416.010 ;
        RECT -55.420 415.520 -54.410 415.750 ;
        RECT -60.970 415.280 -57.970 415.510 ;
        RECT -54.650 415.260 -54.410 415.520 ;
        RECT -54.650 415.030 -53.765 415.260 ;
        RECT -60.970 414.790 -57.970 415.020 ;
        RECT -54.640 414.770 -54.410 415.030 ;
        RECT -55.420 414.540 -54.410 414.770 ;
        RECT -60.970 413.735 -57.970 413.965 ;
        RECT -52.730 412.965 -50.815 413.195 ;
        RECT -59.420 411.735 -59.190 412.730 ;
        RECT -55.415 412.475 -51.230 412.705 ;
        RECT -51.050 412.215 -50.815 412.965 ;
        RECT -52.730 411.985 -50.815 412.215 ;
        RECT -59.420 411.505 -58.410 411.735 ;
        RECT -59.420 411.245 -59.190 411.505 ;
        RECT -55.415 411.495 -53.915 411.725 ;
        RECT -60.065 411.015 -59.180 411.245 ;
        RECT -59.420 410.755 -59.180 411.015 ;
        RECT -53.685 410.925 -53.395 411.320 ;
        RECT -51.050 411.235 -50.815 411.985 ;
        RECT -46.320 411.630 -44.820 411.860 ;
        RECT -43.850 411.385 -43.540 417.250 ;
        RECT -52.730 411.005 -50.815 411.235 ;
        RECT -43.895 411.055 -43.480 411.385 ;
        RECT -41.340 411.140 -39.840 411.370 ;
        RECT -51.235 411.000 -50.815 411.005 ;
        RECT -59.420 410.525 -58.410 410.755 ;
        RECT -53.685 410.655 -52.850 410.925 ;
        RECT -53.685 410.525 -53.395 410.655 ;
        RECT -59.420 410.265 -59.180 410.525 ;
        RECT -60.065 410.035 -59.180 410.265 ;
        RECT -59.420 409.775 -59.190 410.035 ;
        RECT -59.420 409.545 -58.410 409.775 ;
        RECT -53.490 408.820 -53.260 409.815 ;
        RECT -53.120 409.555 -52.850 410.655 ;
        RECT -46.320 410.490 -43.820 410.720 ;
        RECT -46.320 410.000 -43.820 410.230 ;
        RECT -43.465 410.195 -42.775 410.465 ;
        RECT -53.120 409.285 -51.130 409.555 ;
        RECT -54.770 408.590 -53.260 408.820 ;
        RECT -53.490 408.330 -53.260 408.590 ;
        RECT -63.015 407.970 -61.100 408.200 ;
        RECT -53.500 408.100 -52.120 408.330 ;
        RECT -63.015 407.220 -62.780 407.970 ;
        RECT -53.500 407.840 -53.260 408.100 ;
        RECT -62.600 407.480 -58.415 407.710 ;
        RECT -54.770 407.610 -53.260 407.840 ;
        RECT -53.500 407.350 -53.260 407.610 ;
        RECT -63.015 406.990 -61.100 407.220 ;
        RECT -53.500 407.120 -52.120 407.350 ;
        RECT -63.015 406.240 -62.780 406.990 ;
        RECT -53.490 406.860 -53.260 407.120 ;
        RECT -59.915 406.500 -58.415 406.730 ;
        RECT -54.770 406.630 -53.260 406.860 ;
        RECT -63.015 406.010 -61.100 406.240 ;
        RECT -63.015 406.005 -62.595 406.010 ;
        RECT -53.600 405.720 -52.850 405.850 ;
        RECT -60.890 405.450 -52.850 405.720 ;
        RECT -60.890 404.735 -60.620 405.450 ;
        RECT -53.600 405.200 -52.850 405.450 ;
        RECT -51.400 404.495 -51.130 409.285 ;
        RECT -43.360 408.960 -43.140 410.195 ;
        RECT -42.340 410.000 -39.840 410.230 ;
        RECT -46.320 408.370 -43.820 408.600 ;
        RECT -43.390 408.270 -43.120 408.960 ;
        RECT -42.340 408.370 -39.840 408.600 ;
        RECT -46.320 407.745 -43.820 407.975 ;
        RECT -46.320 407.255 -43.820 407.485 ;
        RECT -46.320 405.395 -44.820 405.625 ;
        RECT -43.360 404.930 -43.140 408.270 ;
        RECT -42.340 407.720 -39.840 407.950 ;
        RECT -42.340 407.230 -39.840 407.460 ;
        RECT -42.340 406.740 -39.840 406.970 ;
        RECT -42.340 405.395 -39.840 405.625 ;
        RECT -51.430 404.010 -51.100 404.495 ;
        RECT -43.390 404.240 -43.120 404.930 ;
        RECT -45.075 403.890 -44.620 403.950 ;
        RECT -48.635 403.495 -44.620 403.890 ;
        RECT -50.895 401.390 -50.410 401.445 ;
        RECT -48.635 401.390 -48.240 403.495 ;
        RECT -45.075 403.435 -44.620 403.495 ;
        RECT -50.895 400.995 -48.240 401.390 ;
        RECT -50.895 400.865 -50.410 400.995 ;
        RECT -61.470 400.000 -61.110 400.170 ;
        RECT -44.205 400.040 -43.845 400.210 ;
        RECT -62.210 399.675 -61.110 400.000 ;
        RECT -63.875 398.075 -62.375 398.305 ;
        RECT -63.875 395.885 -62.375 396.115 ;
        RECT -62.210 394.900 -61.885 399.675 ;
        RECT -61.470 399.645 -61.110 399.675 ;
        RECT -44.945 399.715 -43.845 400.040 ;
        RECT -60.815 398.490 -57.815 398.720 ;
        RECT -54.485 398.390 -54.255 399.385 ;
        RECT -55.265 398.160 -54.255 398.390 ;
        RECT -54.485 397.900 -54.255 398.160 ;
        RECT -46.610 398.115 -45.110 398.345 ;
        RECT -54.495 397.670 -53.610 397.900 ;
        RECT -60.815 397.430 -57.815 397.660 ;
        RECT -54.495 397.410 -54.255 397.670 ;
        RECT -55.265 397.180 -54.255 397.410 ;
        RECT -60.815 396.940 -57.815 397.170 ;
        RECT -54.495 396.920 -54.255 397.180 ;
        RECT -54.495 396.690 -53.610 396.920 ;
        RECT -60.815 396.450 -57.815 396.680 ;
        RECT -54.485 396.430 -54.255 396.690 ;
        RECT -55.265 396.200 -54.255 396.430 ;
        RECT -46.610 395.925 -45.110 396.155 ;
        RECT -60.815 395.395 -57.815 395.625 ;
        RECT -44.945 394.940 -44.620 399.715 ;
        RECT -44.205 399.685 -43.845 399.715 ;
        RECT -43.550 398.530 -40.550 398.760 ;
        RECT -37.220 398.430 -36.990 399.425 ;
        RECT -38.000 398.200 -36.990 398.430 ;
        RECT -37.220 397.940 -36.990 398.200 ;
        RECT -37.230 397.710 -36.345 397.940 ;
        RECT -43.550 397.470 -40.550 397.700 ;
        RECT -37.230 397.450 -36.990 397.710 ;
        RECT -38.000 397.220 -36.990 397.450 ;
        RECT -43.550 396.980 -40.550 397.210 ;
        RECT -37.230 396.960 -36.990 397.220 ;
        RECT -37.230 396.730 -36.345 396.960 ;
        RECT -43.550 396.490 -40.550 396.720 ;
        RECT -37.220 396.470 -36.990 396.730 ;
        RECT -38.000 396.240 -36.990 396.470 ;
        RECT -43.550 395.435 -40.550 395.665 ;
        RECT -52.575 394.625 -50.660 394.855 ;
        RECT -35.310 394.665 -33.395 394.895 ;
        RECT -59.265 393.395 -59.035 394.390 ;
        RECT -55.260 394.135 -51.075 394.365 ;
        RECT -50.895 393.875 -50.660 394.625 ;
        RECT -52.575 393.645 -50.660 393.875 ;
        RECT -59.265 393.165 -58.255 393.395 ;
        RECT -59.265 392.905 -59.035 393.165 ;
        RECT -55.260 393.155 -53.760 393.385 ;
        RECT -59.910 392.675 -59.025 392.905 ;
        RECT -59.265 392.415 -59.025 392.675 ;
        RECT -53.530 392.585 -53.240 392.980 ;
        RECT -50.895 392.895 -50.660 393.645 ;
        RECT -42.000 393.435 -41.770 394.430 ;
        RECT -37.995 394.175 -33.810 394.405 ;
        RECT -33.630 393.915 -33.395 394.665 ;
        RECT -35.310 393.685 -33.395 393.915 ;
        RECT -42.000 393.205 -40.990 393.435 ;
        RECT -42.000 392.945 -41.770 393.205 ;
        RECT -37.995 393.195 -36.495 393.425 ;
        RECT -52.575 392.665 -50.660 392.895 ;
        RECT -42.645 392.715 -41.760 392.945 ;
        RECT -51.080 392.660 -50.660 392.665 ;
        RECT -59.265 392.185 -58.255 392.415 ;
        RECT -53.530 392.315 -52.695 392.585 ;
        RECT -53.530 392.185 -53.240 392.315 ;
        RECT -59.265 391.925 -59.025 392.185 ;
        RECT -59.910 391.695 -59.025 391.925 ;
        RECT -59.265 391.435 -59.035 391.695 ;
        RECT -59.265 391.205 -58.255 391.435 ;
        RECT -53.335 390.480 -53.105 391.475 ;
        RECT -52.965 391.215 -52.695 392.315 ;
        RECT -42.000 392.455 -41.760 392.715 ;
        RECT -36.265 392.625 -35.975 393.020 ;
        RECT -33.630 392.935 -33.395 393.685 ;
        RECT -35.310 392.705 -33.395 392.935 ;
        RECT -33.815 392.700 -33.395 392.705 ;
        RECT -42.000 392.225 -40.990 392.455 ;
        RECT -36.265 392.355 -35.430 392.625 ;
        RECT -36.265 392.225 -35.975 392.355 ;
        RECT -42.000 391.965 -41.760 392.225 ;
        RECT -42.645 391.735 -41.760 391.965 ;
        RECT -42.000 391.475 -41.770 391.735 ;
        RECT -42.000 391.245 -40.990 391.475 ;
        RECT -52.965 390.945 -50.975 391.215 ;
        RECT -54.615 390.250 -53.105 390.480 ;
        RECT -53.335 389.990 -53.105 390.250 ;
        RECT -62.860 389.630 -60.945 389.860 ;
        RECT -53.345 389.760 -51.965 389.990 ;
        RECT -62.860 388.880 -62.625 389.630 ;
        RECT -53.345 389.500 -53.105 389.760 ;
        RECT -62.445 389.140 -58.260 389.370 ;
        RECT -54.615 389.270 -53.105 389.500 ;
        RECT -53.345 389.010 -53.105 389.270 ;
        RECT -62.860 388.650 -60.945 388.880 ;
        RECT -53.345 388.780 -51.965 389.010 ;
        RECT -62.860 387.900 -62.625 388.650 ;
        RECT -53.335 388.520 -53.105 388.780 ;
        RECT -59.760 388.160 -58.260 388.390 ;
        RECT -54.615 388.290 -53.105 388.520 ;
        RECT -62.860 387.670 -60.945 387.900 ;
        RECT -62.860 387.665 -62.440 387.670 ;
        RECT -53.445 387.380 -52.695 387.510 ;
        RECT -60.735 387.110 -52.695 387.380 ;
        RECT -60.735 386.395 -60.465 387.110 ;
        RECT -53.445 386.860 -52.695 387.110 ;
        RECT -51.245 385.105 -50.975 390.945 ;
        RECT -36.070 390.520 -35.840 391.515 ;
        RECT -35.700 391.255 -35.430 392.355 ;
        RECT -35.700 390.985 -33.710 391.255 ;
        RECT -37.350 390.290 -35.840 390.520 ;
        RECT -36.070 390.030 -35.840 390.290 ;
        RECT -45.595 389.670 -43.680 389.900 ;
        RECT -36.080 389.800 -34.700 390.030 ;
        RECT -45.595 388.920 -45.360 389.670 ;
        RECT -36.080 389.540 -35.840 389.800 ;
        RECT -45.180 389.180 -40.995 389.410 ;
        RECT -37.350 389.310 -35.840 389.540 ;
        RECT -36.080 389.050 -35.840 389.310 ;
        RECT -45.595 388.690 -43.680 388.920 ;
        RECT -36.080 388.820 -34.700 389.050 ;
        RECT -45.595 387.940 -45.360 388.690 ;
        RECT -36.070 388.560 -35.840 388.820 ;
        RECT -42.495 388.200 -40.995 388.430 ;
        RECT -37.350 388.330 -35.840 388.560 ;
        RECT -45.595 387.710 -43.680 387.940 ;
        RECT -45.595 387.705 -45.175 387.710 ;
        RECT -36.180 387.420 -35.430 387.550 ;
        RECT -43.470 387.150 -35.430 387.420 ;
        RECT -43.470 386.435 -43.200 387.150 ;
        RECT -36.180 386.900 -35.430 387.150 ;
        RECT -33.980 385.360 -33.710 390.985 ;
        RECT -51.720 379.465 -50.710 385.105 ;
        RECT -34.390 383.875 -33.280 385.360 ;
        RECT -31.760 379.465 -30.750 417.250 ;
        RECT -51.720 378.455 -30.750 379.465 ;
        RECT -62.785 377.570 -61.130 377.930 ;
        RECT -62.785 376.245 -23.140 377.570 ;
        RECT -83.945 374.280 -71.620 375.780 ;
        RECT -69.045 374.450 -67.590 376.035 ;
        RECT -83.945 292.695 -82.445 374.280 ;
        RECT -73.505 374.235 -71.620 374.280 ;
        RECT -61.430 374.025 -61.070 374.195 ;
        RECT -62.170 373.700 -61.070 374.025 ;
        RECT -63.835 372.100 -62.335 372.330 ;
        RECT -63.835 369.910 -62.335 370.140 ;
        RECT -62.170 368.925 -61.845 373.700 ;
        RECT -61.430 373.670 -61.070 373.700 ;
        RECT -60.775 372.515 -57.775 372.745 ;
        RECT -54.445 372.415 -54.215 373.410 ;
        RECT -55.225 372.185 -54.215 372.415 ;
        RECT -54.445 371.925 -54.215 372.185 ;
        RECT -54.455 371.695 -53.570 371.925 ;
        RECT -60.775 371.455 -57.775 371.685 ;
        RECT -54.455 371.435 -54.215 371.695 ;
        RECT -55.225 371.205 -54.215 371.435 ;
        RECT -60.775 370.965 -57.775 371.195 ;
        RECT -54.455 370.945 -54.215 371.205 ;
        RECT -43.655 371.385 -43.345 374.850 ;
        RECT -54.455 370.715 -53.570 370.945 ;
        RECT -60.775 370.475 -57.775 370.705 ;
        RECT -54.445 370.455 -54.215 370.715 ;
        RECT -55.225 370.225 -54.215 370.455 ;
        RECT -43.655 370.305 -30.840 371.385 ;
        RECT -60.775 369.420 -57.775 369.650 ;
        RECT -52.535 368.650 -50.620 368.880 ;
        RECT -59.225 367.420 -58.995 368.415 ;
        RECT -55.220 368.160 -51.035 368.390 ;
        RECT -50.855 367.900 -50.620 368.650 ;
        RECT -52.535 367.670 -50.620 367.900 ;
        RECT -59.225 367.190 -58.215 367.420 ;
        RECT -59.225 366.930 -58.995 367.190 ;
        RECT -55.220 367.180 -53.720 367.410 ;
        RECT -59.870 366.700 -58.985 366.930 ;
        RECT -59.225 366.440 -58.985 366.700 ;
        RECT -53.490 366.610 -53.200 367.005 ;
        RECT -50.855 366.920 -50.620 367.670 ;
        RECT -46.125 367.315 -44.625 367.545 ;
        RECT -43.655 367.070 -43.345 370.305 ;
        RECT -52.535 366.690 -50.620 366.920 ;
        RECT -43.700 366.740 -43.285 367.070 ;
        RECT -41.145 366.825 -39.645 367.055 ;
        RECT -51.040 366.685 -50.620 366.690 ;
        RECT -59.225 366.210 -58.215 366.440 ;
        RECT -53.490 366.340 -52.655 366.610 ;
        RECT -53.490 366.210 -53.200 366.340 ;
        RECT -59.225 365.950 -58.985 366.210 ;
        RECT -59.870 365.720 -58.985 365.950 ;
        RECT -59.225 365.460 -58.995 365.720 ;
        RECT -59.225 365.230 -58.215 365.460 ;
        RECT -53.295 364.505 -53.065 365.500 ;
        RECT -52.925 365.240 -52.655 366.340 ;
        RECT -46.125 366.175 -43.625 366.405 ;
        RECT -46.125 365.685 -43.625 365.915 ;
        RECT -43.270 365.880 -42.580 366.150 ;
        RECT -52.925 364.970 -50.935 365.240 ;
        RECT -54.575 364.275 -53.065 364.505 ;
        RECT -53.295 364.015 -53.065 364.275 ;
        RECT -62.820 363.655 -60.905 363.885 ;
        RECT -53.305 363.785 -51.925 364.015 ;
        RECT -62.820 362.905 -62.585 363.655 ;
        RECT -53.305 363.525 -53.065 363.785 ;
        RECT -62.405 363.165 -58.220 363.395 ;
        RECT -54.575 363.295 -53.065 363.525 ;
        RECT -53.305 363.035 -53.065 363.295 ;
        RECT -62.820 362.675 -60.905 362.905 ;
        RECT -53.305 362.805 -51.925 363.035 ;
        RECT -62.820 361.925 -62.585 362.675 ;
        RECT -53.295 362.545 -53.065 362.805 ;
        RECT -59.720 362.185 -58.220 362.415 ;
        RECT -54.575 362.315 -53.065 362.545 ;
        RECT -62.820 361.695 -60.905 361.925 ;
        RECT -62.820 361.690 -62.400 361.695 ;
        RECT -53.405 361.405 -52.655 361.535 ;
        RECT -60.695 361.135 -52.655 361.405 ;
        RECT -60.695 360.420 -60.425 361.135 ;
        RECT -53.405 360.885 -52.655 361.135 ;
        RECT -51.205 360.180 -50.935 364.970 ;
        RECT -43.165 364.645 -42.945 365.880 ;
        RECT -42.145 365.685 -39.645 365.915 ;
        RECT -46.125 364.055 -43.625 364.285 ;
        RECT -43.195 363.955 -42.925 364.645 ;
        RECT -42.145 364.055 -39.645 364.285 ;
        RECT -46.125 363.430 -43.625 363.660 ;
        RECT -46.125 362.940 -43.625 363.170 ;
        RECT -46.125 361.080 -44.625 361.310 ;
        RECT -43.165 360.615 -42.945 363.955 ;
        RECT -42.145 363.405 -39.645 363.635 ;
        RECT -42.145 362.915 -39.645 363.145 ;
        RECT -42.145 362.425 -39.645 362.655 ;
        RECT -42.145 361.080 -39.645 361.310 ;
        RECT -51.235 359.695 -50.905 360.180 ;
        RECT -43.195 359.925 -42.925 360.615 ;
        RECT -44.880 359.575 -44.425 359.635 ;
        RECT -48.440 359.180 -44.425 359.575 ;
        RECT -50.700 357.075 -50.215 357.130 ;
        RECT -48.440 357.075 -48.045 359.180 ;
        RECT -44.880 359.120 -44.425 359.180 ;
        RECT -50.700 356.680 -48.045 357.075 ;
        RECT -50.700 356.550 -50.215 356.680 ;
        RECT -61.275 355.685 -60.915 355.855 ;
        RECT -44.010 355.725 -43.650 355.895 ;
        RECT -62.015 355.360 -60.915 355.685 ;
        RECT -63.680 353.760 -62.180 353.990 ;
        RECT -63.680 351.570 -62.180 351.800 ;
        RECT -62.015 350.585 -61.690 355.360 ;
        RECT -61.275 355.330 -60.915 355.360 ;
        RECT -44.750 355.400 -43.650 355.725 ;
        RECT -60.620 354.175 -57.620 354.405 ;
        RECT -54.290 354.075 -54.060 355.070 ;
        RECT -55.070 353.845 -54.060 354.075 ;
        RECT -54.290 353.585 -54.060 353.845 ;
        RECT -46.415 353.800 -44.915 354.030 ;
        RECT -54.300 353.355 -53.415 353.585 ;
        RECT -60.620 353.115 -57.620 353.345 ;
        RECT -54.300 353.095 -54.060 353.355 ;
        RECT -55.070 352.865 -54.060 353.095 ;
        RECT -60.620 352.625 -57.620 352.855 ;
        RECT -54.300 352.605 -54.060 352.865 ;
        RECT -54.300 352.375 -53.415 352.605 ;
        RECT -60.620 352.135 -57.620 352.365 ;
        RECT -54.290 352.115 -54.060 352.375 ;
        RECT -55.070 351.885 -54.060 352.115 ;
        RECT -46.415 351.610 -44.915 351.840 ;
        RECT -60.620 351.080 -57.620 351.310 ;
        RECT -44.750 350.625 -44.425 355.400 ;
        RECT -44.010 355.370 -43.650 355.400 ;
        RECT -43.355 354.215 -40.355 354.445 ;
        RECT -37.025 354.115 -36.795 355.110 ;
        RECT -37.805 353.885 -36.795 354.115 ;
        RECT -37.025 353.625 -36.795 353.885 ;
        RECT -37.035 353.395 -36.150 353.625 ;
        RECT -43.355 353.155 -40.355 353.385 ;
        RECT -37.035 353.135 -36.795 353.395 ;
        RECT -37.805 352.905 -36.795 353.135 ;
        RECT -43.355 352.665 -40.355 352.895 ;
        RECT -37.035 352.645 -36.795 352.905 ;
        RECT -37.035 352.415 -36.150 352.645 ;
        RECT -43.355 352.175 -40.355 352.405 ;
        RECT -37.025 352.155 -36.795 352.415 ;
        RECT -37.805 351.925 -36.795 352.155 ;
        RECT -43.355 351.120 -40.355 351.350 ;
        RECT -52.380 350.310 -50.465 350.540 ;
        RECT -35.115 350.350 -33.200 350.580 ;
        RECT -59.070 349.080 -58.840 350.075 ;
        RECT -55.065 349.820 -50.880 350.050 ;
        RECT -50.700 349.560 -50.465 350.310 ;
        RECT -52.380 349.330 -50.465 349.560 ;
        RECT -59.070 348.850 -58.060 349.080 ;
        RECT -59.070 348.590 -58.840 348.850 ;
        RECT -55.065 348.840 -53.565 349.070 ;
        RECT -59.715 348.360 -58.830 348.590 ;
        RECT -59.070 348.100 -58.830 348.360 ;
        RECT -53.335 348.270 -53.045 348.665 ;
        RECT -50.700 348.580 -50.465 349.330 ;
        RECT -41.805 349.120 -41.575 350.115 ;
        RECT -37.800 349.860 -33.615 350.090 ;
        RECT -33.435 349.600 -33.200 350.350 ;
        RECT -35.115 349.370 -33.200 349.600 ;
        RECT -41.805 348.890 -40.795 349.120 ;
        RECT -41.805 348.630 -41.575 348.890 ;
        RECT -37.800 348.880 -36.300 349.110 ;
        RECT -52.380 348.350 -50.465 348.580 ;
        RECT -42.450 348.400 -41.565 348.630 ;
        RECT -50.885 348.345 -50.465 348.350 ;
        RECT -59.070 347.870 -58.060 348.100 ;
        RECT -53.335 348.000 -52.500 348.270 ;
        RECT -53.335 347.870 -53.045 348.000 ;
        RECT -59.070 347.610 -58.830 347.870 ;
        RECT -59.715 347.380 -58.830 347.610 ;
        RECT -59.070 347.120 -58.840 347.380 ;
        RECT -59.070 346.890 -58.060 347.120 ;
        RECT -53.140 346.165 -52.910 347.160 ;
        RECT -52.770 346.900 -52.500 348.000 ;
        RECT -41.805 348.140 -41.565 348.400 ;
        RECT -36.070 348.310 -35.780 348.705 ;
        RECT -33.435 348.620 -33.200 349.370 ;
        RECT -35.115 348.390 -33.200 348.620 ;
        RECT -33.620 348.385 -33.200 348.390 ;
        RECT -41.805 347.910 -40.795 348.140 ;
        RECT -36.070 348.040 -35.235 348.310 ;
        RECT -36.070 347.910 -35.780 348.040 ;
        RECT -41.805 347.650 -41.565 347.910 ;
        RECT -42.450 347.420 -41.565 347.650 ;
        RECT -41.805 347.160 -41.575 347.420 ;
        RECT -41.805 346.930 -40.795 347.160 ;
        RECT -52.770 346.630 -50.780 346.900 ;
        RECT -54.420 345.935 -52.910 346.165 ;
        RECT -53.140 345.675 -52.910 345.935 ;
        RECT -62.665 345.315 -60.750 345.545 ;
        RECT -53.150 345.445 -51.770 345.675 ;
        RECT -62.665 344.565 -62.430 345.315 ;
        RECT -53.150 345.185 -52.910 345.445 ;
        RECT -62.250 344.825 -58.065 345.055 ;
        RECT -54.420 344.955 -52.910 345.185 ;
        RECT -53.150 344.695 -52.910 344.955 ;
        RECT -62.665 344.335 -60.750 344.565 ;
        RECT -53.150 344.465 -51.770 344.695 ;
        RECT -62.665 343.585 -62.430 344.335 ;
        RECT -53.140 344.205 -52.910 344.465 ;
        RECT -59.565 343.845 -58.065 344.075 ;
        RECT -54.420 343.975 -52.910 344.205 ;
        RECT -62.665 343.355 -60.750 343.585 ;
        RECT -62.665 343.350 -62.245 343.355 ;
        RECT -53.250 343.065 -52.500 343.195 ;
        RECT -60.540 342.795 -52.500 343.065 ;
        RECT -60.540 342.080 -60.270 342.795 ;
        RECT -53.250 342.545 -52.500 342.795 ;
        RECT -51.050 340.225 -50.780 346.630 ;
        RECT -35.875 346.205 -35.645 347.200 ;
        RECT -35.505 346.940 -35.235 348.040 ;
        RECT -35.505 346.670 -33.515 346.940 ;
        RECT -37.155 345.975 -35.645 346.205 ;
        RECT -35.875 345.715 -35.645 345.975 ;
        RECT -45.400 345.355 -43.485 345.585 ;
        RECT -35.885 345.485 -34.505 345.715 ;
        RECT -45.400 344.605 -45.165 345.355 ;
        RECT -35.885 345.225 -35.645 345.485 ;
        RECT -44.985 344.865 -40.800 345.095 ;
        RECT -37.155 344.995 -35.645 345.225 ;
        RECT -35.885 344.735 -35.645 344.995 ;
        RECT -45.400 344.375 -43.485 344.605 ;
        RECT -35.885 344.505 -34.505 344.735 ;
        RECT -45.400 343.625 -45.165 344.375 ;
        RECT -35.875 344.245 -35.645 344.505 ;
        RECT -42.300 343.885 -40.800 344.115 ;
        RECT -37.155 344.015 -35.645 344.245 ;
        RECT -45.400 343.395 -43.485 343.625 ;
        RECT -45.400 343.390 -44.980 343.395 ;
        RECT -35.985 343.105 -35.235 343.235 ;
        RECT -43.275 342.835 -35.235 343.105 ;
        RECT -43.275 342.120 -43.005 342.835 ;
        RECT -35.985 342.585 -35.235 342.835 ;
        RECT -33.785 341.140 -33.515 346.670 ;
        RECT -68.910 295.950 -68.005 339.950 ;
        RECT -51.320 336.930 -50.365 340.225 ;
        RECT -34.170 339.355 -32.835 341.140 ;
        RECT -31.795 336.930 -30.840 370.305 ;
        RECT -51.320 335.975 -30.840 336.930 ;
        RECT -33.615 335.250 -33.345 335.280 ;
        RECT -34.000 335.165 -32.665 335.250 ;
        RECT -61.445 335.115 -25.250 335.165 ;
        RECT -62.290 334.000 -25.250 335.115 ;
        RECT -61.445 333.920 -25.250 334.000 ;
        RECT -34.000 333.465 -32.665 333.920 ;
        RECT -61.375 331.825 -61.015 331.995 ;
        RECT -62.115 331.500 -61.015 331.825 ;
        RECT -63.780 329.900 -62.280 330.130 ;
        RECT -63.780 327.710 -62.280 327.940 ;
        RECT -62.115 326.725 -61.790 331.500 ;
        RECT -61.375 331.470 -61.015 331.500 ;
        RECT -60.720 330.315 -57.720 330.545 ;
        RECT -54.390 330.215 -54.160 331.210 ;
        RECT -55.170 329.985 -54.160 330.215 ;
        RECT -54.390 329.725 -54.160 329.985 ;
        RECT -54.400 329.495 -53.515 329.725 ;
        RECT -60.720 329.255 -57.720 329.485 ;
        RECT -54.400 329.235 -54.160 329.495 ;
        RECT -55.170 329.005 -54.160 329.235 ;
        RECT -60.720 328.765 -57.720 328.995 ;
        RECT -54.400 328.745 -54.160 329.005 ;
        RECT -54.400 328.515 -53.515 328.745 ;
        RECT -60.720 328.275 -57.720 328.505 ;
        RECT -54.390 328.255 -54.160 328.515 ;
        RECT -55.170 328.025 -54.160 328.255 ;
        RECT -43.600 328.385 -43.290 332.650 ;
        RECT -43.600 327.540 -31.210 328.385 ;
        RECT -60.720 327.220 -57.720 327.450 ;
        RECT -52.480 326.450 -50.565 326.680 ;
        RECT -59.170 325.220 -58.940 326.215 ;
        RECT -55.165 325.960 -50.980 326.190 ;
        RECT -50.800 325.700 -50.565 326.450 ;
        RECT -52.480 325.470 -50.565 325.700 ;
        RECT -59.170 324.990 -58.160 325.220 ;
        RECT -59.170 324.730 -58.940 324.990 ;
        RECT -55.165 324.980 -53.665 325.210 ;
        RECT -59.815 324.500 -58.930 324.730 ;
        RECT -59.170 324.240 -58.930 324.500 ;
        RECT -53.435 324.410 -53.145 324.805 ;
        RECT -50.800 324.720 -50.565 325.470 ;
        RECT -46.070 325.115 -44.570 325.345 ;
        RECT -43.600 324.870 -43.290 327.540 ;
        RECT -52.480 324.490 -50.565 324.720 ;
        RECT -43.645 324.540 -43.230 324.870 ;
        RECT -41.090 324.625 -39.590 324.855 ;
        RECT -50.985 324.485 -50.565 324.490 ;
        RECT -59.170 324.010 -58.160 324.240 ;
        RECT -53.435 324.140 -52.600 324.410 ;
        RECT -53.435 324.010 -53.145 324.140 ;
        RECT -59.170 323.750 -58.930 324.010 ;
        RECT -59.815 323.520 -58.930 323.750 ;
        RECT -59.170 323.260 -58.940 323.520 ;
        RECT -59.170 323.030 -58.160 323.260 ;
        RECT -53.240 322.305 -53.010 323.300 ;
        RECT -52.870 323.040 -52.600 324.140 ;
        RECT -46.070 323.975 -43.570 324.205 ;
        RECT -46.070 323.485 -43.570 323.715 ;
        RECT -43.215 323.680 -42.525 323.950 ;
        RECT -52.870 322.770 -50.880 323.040 ;
        RECT -54.520 322.075 -53.010 322.305 ;
        RECT -53.240 321.815 -53.010 322.075 ;
        RECT -62.765 321.455 -60.850 321.685 ;
        RECT -53.250 321.585 -51.870 321.815 ;
        RECT -62.765 320.705 -62.530 321.455 ;
        RECT -53.250 321.325 -53.010 321.585 ;
        RECT -62.350 320.965 -58.165 321.195 ;
        RECT -54.520 321.095 -53.010 321.325 ;
        RECT -53.250 320.835 -53.010 321.095 ;
        RECT -62.765 320.475 -60.850 320.705 ;
        RECT -53.250 320.605 -51.870 320.835 ;
        RECT -62.765 319.725 -62.530 320.475 ;
        RECT -53.240 320.345 -53.010 320.605 ;
        RECT -59.665 319.985 -58.165 320.215 ;
        RECT -54.520 320.115 -53.010 320.345 ;
        RECT -62.765 319.495 -60.850 319.725 ;
        RECT -62.765 319.490 -62.345 319.495 ;
        RECT -53.350 319.205 -52.600 319.335 ;
        RECT -60.640 318.935 -52.600 319.205 ;
        RECT -60.640 318.220 -60.370 318.935 ;
        RECT -53.350 318.685 -52.600 318.935 ;
        RECT -51.150 317.980 -50.880 322.770 ;
        RECT -43.110 322.445 -42.890 323.680 ;
        RECT -42.090 323.485 -39.590 323.715 ;
        RECT -46.070 321.855 -43.570 322.085 ;
        RECT -43.140 321.755 -42.870 322.445 ;
        RECT -42.090 321.855 -39.590 322.085 ;
        RECT -46.070 321.230 -43.570 321.460 ;
        RECT -46.070 320.740 -43.570 320.970 ;
        RECT -46.070 318.880 -44.570 319.110 ;
        RECT -43.110 318.415 -42.890 321.755 ;
        RECT -42.090 321.205 -39.590 321.435 ;
        RECT -42.090 320.715 -39.590 320.945 ;
        RECT -42.090 320.225 -39.590 320.455 ;
        RECT -42.090 318.880 -39.590 319.110 ;
        RECT -51.180 317.495 -50.850 317.980 ;
        RECT -43.140 317.725 -42.870 318.415 ;
        RECT -44.825 317.375 -44.370 317.435 ;
        RECT -48.385 316.980 -44.370 317.375 ;
        RECT -50.645 314.875 -50.160 314.930 ;
        RECT -48.385 314.875 -47.990 316.980 ;
        RECT -44.825 316.920 -44.370 316.980 ;
        RECT -50.645 314.480 -47.990 314.875 ;
        RECT -50.645 314.350 -50.160 314.480 ;
        RECT -61.220 313.485 -60.860 313.655 ;
        RECT -43.955 313.525 -43.595 313.695 ;
        RECT -61.960 313.160 -60.860 313.485 ;
        RECT -63.625 311.560 -62.125 311.790 ;
        RECT -63.625 309.370 -62.125 309.600 ;
        RECT -61.960 308.385 -61.635 313.160 ;
        RECT -61.220 313.130 -60.860 313.160 ;
        RECT -44.695 313.200 -43.595 313.525 ;
        RECT -60.565 311.975 -57.565 312.205 ;
        RECT -54.235 311.875 -54.005 312.870 ;
        RECT -55.015 311.645 -54.005 311.875 ;
        RECT -54.235 311.385 -54.005 311.645 ;
        RECT -46.360 311.600 -44.860 311.830 ;
        RECT -54.245 311.155 -53.360 311.385 ;
        RECT -60.565 310.915 -57.565 311.145 ;
        RECT -54.245 310.895 -54.005 311.155 ;
        RECT -55.015 310.665 -54.005 310.895 ;
        RECT -60.565 310.425 -57.565 310.655 ;
        RECT -54.245 310.405 -54.005 310.665 ;
        RECT -54.245 310.175 -53.360 310.405 ;
        RECT -60.565 309.935 -57.565 310.165 ;
        RECT -54.235 309.915 -54.005 310.175 ;
        RECT -55.015 309.685 -54.005 309.915 ;
        RECT -46.360 309.410 -44.860 309.640 ;
        RECT -60.565 308.880 -57.565 309.110 ;
        RECT -44.695 308.425 -44.370 313.200 ;
        RECT -43.955 313.170 -43.595 313.200 ;
        RECT -43.300 312.015 -40.300 312.245 ;
        RECT -36.970 311.915 -36.740 312.910 ;
        RECT -37.750 311.685 -36.740 311.915 ;
        RECT -36.970 311.425 -36.740 311.685 ;
        RECT -36.980 311.195 -36.095 311.425 ;
        RECT -43.300 310.955 -40.300 311.185 ;
        RECT -36.980 310.935 -36.740 311.195 ;
        RECT -37.750 310.705 -36.740 310.935 ;
        RECT -43.300 310.465 -40.300 310.695 ;
        RECT -36.980 310.445 -36.740 310.705 ;
        RECT -36.980 310.215 -36.095 310.445 ;
        RECT -43.300 309.975 -40.300 310.205 ;
        RECT -36.970 309.955 -36.740 310.215 ;
        RECT -37.750 309.725 -36.740 309.955 ;
        RECT -43.300 308.920 -40.300 309.150 ;
        RECT -52.325 308.110 -50.410 308.340 ;
        RECT -35.060 308.150 -33.145 308.380 ;
        RECT -59.015 306.880 -58.785 307.875 ;
        RECT -55.010 307.620 -50.825 307.850 ;
        RECT -50.645 307.360 -50.410 308.110 ;
        RECT -52.325 307.130 -50.410 307.360 ;
        RECT -59.015 306.650 -58.005 306.880 ;
        RECT -59.015 306.390 -58.785 306.650 ;
        RECT -55.010 306.640 -53.510 306.870 ;
        RECT -59.660 306.160 -58.775 306.390 ;
        RECT -59.015 305.900 -58.775 306.160 ;
        RECT -53.280 306.070 -52.990 306.465 ;
        RECT -50.645 306.380 -50.410 307.130 ;
        RECT -41.750 306.920 -41.520 307.915 ;
        RECT -37.745 307.660 -33.560 307.890 ;
        RECT -33.380 307.400 -33.145 308.150 ;
        RECT -35.060 307.170 -33.145 307.400 ;
        RECT -41.750 306.690 -40.740 306.920 ;
        RECT -41.750 306.430 -41.520 306.690 ;
        RECT -37.745 306.680 -36.245 306.910 ;
        RECT -52.325 306.150 -50.410 306.380 ;
        RECT -42.395 306.200 -41.510 306.430 ;
        RECT -33.380 306.420 -33.145 307.170 ;
        RECT -50.830 306.145 -50.410 306.150 ;
        RECT -59.015 305.670 -58.005 305.900 ;
        RECT -53.280 305.800 -52.445 306.070 ;
        RECT -53.280 305.670 -52.990 305.800 ;
        RECT -59.015 305.410 -58.775 305.670 ;
        RECT -59.660 305.180 -58.775 305.410 ;
        RECT -59.015 304.920 -58.785 305.180 ;
        RECT -59.015 304.690 -58.005 304.920 ;
        RECT -53.085 303.965 -52.855 304.960 ;
        RECT -52.715 304.700 -52.445 305.800 ;
        RECT -41.750 305.940 -41.510 306.200 ;
        RECT -35.060 306.190 -33.145 306.420 ;
        RECT -33.565 306.185 -33.145 306.190 ;
        RECT -41.750 305.710 -40.740 305.940 ;
        RECT -41.750 305.450 -41.510 305.710 ;
        RECT -42.395 305.220 -41.510 305.450 ;
        RECT -41.750 304.960 -41.520 305.220 ;
        RECT -41.750 304.730 -40.740 304.960 ;
        RECT -52.715 304.430 -50.725 304.700 ;
        RECT -54.365 303.735 -52.855 303.965 ;
        RECT -53.085 303.475 -52.855 303.735 ;
        RECT -62.610 303.115 -60.695 303.345 ;
        RECT -53.095 303.245 -51.715 303.475 ;
        RECT -62.610 302.365 -62.375 303.115 ;
        RECT -53.095 302.985 -52.855 303.245 ;
        RECT -62.195 302.625 -58.010 302.855 ;
        RECT -54.365 302.755 -52.855 302.985 ;
        RECT -53.095 302.495 -52.855 302.755 ;
        RECT -62.610 302.135 -60.695 302.365 ;
        RECT -53.095 302.265 -51.715 302.495 ;
        RECT -62.610 301.385 -62.375 302.135 ;
        RECT -53.085 302.005 -52.855 302.265 ;
        RECT -59.510 301.645 -58.010 301.875 ;
        RECT -54.365 301.775 -52.855 302.005 ;
        RECT -62.610 301.155 -60.695 301.385 ;
        RECT -62.610 301.150 -62.190 301.155 ;
        RECT -53.195 300.865 -52.445 300.995 ;
        RECT -60.485 300.595 -52.445 300.865 ;
        RECT -60.485 299.880 -60.215 300.595 ;
        RECT -53.195 300.345 -52.445 300.595 ;
        RECT -50.995 297.810 -50.725 304.430 ;
        RECT -35.820 304.005 -35.590 305.000 ;
        RECT -37.100 303.775 -35.590 304.005 ;
        RECT -35.820 303.515 -35.590 303.775 ;
        RECT -45.345 303.155 -43.430 303.385 ;
        RECT -35.830 303.285 -34.450 303.515 ;
        RECT -45.345 302.405 -45.110 303.155 ;
        RECT -35.830 303.025 -35.590 303.285 ;
        RECT -44.930 302.665 -40.745 302.895 ;
        RECT -37.100 302.795 -35.590 303.025 ;
        RECT -35.830 302.535 -35.590 302.795 ;
        RECT -45.345 302.175 -43.430 302.405 ;
        RECT -35.830 302.305 -34.450 302.535 ;
        RECT -45.345 301.425 -45.110 302.175 ;
        RECT -35.820 302.045 -35.590 302.305 ;
        RECT -42.245 301.685 -40.745 301.915 ;
        RECT -37.100 301.815 -35.590 302.045 ;
        RECT -45.345 301.195 -43.430 301.425 ;
        RECT -45.345 301.190 -44.925 301.195 ;
        RECT -35.930 300.905 -35.180 301.035 ;
        RECT -43.220 300.635 -35.180 300.905 ;
        RECT -43.220 299.920 -42.950 300.635 ;
        RECT -35.930 300.385 -35.180 300.635 ;
        RECT -51.140 296.905 -50.295 297.810 ;
        RECT -32.055 296.905 -31.210 327.540 ;
        RECT -51.140 296.060 -31.210 296.905 ;
        RECT -83.945 292.090 -52.110 292.695 ;
        RECT -83.945 286.890 -82.445 292.090 ;
        RECT -71.240 291.425 -57.350 291.555 ;
        RECT -71.240 291.255 -56.540 291.425 ;
        RECT -71.240 290.950 -57.350 291.255 ;
        RECT -86.060 285.155 -85.455 285.865 ;
        RECT -71.240 285.155 -70.635 290.950 ;
        RECT -68.990 288.470 -67.890 289.380 ;
        RECT -57.035 288.470 -56.865 290.985 ;
        RECT -68.990 288.120 -56.865 288.470 ;
        RECT -68.990 287.525 -67.890 288.120 ;
        RECT -86.060 284.550 -70.635 285.155 ;
        RECT -57.035 280.505 -56.865 288.120 ;
        RECT -56.710 285.055 -56.540 291.255 ;
        RECT -52.450 289.925 -52.225 292.090 ;
        RECT -48.275 291.265 -35.205 292.040 ;
        RECT -52.495 289.335 -52.205 289.925 ;
        RECT -56.365 288.900 -52.865 289.130 ;
        RECT -51.940 288.900 -48.440 289.130 ;
        RECT -56.365 286.900 -52.865 287.130 ;
        RECT -51.940 286.900 -48.440 287.130 ;
        RECT -48.275 286.130 -47.925 291.265 ;
        RECT -41.990 290.340 -41.670 290.955 ;
        RECT -51.930 285.780 -47.925 286.130 ;
        RECT -52.555 285.055 -52.265 285.445 ;
        RECT -56.710 284.885 -52.265 285.055 ;
        RECT -52.555 284.855 -52.265 284.885 ;
        RECT -56.365 283.900 -52.865 284.130 ;
        RECT -51.940 283.900 -48.440 284.130 ;
        RECT -56.365 281.900 -52.865 282.130 ;
        RECT -51.940 281.900 -48.440 282.130 ;
        RECT -48.275 281.175 -47.925 285.780 ;
        RECT -51.925 280.825 -47.925 281.175 ;
        RECT -57.035 280.335 -52.190 280.505 ;
        RECT -52.360 280.060 -52.190 280.335 ;
        RECT -52.420 279.470 -52.130 280.060 ;
        RECT -56.365 278.900 -52.865 279.130 ;
        RECT -51.940 278.900 -48.440 279.130 ;
        RECT -56.365 276.900 -52.865 277.130 ;
        RECT -51.940 276.900 -48.440 277.130 ;
        RECT -48.275 275.955 -47.925 280.825 ;
        RECT -49.170 275.605 -47.925 275.955 ;
        RECT -46.790 289.910 -41.670 290.340 ;
        RECT -46.790 289.890 -41.435 289.910 ;
        RECT -56.720 274.460 -55.720 274.690 ;
        RECT -54.820 274.460 -54.320 274.690 ;
        RECT -51.150 274.625 -47.585 274.910 ;
        RECT -51.150 274.480 -50.480 274.625 ;
        RECT -52.485 273.800 -51.485 274.030 ;
        RECT -50.215 273.730 -48.215 273.960 ;
        RECT -56.720 273.480 -55.720 273.710 ;
        RECT -54.820 273.480 -54.320 273.710 ;
        RECT -52.485 273.310 -51.485 273.540 ;
        RECT -52.485 272.750 -51.485 272.980 ;
        RECT -50.215 272.750 -48.215 272.980 ;
        RECT -56.720 272.500 -55.720 272.730 ;
        RECT -54.820 272.500 -54.320 272.730 ;
        RECT -51.235 272.210 -50.945 272.215 ;
        RECT -55.310 270.805 -55.010 272.140 ;
        RECT -51.240 270.805 -50.940 272.210 ;
        RECT -48.820 270.805 -48.160 270.965 ;
        RECT -55.310 270.505 -48.160 270.805 ;
        RECT -54.460 270.110 -54.160 270.270 ;
        RECT -50.735 270.110 -50.435 270.310 ;
        RECT -48.820 270.165 -48.160 270.505 ;
        RECT -54.460 269.810 -50.435 270.110 ;
        RECT -54.460 269.615 -54.160 269.810 ;
        RECT -50.735 269.650 -50.435 269.810 ;
        RECT -56.755 268.855 -55.755 269.085 ;
        RECT -53.215 268.855 -52.215 269.085 ;
        RECT -53.715 266.790 -52.215 267.020 ;
        RECT -53.715 266.300 -52.215 266.530 ;
        RECT -53.715 265.810 -52.215 266.040 ;
        RECT -56.755 265.165 -55.755 265.395 ;
        RECT -53.715 265.245 -52.215 265.475 ;
        RECT -53.715 264.755 -52.215 264.985 ;
        RECT -56.755 264.185 -55.755 264.415 ;
        RECT -53.715 264.265 -52.215 264.495 ;
        RECT -53.720 263.695 -52.220 263.925 ;
        RECT -56.755 263.205 -55.755 263.435 ;
        RECT -53.720 262.715 -52.220 262.945 ;
        RECT -55.975 261.950 -55.315 262.000 ;
        RECT -55.975 261.740 -50.695 261.950 ;
        RECT -55.975 261.700 -55.315 261.740 ;
        RECT -54.725 261.125 -54.065 261.425 ;
        RECT -56.585 260.660 -54.585 260.890 ;
        RECT -56.585 260.170 -54.585 260.400 ;
        RECT -56.585 259.680 -54.585 259.910 ;
        RECT -56.585 258.625 -54.585 258.855 ;
        RECT -54.425 256.590 -54.215 261.125 ;
        RECT -54.020 259.300 -53.720 259.960 ;
        RECT -53.985 257.365 -53.775 259.300 ;
        RECT -53.125 259.115 -52.125 259.345 ;
        RECT -53.620 258.185 -53.320 258.845 ;
        RECT -50.905 258.310 -50.695 261.740 ;
        RECT -47.870 258.835 -47.585 274.625 ;
        RECT -46.790 270.980 -46.340 289.890 ;
        RECT -42.120 289.610 -41.435 289.890 ;
        RECT -45.455 289.110 -44.455 289.340 ;
        RECT -43.555 289.110 -43.055 289.340 ;
        RECT -40.265 288.620 -39.765 288.850 ;
        RECT -38.865 288.620 -37.865 288.850 ;
        RECT -45.455 288.130 -44.455 288.360 ;
        RECT -43.555 288.130 -43.055 288.360 ;
        RECT -40.265 287.640 -39.765 287.870 ;
        RECT -38.865 287.640 -37.865 287.870 ;
        RECT -45.455 287.150 -44.455 287.380 ;
        RECT -43.555 287.150 -43.055 287.380 ;
        RECT -40.265 286.660 -39.765 286.890 ;
        RECT -38.865 286.660 -37.865 286.890 ;
        RECT -42.270 286.045 -41.970 286.225 ;
        RECT -42.270 285.745 -39.635 286.045 ;
        RECT -42.270 285.565 -41.970 285.745 ;
        RECT -39.415 285.455 -37.955 285.740 ;
        RECT -43.080 285.150 -42.070 285.160 ;
        RECT -45.380 284.920 -44.880 285.150 ;
        RECT -43.305 284.920 -42.070 285.150 ;
        RECT -45.380 284.430 -44.880 284.660 ;
        RECT -43.305 284.430 -42.805 284.660 ;
        RECT -42.310 284.200 -42.070 284.920 ;
        RECT -40.265 284.435 -39.765 284.665 ;
        RECT -42.900 284.170 -42.070 284.200 ;
        RECT -45.380 283.940 -44.880 284.170 ;
        RECT -43.305 283.940 -42.070 284.170 ;
        RECT -42.900 283.895 -42.070 283.940 ;
        RECT -45.380 283.450 -44.880 283.680 ;
        RECT -43.305 283.450 -42.805 283.680 ;
        RECT -42.310 283.220 -42.070 283.895 ;
        RECT -40.265 283.455 -39.765 283.685 ;
        RECT -42.910 283.190 -42.070 283.220 ;
        RECT -45.380 282.960 -44.880 283.190 ;
        RECT -43.305 282.960 -42.070 283.190 ;
        RECT -42.910 282.915 -42.070 282.960 ;
        RECT -45.380 282.470 -44.880 282.700 ;
        RECT -43.305 282.470 -42.805 282.700 ;
        RECT -45.380 281.980 -44.880 282.210 ;
        RECT -45.380 281.490 -44.880 281.720 ;
        RECT -44.240 281.505 -43.870 282.350 ;
        RECT -42.310 282.265 -42.070 282.915 ;
        RECT -40.265 282.475 -39.765 282.705 ;
        RECT -42.900 282.210 -42.070 282.265 ;
        RECT -43.305 281.980 -42.070 282.210 ;
        RECT -42.900 281.960 -42.070 281.980 ;
        RECT -45.455 280.395 -44.455 280.625 ;
        RECT -45.455 279.415 -44.455 279.645 ;
        RECT -45.455 278.435 -44.455 278.665 ;
        RECT -44.190 277.645 -43.905 281.505 ;
        RECT -43.305 281.490 -42.805 281.720 ;
        RECT -43.555 280.395 -43.055 280.625 ;
        RECT -43.555 279.415 -43.055 279.645 ;
        RECT -43.555 278.435 -43.055 278.665 ;
        RECT -45.365 277.360 -43.905 277.645 ;
        RECT -42.310 277.710 -42.070 281.960 ;
        RECT -40.515 281.380 -40.015 281.610 ;
        RECT -39.415 281.595 -39.130 285.455 ;
        RECT -38.865 284.435 -37.865 284.665 ;
        RECT -38.865 283.455 -37.865 283.685 ;
        RECT -38.865 282.475 -37.865 282.705 ;
        RECT -40.515 280.890 -40.015 281.120 ;
        RECT -39.450 280.750 -39.080 281.595 ;
        RECT -38.440 281.380 -37.940 281.610 ;
        RECT -38.440 280.890 -37.940 281.120 ;
        RECT -40.515 280.400 -40.015 280.630 ;
        RECT -38.440 280.400 -37.940 280.630 ;
        RECT -40.515 279.910 -40.015 280.140 ;
        RECT -38.440 279.910 -37.940 280.140 ;
        RECT -40.515 279.420 -40.015 279.650 ;
        RECT -38.440 279.420 -37.940 279.650 ;
        RECT -40.515 278.930 -40.015 279.160 ;
        RECT -38.440 278.930 -37.940 279.160 ;
        RECT -40.515 278.440 -40.015 278.670 ;
        RECT -38.440 278.440 -37.940 278.670 ;
        RECT -40.515 277.950 -40.015 278.180 ;
        RECT -39.645 277.710 -39.345 278.185 ;
        RECT -38.440 277.950 -37.940 278.180 ;
        RECT -42.310 277.505 -39.340 277.710 ;
        RECT -39.645 277.500 -39.345 277.505 ;
        RECT -43.940 276.535 -43.280 276.540 ;
        RECT -43.940 276.240 -39.210 276.535 ;
        RECT -43.505 276.235 -39.210 276.240 ;
        RECT -45.455 275.610 -44.455 275.840 ;
        RECT -43.555 275.610 -43.055 275.840 ;
        RECT -39.540 275.820 -39.240 276.235 ;
        RECT -40.265 275.120 -39.765 275.350 ;
        RECT -38.865 275.120 -37.865 275.350 ;
        RECT -45.455 274.630 -44.455 274.860 ;
        RECT -43.555 274.630 -43.055 274.860 ;
        RECT -40.265 274.140 -39.765 274.370 ;
        RECT -38.865 274.140 -37.865 274.370 ;
        RECT -45.455 273.650 -44.455 273.880 ;
        RECT -43.555 273.650 -43.055 273.880 ;
        RECT -40.265 273.160 -39.765 273.390 ;
        RECT -38.865 273.160 -37.865 273.390 ;
        RECT -39.415 271.955 -37.955 272.240 ;
        RECT -45.380 271.420 -44.880 271.650 ;
        RECT -43.305 271.635 -42.805 271.650 ;
        RECT -43.305 271.405 -42.090 271.635 ;
        RECT -47.245 270.180 -46.340 270.980 ;
        RECT -45.380 270.930 -44.880 271.160 ;
        RECT -43.305 270.930 -42.805 271.160 ;
        RECT -45.380 270.440 -44.880 270.670 ;
        RECT -43.305 270.660 -42.805 270.670 ;
        RECT -42.320 270.660 -42.090 271.405 ;
        RECT -40.265 270.935 -39.765 271.165 ;
        RECT -43.305 270.450 -42.090 270.660 ;
        RECT -43.305 270.440 -42.805 270.450 ;
        RECT -45.380 269.950 -44.880 270.180 ;
        RECT -43.305 269.950 -42.805 270.180 ;
        RECT -45.380 269.460 -44.880 269.690 ;
        RECT -43.305 269.685 -42.805 269.690 ;
        RECT -42.320 269.685 -42.090 270.450 ;
        RECT -40.265 269.955 -39.765 270.185 ;
        RECT -43.305 269.475 -42.090 269.685 ;
        RECT -43.305 269.460 -42.805 269.475 ;
        RECT -45.380 268.970 -44.880 269.200 ;
        RECT -43.305 268.970 -42.805 269.200 ;
        RECT -45.380 268.480 -44.880 268.710 ;
        RECT -45.380 267.990 -44.880 268.220 ;
        RECT -44.240 268.005 -43.870 268.850 ;
        RECT -43.305 268.705 -42.805 268.710 ;
        RECT -42.320 268.705 -42.090 269.475 ;
        RECT -40.265 268.975 -39.765 269.205 ;
        RECT -43.305 268.495 -42.090 268.705 ;
        RECT -43.305 268.480 -42.805 268.495 ;
        RECT -45.455 266.895 -44.455 267.125 ;
        RECT -45.455 265.915 -44.455 266.145 ;
        RECT -45.455 264.935 -44.455 265.165 ;
        RECT -44.190 264.145 -43.905 268.005 ;
        RECT -43.305 267.990 -42.805 268.220 ;
        RECT -42.320 268.065 -42.090 268.495 ;
        RECT -42.320 267.835 -41.030 268.065 ;
        RECT -40.515 267.880 -40.015 268.110 ;
        RECT -39.415 268.095 -39.130 271.955 ;
        RECT -38.865 270.935 -37.865 271.165 ;
        RECT -38.865 269.955 -37.865 270.185 ;
        RECT -38.865 268.975 -37.865 269.205 ;
        RECT -43.555 266.895 -43.055 267.125 ;
        RECT -43.555 265.915 -43.055 266.145 ;
        RECT -43.555 264.935 -43.055 265.165 ;
        RECT -41.260 264.200 -41.030 267.835 ;
        RECT -40.515 267.390 -40.015 267.620 ;
        RECT -39.450 267.250 -39.080 268.095 ;
        RECT -38.440 267.880 -37.940 268.110 ;
        RECT -38.440 267.390 -37.940 267.620 ;
        RECT -40.515 266.900 -40.015 267.130 ;
        RECT -38.440 266.900 -37.940 267.130 ;
        RECT -40.515 266.410 -40.015 266.640 ;
        RECT -38.440 266.410 -37.940 266.640 ;
        RECT -40.515 265.920 -40.015 266.150 ;
        RECT -38.440 265.920 -37.940 266.150 ;
        RECT -40.515 265.430 -40.015 265.660 ;
        RECT -38.440 265.430 -37.940 265.660 ;
        RECT -40.515 264.940 -40.015 265.170 ;
        RECT -38.440 264.940 -37.940 265.170 ;
        RECT -40.515 264.450 -40.015 264.680 ;
        RECT -39.655 264.200 -39.355 264.740 ;
        RECT -38.440 264.450 -37.940 264.680 ;
        RECT -45.365 263.860 -41.435 264.145 ;
        RECT -41.260 264.010 -39.355 264.200 ;
        RECT -41.255 263.970 -39.355 264.010 ;
        RECT -44.060 263.445 -43.400 263.455 ;
        RECT -42.260 263.445 -41.960 263.610 ;
        RECT -44.060 263.155 -41.960 263.445 ;
        RECT -42.260 262.950 -41.960 263.155 ;
        RECT -41.720 263.100 -41.435 263.860 ;
        RECT -41.720 262.815 -40.545 263.100 ;
        RECT -45.455 262.485 -44.455 262.715 ;
        RECT -43.555 262.485 -43.055 262.715 ;
        RECT -45.455 261.505 -44.455 261.735 ;
        RECT -43.555 261.505 -43.055 261.735 ;
        RECT -45.455 260.525 -44.455 260.755 ;
        RECT -43.555 260.525 -43.055 260.755 ;
        RECT -40.830 258.835 -40.545 262.815 ;
        RECT -47.870 258.550 -40.545 258.835 ;
        RECT -40.525 258.310 -40.225 258.350 ;
        RECT -53.565 257.815 -53.355 258.185 ;
        RECT -50.905 258.100 -40.205 258.310 ;
        RECT -53.565 257.605 -50.340 257.815 ;
        RECT -53.985 257.155 -50.710 257.365 ;
        RECT -53.650 256.590 -53.350 256.605 ;
        RECT -54.425 256.380 -53.350 256.590 ;
        RECT -56.585 255.930 -54.585 256.160 ;
        RECT -53.650 255.945 -53.350 256.380 ;
        RECT -56.585 255.440 -54.585 255.670 ;
        RECT -56.585 254.950 -54.585 255.180 ;
        RECT -53.125 254.385 -52.125 254.615 ;
        RECT -56.585 253.895 -54.585 254.125 ;
        RECT -83.320 250.610 -64.110 251.250 ;
        RECT -83.320 250.585 -82.640 250.610 ;
        RECT -64.430 249.270 -64.110 250.610 ;
        RECT -50.920 250.310 -50.710 257.155 ;
        RECT -50.550 253.655 -50.340 257.605 ;
        RECT -44.855 257.505 -41.855 257.735 ;
        RECT -40.525 257.690 -40.225 258.100 ;
        RECT -44.855 257.015 -41.855 257.245 ;
        RECT -44.855 256.525 -41.855 256.755 ;
        RECT -44.855 255.960 -41.855 256.190 ;
        RECT -44.855 255.470 -41.855 255.700 ;
        RECT -40.035 255.390 -39.035 255.620 ;
        RECT -44.855 254.980 -41.855 255.210 ;
        RECT -40.035 254.410 -39.035 254.640 ;
        RECT -44.855 253.920 -41.855 254.150 ;
        RECT -50.550 253.645 -49.570 253.655 ;
        RECT -50.550 252.665 -48.560 253.645 ;
        RECT -50.550 252.630 -50.340 252.665 ;
        RECT -64.665 248.970 -63.980 249.270 ;
        RECT -63.045 248.470 -62.545 248.700 ;
        RECT -61.645 248.470 -60.645 248.700 ;
        RECT -68.235 247.980 -67.235 248.210 ;
        RECT -66.335 247.980 -65.835 248.210 ;
        RECT -63.045 247.490 -62.545 247.720 ;
        RECT -61.645 247.490 -60.645 247.720 ;
        RECT -68.235 247.000 -67.235 247.230 ;
        RECT -66.335 247.000 -65.835 247.230 ;
        RECT -63.045 246.510 -62.545 246.740 ;
        RECT -61.645 246.510 -60.645 246.740 ;
        RECT -68.235 246.020 -67.235 246.250 ;
        RECT -66.335 246.020 -65.835 246.250 ;
        RECT -64.130 245.405 -63.830 245.585 ;
        RECT -66.465 245.105 -63.830 245.405 ;
        RECT -68.145 244.815 -66.685 245.100 ;
        RECT -64.130 244.925 -63.830 245.105 ;
        RECT -68.235 243.795 -67.235 244.025 ;
        RECT -68.235 242.815 -67.235 243.045 ;
        RECT -68.235 241.835 -67.235 242.065 ;
        RECT -68.160 240.740 -67.660 240.970 ;
        RECT -66.970 240.955 -66.685 244.815 ;
        RECT -64.030 244.510 -63.020 244.520 ;
        RECT -64.030 244.280 -62.795 244.510 ;
        RECT -61.220 244.280 -60.720 244.510 ;
        RECT -66.335 243.795 -65.835 244.025 ;
        RECT -64.030 243.560 -63.790 244.280 ;
        RECT -63.295 243.790 -62.795 244.020 ;
        RECT -61.220 243.790 -60.720 244.020 ;
        RECT -64.030 243.530 -63.200 243.560 ;
        RECT -64.030 243.300 -62.795 243.530 ;
        RECT -61.220 243.300 -60.720 243.530 ;
        RECT -64.030 243.255 -63.200 243.300 ;
        RECT -66.335 242.815 -65.835 243.045 ;
        RECT -64.030 242.580 -63.790 243.255 ;
        RECT -63.295 242.810 -62.795 243.040 ;
        RECT -61.220 242.810 -60.720 243.040 ;
        RECT -64.030 242.550 -63.190 242.580 ;
        RECT -64.030 242.320 -62.795 242.550 ;
        RECT -61.220 242.320 -60.720 242.550 ;
        RECT -64.030 242.275 -63.190 242.320 ;
        RECT -66.335 241.835 -65.835 242.065 ;
        RECT -64.030 241.625 -63.790 242.275 ;
        RECT -63.295 241.830 -62.795 242.060 ;
        RECT -61.220 241.830 -60.720 242.060 ;
        RECT -64.030 241.570 -63.200 241.625 ;
        RECT -64.030 241.340 -62.795 241.570 ;
        RECT -64.030 241.320 -63.200 241.340 ;
        RECT -68.160 240.250 -67.660 240.480 ;
        RECT -67.020 240.110 -66.650 240.955 ;
        RECT -66.085 240.740 -65.585 240.970 ;
        RECT -66.085 240.250 -65.585 240.480 ;
        RECT -68.160 239.760 -67.660 239.990 ;
        RECT -66.085 239.760 -65.585 239.990 ;
        RECT -68.160 239.270 -67.660 239.500 ;
        RECT -66.085 239.270 -65.585 239.500 ;
        RECT -68.160 238.780 -67.660 239.010 ;
        RECT -66.085 238.780 -65.585 239.010 ;
        RECT -68.160 238.290 -67.660 238.520 ;
        RECT -66.085 238.290 -65.585 238.520 ;
        RECT -68.160 237.800 -67.660 238.030 ;
        RECT -66.085 237.800 -65.585 238.030 ;
        RECT -68.160 237.310 -67.660 237.540 ;
        RECT -66.755 237.070 -66.455 237.545 ;
        RECT -66.085 237.310 -65.585 237.540 ;
        RECT -64.030 237.070 -63.790 241.320 ;
        RECT -63.295 240.850 -62.795 241.080 ;
        RECT -62.230 240.865 -61.860 241.710 ;
        RECT -61.220 241.340 -60.720 241.570 ;
        RECT -63.045 239.755 -62.545 239.985 ;
        RECT -63.045 238.775 -62.545 239.005 ;
        RECT -63.045 237.795 -62.545 238.025 ;
        RECT -66.760 236.865 -63.790 237.070 ;
        RECT -62.195 237.005 -61.910 240.865 ;
        RECT -61.220 240.850 -60.720 241.080 ;
        RECT -51.095 240.845 -50.645 250.310 ;
        RECT -49.540 243.095 -48.560 252.665 ;
        RECT -38.525 243.785 -37.770 247.920 ;
        RECT -35.980 243.805 -35.205 291.265 ;
        RECT -30.595 244.060 -29.890 246.885 ;
        RECT -36.305 242.470 -34.815 243.805 ;
        RECT -30.595 242.635 -29.895 244.060 ;
        RECT -26.495 243.930 -25.250 333.920 ;
        RECT -24.465 245.340 -23.140 376.245 ;
        RECT -22.065 247.300 -20.935 420.565 ;
        RECT -39.820 240.845 -39.000 240.865 ;
        RECT -19.280 240.845 -18.175 466.535 ;
        RECT -51.095 240.395 -18.175 240.845 ;
        RECT -39.820 240.375 -39.000 240.395 ;
        RECT -61.645 239.755 -60.645 239.985 ;
        RECT -61.645 238.775 -60.645 239.005 ;
        RECT -61.645 237.795 -60.645 238.025 ;
        RECT -66.755 236.860 -66.455 236.865 ;
        RECT -62.195 236.720 -60.735 237.005 ;
        RECT -50.025 236.490 -47.900 236.885 ;
        RECT -16.485 236.490 -15.600 510.300 ;
        RECT -62.820 235.895 -62.160 235.900 ;
        RECT -66.890 235.600 -62.160 235.895 ;
        RECT -66.890 235.595 -62.595 235.600 ;
        RECT -66.860 235.180 -66.560 235.595 ;
        RECT -63.045 234.970 -62.545 235.200 ;
        RECT -61.645 234.970 -60.645 235.200 ;
        RECT -50.025 234.835 -15.600 236.490 ;
        RECT -68.235 234.480 -67.235 234.710 ;
        RECT -66.335 234.480 -65.835 234.710 ;
        RECT -50.025 234.315 -47.900 234.835 ;
        RECT -63.045 233.990 -62.545 234.220 ;
        RECT -61.645 233.990 -60.645 234.220 ;
        RECT -68.235 233.500 -67.235 233.730 ;
        RECT -66.335 233.500 -65.835 233.730 ;
        RECT -63.045 233.010 -62.545 233.240 ;
        RECT -61.645 233.010 -60.645 233.240 ;
        RECT -55.300 233.155 -54.150 233.260 ;
        RECT -14.235 233.155 -12.680 555.970 ;
        RECT -68.235 232.520 -67.235 232.750 ;
        RECT -66.335 232.520 -65.835 232.750 ;
        RECT -55.300 231.900 -12.680 233.155 ;
        RECT -55.300 231.820 -54.150 231.900 ;
        RECT -68.145 231.315 -66.685 231.600 ;
        RECT -68.235 230.295 -67.235 230.525 ;
        RECT -68.235 229.315 -67.235 229.545 ;
        RECT -68.235 228.335 -67.235 228.565 ;
        RECT -68.160 227.240 -67.660 227.470 ;
        RECT -66.970 227.455 -66.685 231.315 ;
        RECT -63.295 230.995 -62.795 231.010 ;
        RECT -64.010 230.765 -62.795 230.995 ;
        RECT -61.220 230.780 -60.720 231.010 ;
        RECT -66.335 230.295 -65.835 230.525 ;
        RECT -64.010 230.020 -63.780 230.765 ;
        RECT -63.295 230.290 -62.795 230.520 ;
        RECT -61.220 230.290 -60.720 230.520 ;
        RECT -63.295 230.020 -62.795 230.030 ;
        RECT -64.010 229.810 -62.795 230.020 ;
        RECT -66.335 229.315 -65.835 229.545 ;
        RECT -64.010 229.045 -63.780 229.810 ;
        RECT -63.295 229.800 -62.795 229.810 ;
        RECT -61.220 229.800 -60.720 230.030 ;
        RECT -63.295 229.310 -62.795 229.540 ;
        RECT -61.220 229.310 -60.720 229.540 ;
        RECT -63.295 229.045 -62.795 229.050 ;
        RECT -64.010 228.835 -62.795 229.045 ;
        RECT -66.335 228.335 -65.835 228.565 ;
        RECT -64.010 228.065 -63.780 228.835 ;
        RECT -63.295 228.820 -62.795 228.835 ;
        RECT -61.220 228.820 -60.720 229.050 ;
        RECT -63.295 228.330 -62.795 228.560 ;
        RECT -61.220 228.330 -60.720 228.560 ;
        RECT -54.405 228.285 -52.700 228.565 ;
        RECT -9.570 228.285 -8.150 603.625 ;
        RECT -63.295 228.065 -62.795 228.070 ;
        RECT -64.010 227.855 -62.795 228.065 ;
        RECT -68.160 226.750 -67.660 226.980 ;
        RECT -67.020 226.610 -66.650 227.455 ;
        RECT -66.085 227.240 -65.585 227.470 ;
        RECT -64.010 227.425 -63.780 227.855 ;
        RECT -63.295 227.840 -62.795 227.855 ;
        RECT -65.070 227.195 -63.780 227.425 ;
        RECT -63.295 227.350 -62.795 227.580 ;
        RECT -62.230 227.365 -61.860 228.210 ;
        RECT -61.220 227.840 -60.720 228.070 ;
        RECT -66.085 226.750 -65.585 226.980 ;
        RECT -68.160 226.260 -67.660 226.490 ;
        RECT -66.085 226.260 -65.585 226.490 ;
        RECT -68.160 225.770 -67.660 226.000 ;
        RECT -66.085 225.770 -65.585 226.000 ;
        RECT -68.160 225.280 -67.660 225.510 ;
        RECT -66.085 225.280 -65.585 225.510 ;
        RECT -68.160 224.790 -67.660 225.020 ;
        RECT -66.085 224.790 -65.585 225.020 ;
        RECT -68.160 224.300 -67.660 224.530 ;
        RECT -66.085 224.300 -65.585 224.530 ;
        RECT -68.160 223.810 -67.660 224.040 ;
        RECT -66.745 223.560 -66.445 224.100 ;
        RECT -66.085 223.810 -65.585 224.040 ;
        RECT -65.070 223.560 -64.840 227.195 ;
        RECT -63.045 226.255 -62.545 226.485 ;
        RECT -63.045 225.275 -62.545 225.505 ;
        RECT -63.045 224.295 -62.545 224.525 ;
        RECT -66.745 223.370 -64.840 223.560 ;
        RECT -62.195 223.505 -61.910 227.365 ;
        RECT -61.220 227.350 -60.720 227.580 ;
        RECT -54.405 226.940 -8.150 228.285 ;
        RECT -54.405 226.635 -52.700 226.940 ;
        RECT -61.645 226.255 -60.645 226.485 ;
        RECT -61.645 225.275 -60.645 225.505 ;
        RECT -61.645 224.295 -60.645 224.525 ;
        RECT -66.745 223.330 -64.845 223.370 ;
        RECT -64.665 223.220 -60.735 223.505 ;
        RECT -64.665 222.460 -64.380 223.220 ;
        RECT -65.555 222.175 -64.380 222.460 ;
        RECT -64.140 222.805 -63.840 222.970 ;
        RECT -62.700 222.805 -62.040 222.815 ;
        RECT -64.140 222.515 -62.040 222.805 ;
        RECT -64.140 222.310 -63.840 222.515 ;
        RECT -65.555 218.620 -65.270 222.175 ;
        RECT -63.045 221.845 -62.545 222.075 ;
        RECT -61.645 221.845 -60.645 222.075 ;
        RECT -63.045 220.865 -62.545 221.095 ;
        RECT -61.645 220.865 -60.645 221.095 ;
        RECT -63.045 219.885 -62.545 220.115 ;
        RECT -61.645 219.885 -60.645 220.115 ;
        RECT -84.505 217.620 -34.990 218.620 ;
        RECT -67.410 214.410 -27.000 214.550 ;
        RECT -67.410 203.895 -67.270 214.410 ;
        RECT -63.895 213.725 -30.515 213.770 ;
        RECT -63.895 213.630 -29.930 213.725 ;
        RECT -67.470 203.200 -67.200 203.895 ;
        RECT -69.050 202.755 -68.050 202.985 ;
        RECT -69.050 201.210 -68.050 201.440 ;
        RECT -67.410 200.820 -67.270 203.200 ;
        RECT -67.130 202.265 -66.900 202.945 ;
        RECT -66.020 202.755 -65.020 202.985 ;
        RECT -67.500 200.125 -67.230 200.820 ;
        RECT -69.050 199.660 -68.050 199.890 ;
        RECT -69.050 198.680 -68.050 198.910 ;
        RECT -67.085 198.775 -66.945 202.265 ;
        RECT -66.410 200.735 -66.180 201.390 ;
        RECT -66.020 201.210 -65.020 201.440 ;
        RECT -67.130 198.080 -66.860 198.775 ;
        RECT -69.050 196.870 -68.050 197.100 ;
        RECT -69.050 196.380 -68.050 196.610 ;
        RECT -69.050 195.890 -68.050 196.120 ;
        RECT -66.350 196.105 -66.210 200.735 ;
        RECT -66.020 200.150 -65.020 200.380 ;
        RECT -66.020 199.660 -65.020 199.890 ;
        RECT -66.020 198.680 -65.020 198.910 ;
        RECT -66.020 198.190 -65.020 198.420 ;
        RECT -66.020 196.870 -65.020 197.100 ;
        RECT -67.215 195.965 -66.210 196.105 ;
        RECT -69.050 195.290 -68.050 195.520 ;
        RECT -67.215 195.030 -67.075 195.965 ;
        RECT -69.050 194.800 -68.050 195.030 ;
        RECT -69.050 194.310 -68.050 194.540 ;
        RECT -67.280 194.335 -67.010 195.030 ;
        RECT -66.020 194.800 -65.020 195.030 ;
        RECT -63.895 193.765 -63.755 213.630 ;
        RECT -39.705 213.005 -39.040 213.065 ;
        RECT -67.410 193.625 -63.755 193.765 ;
        RECT -63.230 212.815 -31.180 213.005 ;
        RECT -63.230 208.990 -63.040 212.815 ;
        RECT -50.815 212.245 -50.225 212.325 ;
        RECT -62.545 212.105 -31.865 212.245 ;
        RECT -63.230 205.590 -63.090 208.990 ;
        RECT -67.410 188.895 -67.270 193.625 ;
        RECT -65.845 192.945 -65.165 192.950 ;
        RECT -63.685 192.945 -63.455 193.140 ;
        RECT -65.845 192.725 -63.455 192.945 ;
        RECT -65.845 192.720 -65.165 192.725 ;
        RECT -63.685 192.460 -63.455 192.725 ;
        RECT -67.470 188.200 -67.200 188.895 ;
        RECT -69.050 187.755 -68.050 187.985 ;
        RECT -69.050 186.210 -68.050 186.440 ;
        RECT -67.410 185.820 -67.270 188.200 ;
        RECT -67.130 187.265 -66.900 187.945 ;
        RECT -66.020 187.755 -65.020 187.985 ;
        RECT -67.500 185.125 -67.230 185.820 ;
        RECT -69.050 184.660 -68.050 184.890 ;
        RECT -69.050 183.680 -68.050 183.910 ;
        RECT -67.085 183.775 -66.945 187.265 ;
        RECT -66.410 185.735 -66.180 186.390 ;
        RECT -66.020 186.210 -65.020 186.440 ;
        RECT -67.130 183.080 -66.860 183.775 ;
        RECT -69.050 181.870 -68.050 182.100 ;
        RECT -69.050 181.380 -68.050 181.610 ;
        RECT -69.050 180.890 -68.050 181.120 ;
        RECT -66.350 181.105 -66.210 185.735 ;
        RECT -66.020 185.150 -65.020 185.380 ;
        RECT -66.020 184.660 -65.020 184.890 ;
        RECT -66.020 183.680 -65.020 183.910 ;
        RECT -66.020 183.190 -65.020 183.420 ;
        RECT -66.020 181.870 -65.020 182.100 ;
        RECT -67.215 180.965 -66.210 181.105 ;
        RECT -69.050 180.290 -68.050 180.520 ;
        RECT -67.215 180.030 -67.075 180.965 ;
        RECT -69.050 179.800 -68.050 180.030 ;
        RECT -69.050 179.310 -68.050 179.540 ;
        RECT -67.280 179.335 -67.010 180.030 ;
        RECT -66.020 179.800 -65.020 180.030 ;
        RECT -65.845 178.420 -65.165 178.425 ;
        RECT -63.605 178.420 -63.375 178.615 ;
        RECT -65.845 178.200 -63.375 178.420 ;
        RECT -65.845 178.195 -65.165 178.200 ;
        RECT -63.605 177.935 -63.375 178.200 ;
        RECT -63.230 177.240 -63.040 205.590 ;
        RECT -67.410 177.100 -63.040 177.240 ;
        RECT -67.410 176.395 -67.270 177.100 ;
        RECT -67.470 175.700 -67.200 176.395 ;
        RECT -69.050 175.255 -68.050 175.485 ;
        RECT -69.050 173.710 -68.050 173.940 ;
        RECT -67.410 173.320 -67.270 175.700 ;
        RECT -67.130 174.765 -66.900 175.445 ;
        RECT -66.020 175.255 -65.020 175.485 ;
        RECT -67.500 172.625 -67.230 173.320 ;
        RECT -69.050 172.160 -68.050 172.390 ;
        RECT -69.050 171.180 -68.050 171.410 ;
        RECT -67.085 171.275 -66.945 174.765 ;
        RECT -66.410 173.235 -66.180 173.890 ;
        RECT -66.020 173.710 -65.020 173.940 ;
        RECT -67.130 170.580 -66.860 171.275 ;
        RECT -69.050 169.370 -68.050 169.600 ;
        RECT -69.050 168.880 -68.050 169.110 ;
        RECT -69.050 168.390 -68.050 168.620 ;
        RECT -66.350 168.605 -66.210 173.235 ;
        RECT -66.020 172.650 -65.020 172.880 ;
        RECT -66.020 172.160 -65.020 172.390 ;
        RECT -66.020 171.180 -65.020 171.410 ;
        RECT -66.020 170.690 -65.020 170.920 ;
        RECT -66.020 169.370 -65.020 169.600 ;
        RECT -67.215 168.465 -66.210 168.605 ;
        RECT -69.050 167.790 -68.050 168.020 ;
        RECT -67.215 167.530 -67.075 168.465 ;
        RECT -69.050 167.300 -68.050 167.530 ;
        RECT -69.050 166.810 -68.050 167.040 ;
        RECT -67.280 166.835 -67.010 167.530 ;
        RECT -66.020 167.300 -65.020 167.530 ;
        RECT -63.920 167.020 -63.690 167.700 ;
        RECT -65.845 166.335 -65.165 166.340 ;
        RECT -63.915 166.335 -63.695 167.020 ;
        RECT -65.845 166.115 -63.695 166.335 ;
        RECT -65.845 166.110 -65.165 166.115 ;
        RECT -62.545 164.865 -62.405 212.105 ;
        RECT -50.815 212.005 -50.225 212.105 ;
        RECT -56.480 211.450 -55.785 211.510 ;
        RECT -61.915 211.195 -32.430 211.450 ;
        RECT -61.915 209.515 -61.725 211.195 ;
        RECT -56.480 211.165 -55.785 211.195 ;
        RECT -52.300 210.670 -51.825 210.695 ;
        RECT -61.880 208.550 -61.725 209.515 ;
        RECT -61.205 210.415 -33.180 210.670 ;
        RECT -61.205 208.550 -60.975 210.415 ;
        RECT -52.300 210.400 -51.825 210.415 ;
        RECT -38.370 208.880 -37.925 208.995 ;
        RECT -67.410 164.725 -62.405 164.865 ;
        RECT -67.410 163.895 -67.270 164.725 ;
        RECT -67.470 163.200 -67.200 163.895 ;
        RECT -69.050 162.755 -68.050 162.985 ;
        RECT -69.050 161.210 -68.050 161.440 ;
        RECT -67.410 160.820 -67.270 163.200 ;
        RECT -67.130 162.265 -66.900 162.945 ;
        RECT -66.020 162.755 -65.020 162.985 ;
        RECT -67.500 160.125 -67.230 160.820 ;
        RECT -69.050 159.660 -68.050 159.890 ;
        RECT -69.050 158.680 -68.050 158.910 ;
        RECT -67.085 158.775 -66.945 162.265 ;
        RECT -66.410 160.735 -66.180 161.390 ;
        RECT -66.020 161.210 -65.020 161.440 ;
        RECT -67.130 158.080 -66.860 158.775 ;
        RECT -69.050 156.870 -68.050 157.100 ;
        RECT -69.050 156.380 -68.050 156.610 ;
        RECT -69.050 155.890 -68.050 156.120 ;
        RECT -66.350 156.105 -66.210 160.735 ;
        RECT -66.020 160.150 -65.020 160.380 ;
        RECT -66.020 159.660 -65.020 159.890 ;
        RECT -66.020 158.680 -65.020 158.910 ;
        RECT -66.020 158.190 -65.020 158.420 ;
        RECT -66.020 156.870 -65.020 157.100 ;
        RECT -67.215 155.965 -66.210 156.105 ;
        RECT -69.050 155.290 -68.050 155.520 ;
        RECT -67.215 155.030 -67.075 155.965 ;
        RECT -69.050 154.800 -68.050 155.030 ;
        RECT -69.050 154.310 -68.050 154.540 ;
        RECT -67.280 154.335 -67.010 155.030 ;
        RECT -66.020 154.800 -65.020 155.030 ;
        RECT -63.985 154.535 -63.755 155.215 ;
        RECT -65.845 153.935 -65.165 153.940 ;
        RECT -63.980 153.935 -63.760 154.535 ;
        RECT -65.845 153.715 -63.760 153.935 ;
        RECT -65.845 153.710 -65.165 153.715 ;
        RECT -63.980 153.710 -63.760 153.715 ;
        RECT -61.980 152.505 -61.725 208.550 ;
        RECT -67.410 152.365 -61.725 152.505 ;
        RECT -67.410 151.395 -67.270 152.365 ;
        RECT -67.470 150.700 -67.200 151.395 ;
        RECT -69.050 150.255 -68.050 150.485 ;
        RECT -69.050 148.710 -68.050 148.940 ;
        RECT -67.410 148.320 -67.270 150.700 ;
        RECT -67.130 149.765 -66.900 150.445 ;
        RECT -66.020 150.255 -65.020 150.485 ;
        RECT -67.500 147.625 -67.230 148.320 ;
        RECT -69.050 147.160 -68.050 147.390 ;
        RECT -69.050 146.180 -68.050 146.410 ;
        RECT -67.085 146.275 -66.945 149.765 ;
        RECT -66.410 148.235 -66.180 148.890 ;
        RECT -66.020 148.710 -65.020 148.940 ;
        RECT -67.130 145.580 -66.860 146.275 ;
        RECT -69.050 144.370 -68.050 144.600 ;
        RECT -69.050 143.880 -68.050 144.110 ;
        RECT -69.050 143.390 -68.050 143.620 ;
        RECT -66.350 143.605 -66.210 148.235 ;
        RECT -66.020 147.650 -65.020 147.880 ;
        RECT -66.020 147.160 -65.020 147.390 ;
        RECT -66.020 146.180 -65.020 146.410 ;
        RECT -66.020 145.690 -65.020 145.920 ;
        RECT -66.020 144.370 -65.020 144.600 ;
        RECT -67.215 143.465 -66.210 143.605 ;
        RECT -69.050 142.790 -68.050 143.020 ;
        RECT -67.215 142.530 -67.075 143.465 ;
        RECT -69.050 142.300 -68.050 142.530 ;
        RECT -69.050 141.810 -68.050 142.040 ;
        RECT -67.280 141.835 -67.010 142.530 ;
        RECT -66.020 142.300 -65.020 142.530 ;
        RECT -65.865 141.195 -65.185 141.200 ;
        RECT -62.335 141.195 -61.655 141.200 ;
        RECT -65.865 140.975 -61.655 141.195 ;
        RECT -65.865 140.970 -65.185 140.975 ;
        RECT -62.335 140.970 -61.655 140.975 ;
        RECT -61.230 139.650 -60.975 208.550 ;
        RECT -56.190 208.740 -37.925 208.880 ;
        RECT -56.190 204.450 -56.050 208.740 ;
        RECT -38.370 207.905 -37.925 208.740 ;
        RECT -38.360 204.450 -38.220 207.905 ;
        RECT -56.190 203.945 -56.015 204.450 ;
        RECT -38.395 203.945 -38.220 204.450 ;
        RECT -56.215 203.250 -55.945 203.945 ;
        RECT -38.465 203.250 -38.195 203.945 ;
        RECT -57.795 202.805 -56.795 203.035 ;
        RECT -57.795 201.260 -56.795 201.490 ;
        RECT -56.155 200.870 -56.015 203.250 ;
        RECT -55.875 202.315 -55.645 202.995 ;
        RECT -54.765 202.805 -53.765 203.035 ;
        RECT -40.645 202.805 -39.645 203.035 ;
        RECT -38.765 202.315 -38.535 202.995 ;
        RECT -56.245 200.175 -55.975 200.870 ;
        RECT -57.795 199.710 -56.795 199.940 ;
        RECT -57.795 198.730 -56.795 198.960 ;
        RECT -55.830 198.825 -55.690 202.315 ;
        RECT -55.155 200.785 -54.925 201.440 ;
        RECT -54.765 201.260 -53.765 201.490 ;
        RECT -40.645 201.260 -39.645 201.490 ;
        RECT -39.485 200.785 -39.255 201.440 ;
        RECT -55.875 198.130 -55.605 198.825 ;
        RECT -57.795 196.920 -56.795 197.150 ;
        RECT -57.795 196.430 -56.795 196.660 ;
        RECT -57.795 195.940 -56.795 196.170 ;
        RECT -55.095 196.155 -54.955 200.785 ;
        RECT -54.765 200.200 -53.765 200.430 ;
        RECT -40.645 200.200 -39.645 200.430 ;
        RECT -54.765 199.710 -53.765 199.940 ;
        RECT -40.645 199.710 -39.645 199.940 ;
        RECT -54.765 198.730 -53.765 198.960 ;
        RECT -40.645 198.730 -39.645 198.960 ;
        RECT -54.765 198.240 -53.765 198.470 ;
        RECT -40.645 198.240 -39.645 198.470 ;
        RECT -54.765 196.920 -53.765 197.150 ;
        RECT -40.645 196.920 -39.645 197.150 ;
        RECT -55.960 196.015 -54.955 196.155 ;
        RECT -39.455 196.155 -39.315 200.785 ;
        RECT -38.720 198.825 -38.580 202.315 ;
        RECT -38.395 200.870 -38.255 203.250 ;
        RECT -37.615 202.805 -36.615 203.035 ;
        RECT -37.615 201.260 -36.615 201.490 ;
        RECT -38.435 200.175 -38.165 200.870 ;
        RECT -37.615 199.710 -36.615 199.940 ;
        RECT -38.805 198.130 -38.535 198.825 ;
        RECT -37.615 198.730 -36.615 198.960 ;
        RECT -37.615 196.920 -36.615 197.150 ;
        RECT -37.615 196.430 -36.615 196.660 ;
        RECT -39.455 196.015 -38.450 196.155 ;
        RECT -57.795 195.340 -56.795 195.570 ;
        RECT -55.960 195.080 -55.820 196.015 ;
        RECT -38.590 195.080 -38.450 196.015 ;
        RECT -37.615 195.940 -36.615 196.170 ;
        RECT -37.615 195.340 -36.615 195.570 ;
        RECT -57.795 194.850 -56.410 195.080 ;
        RECT -57.795 194.360 -56.795 194.590 ;
        RECT -56.640 193.020 -56.410 194.850 ;
        RECT -56.025 194.385 -55.755 195.080 ;
        RECT -54.765 194.850 -53.765 195.080 ;
        RECT -40.645 194.850 -39.645 195.080 ;
        RECT -38.655 194.385 -38.385 195.080 ;
        RECT -38.000 194.850 -36.615 195.080 ;
        RECT -38.000 193.020 -37.770 194.850 ;
        RECT -37.615 194.360 -36.615 194.590 ;
        RECT -56.640 192.340 -56.365 193.020 ;
        RECT -54.815 192.435 -53.315 192.665 ;
        RECT -41.095 192.435 -39.595 192.665 ;
        RECT -38.045 192.340 -37.770 193.020 ;
        RECT -56.640 192.320 -56.410 192.340 ;
        RECT -38.000 192.320 -37.770 192.340 ;
        RECT -57.850 191.945 -56.850 192.175 ;
        RECT -37.560 191.945 -36.560 192.175 ;
        RECT -54.815 191.455 -53.315 191.685 ;
        RECT -41.095 191.455 -39.595 191.685 ;
        RECT -57.850 190.965 -56.850 191.195 ;
        RECT -54.810 190.885 -53.310 191.115 ;
        RECT -41.100 190.885 -39.600 191.115 ;
        RECT -37.560 190.965 -36.560 191.195 ;
        RECT -54.810 190.395 -53.310 190.625 ;
        RECT -41.100 190.395 -39.600 190.625 ;
        RECT -57.850 189.985 -56.850 190.215 ;
        RECT -54.810 189.905 -53.310 190.135 ;
        RECT -41.100 189.905 -39.600 190.135 ;
        RECT -37.560 189.985 -36.560 190.215 ;
        RECT -54.810 189.340 -53.310 189.570 ;
        RECT -41.100 189.340 -39.600 189.570 ;
        RECT -54.810 188.850 -53.310 189.080 ;
        RECT -41.100 188.850 -39.600 189.080 ;
        RECT -54.810 188.360 -53.310 188.590 ;
        RECT -41.100 188.360 -39.600 188.590 ;
        RECT -57.850 186.295 -56.850 186.525 ;
        RECT -54.310 186.295 -53.310 186.525 ;
        RECT -41.100 186.295 -40.100 186.525 ;
        RECT -37.560 186.295 -36.560 186.525 ;
        RECT -53.545 183.900 -53.125 183.905 ;
        RECT -55.040 183.670 -53.125 183.900 ;
        RECT -57.725 183.180 -56.225 183.410 ;
        RECT -53.360 182.920 -53.125 183.670 ;
        RECT -55.040 182.690 -53.125 182.920 ;
        RECT -57.725 182.200 -53.540 182.430 ;
        RECT -53.360 181.940 -53.125 182.690 ;
        RECT -55.040 181.710 -53.125 181.940 ;
        RECT -57.730 180.135 -56.720 180.365 ;
        RECT -56.950 179.875 -56.720 180.135 ;
        RECT -56.960 179.645 -56.075 179.875 ;
        RECT -56.960 179.385 -56.720 179.645 ;
        RECT -57.730 179.155 -56.720 179.385 ;
        RECT -56.960 178.895 -56.720 179.155 ;
        RECT -56.960 178.665 -56.075 178.895 ;
        RECT -56.950 178.405 -56.720 178.665 ;
        RECT -57.730 178.175 -56.720 178.405 ;
        RECT -56.950 178.050 -56.720 178.175 ;
        RECT -60.400 176.230 -60.170 176.910 ;
        RECT -60.380 141.665 -60.170 176.230 ;
        RECT -59.980 175.710 -59.750 176.485 ;
        RECT -53.555 175.875 -53.135 175.880 ;
        RECT -60.390 140.985 -60.160 141.665 ;
        RECT -67.410 139.510 -60.975 139.650 ;
        RECT -67.410 138.895 -67.270 139.510 ;
        RECT -67.470 138.200 -67.200 138.895 ;
        RECT -69.050 137.755 -68.050 137.985 ;
        RECT -69.050 136.210 -68.050 136.440 ;
        RECT -67.410 135.820 -67.270 138.200 ;
        RECT -67.130 137.265 -66.900 137.945 ;
        RECT -66.020 137.755 -65.020 137.985 ;
        RECT -67.500 135.125 -67.230 135.820 ;
        RECT -69.050 134.660 -68.050 134.890 ;
        RECT -69.050 133.680 -68.050 133.910 ;
        RECT -67.085 133.775 -66.945 137.265 ;
        RECT -66.410 135.735 -66.180 136.390 ;
        RECT -66.020 136.210 -65.020 136.440 ;
        RECT -67.130 133.080 -66.860 133.775 ;
        RECT -69.050 131.870 -68.050 132.100 ;
        RECT -69.050 131.380 -68.050 131.610 ;
        RECT -69.050 130.890 -68.050 131.120 ;
        RECT -66.350 131.105 -66.210 135.735 ;
        RECT -66.020 135.150 -65.020 135.380 ;
        RECT -66.020 134.660 -65.020 134.890 ;
        RECT -66.020 133.680 -65.020 133.910 ;
        RECT -66.020 133.190 -65.020 133.420 ;
        RECT -66.020 131.870 -65.020 132.100 ;
        RECT -67.215 130.965 -66.210 131.105 ;
        RECT -69.050 130.290 -68.050 130.520 ;
        RECT -67.215 130.030 -67.075 130.965 ;
        RECT -69.050 129.800 -68.050 130.030 ;
        RECT -69.050 129.310 -68.050 129.540 ;
        RECT -67.280 129.335 -67.010 130.030 ;
        RECT -66.020 129.800 -65.020 130.030 ;
        RECT -59.970 129.265 -59.760 175.710 ;
        RECT -55.050 175.645 -53.135 175.875 ;
        RECT -57.735 175.155 -56.235 175.385 ;
        RECT -53.370 174.895 -53.135 175.645 ;
        RECT -55.050 174.665 -53.135 174.895 ;
        RECT -57.735 174.175 -53.550 174.405 ;
        RECT -53.370 173.915 -53.135 174.665 ;
        RECT -55.050 173.685 -53.135 173.915 ;
        RECT -57.740 172.110 -56.730 172.340 ;
        RECT -56.960 171.850 -56.730 172.110 ;
        RECT -56.970 171.620 -56.085 171.850 ;
        RECT -56.970 171.360 -56.730 171.620 ;
        RECT -57.740 171.130 -56.730 171.360 ;
        RECT -56.970 170.870 -56.730 171.130 ;
        RECT -56.970 170.640 -56.085 170.870 ;
        RECT -56.960 170.380 -56.730 170.640 ;
        RECT -57.740 170.150 -56.730 170.380 ;
        RECT -56.960 170.025 -56.730 170.150 ;
        RECT -56.140 169.220 -55.910 169.350 ;
        RECT -52.865 169.220 -52.635 177.735 ;
        RECT -56.140 168.990 -52.635 169.220 ;
        RECT -56.140 168.670 -55.910 168.990 ;
        RECT -57.010 168.455 -56.330 168.495 ;
        RECT -52.305 168.455 -52.075 185.575 ;
        RECT -57.010 168.265 -52.075 168.455 ;
        RECT -57.000 168.225 -52.075 168.265 ;
        RECT -42.335 168.455 -42.105 185.575 ;
        RECT -41.285 183.900 -40.865 183.905 ;
        RECT -41.285 183.670 -39.370 183.900 ;
        RECT -41.285 182.920 -41.050 183.670 ;
        RECT -38.185 183.180 -36.685 183.410 ;
        RECT -41.285 182.690 -39.370 182.920 ;
        RECT -41.285 181.940 -41.050 182.690 ;
        RECT -40.870 182.200 -36.685 182.430 ;
        RECT -41.285 181.710 -39.370 181.940 ;
        RECT -37.690 180.135 -36.680 180.365 ;
        RECT -37.690 179.875 -37.460 180.135 ;
        RECT -38.335 179.645 -37.450 179.875 ;
        RECT -37.690 179.385 -37.450 179.645 ;
        RECT -37.690 179.155 -36.680 179.385 ;
        RECT -37.690 178.895 -37.450 179.155 ;
        RECT -38.335 178.665 -37.450 178.895 ;
        RECT -37.690 178.405 -37.460 178.665 ;
        RECT -37.690 178.175 -36.680 178.405 ;
        RECT -37.690 178.050 -37.460 178.175 ;
        RECT -41.775 169.220 -41.545 177.735 ;
        RECT -41.275 175.875 -40.855 175.880 ;
        RECT -41.275 175.645 -39.360 175.875 ;
        RECT -34.660 175.710 -34.430 176.485 ;
        RECT -34.240 176.230 -34.010 176.910 ;
        RECT -41.275 174.895 -41.040 175.645 ;
        RECT -38.175 175.155 -36.675 175.385 ;
        RECT -41.275 174.665 -39.360 174.895 ;
        RECT -41.275 173.915 -41.040 174.665 ;
        RECT -40.860 174.175 -36.675 174.405 ;
        RECT -41.275 173.685 -39.360 173.915 ;
        RECT -37.680 172.110 -36.670 172.340 ;
        RECT -37.680 171.850 -37.450 172.110 ;
        RECT -38.325 171.620 -37.440 171.850 ;
        RECT -37.680 171.360 -37.440 171.620 ;
        RECT -37.680 171.130 -36.670 171.360 ;
        RECT -37.680 170.870 -37.440 171.130 ;
        RECT -38.325 170.640 -37.440 170.870 ;
        RECT -37.680 170.380 -37.450 170.640 ;
        RECT -37.680 170.150 -36.670 170.380 ;
        RECT -37.680 170.025 -37.450 170.150 ;
        RECT -38.500 169.220 -38.270 169.350 ;
        RECT -41.775 168.990 -38.270 169.220 ;
        RECT -38.500 168.670 -38.270 168.990 ;
        RECT -38.080 168.455 -37.400 168.495 ;
        RECT -42.335 168.265 -37.400 168.455 ;
        RECT -42.335 168.225 -37.410 168.265 ;
        RECT -54.770 167.625 -53.270 167.855 ;
        RECT -41.140 167.625 -39.640 167.855 ;
        RECT -57.805 167.135 -56.805 167.365 ;
        RECT -37.605 167.135 -36.605 167.365 ;
        RECT -54.770 166.645 -53.270 166.875 ;
        RECT -41.140 166.645 -39.640 166.875 ;
        RECT -57.805 166.155 -56.805 166.385 ;
        RECT -54.765 166.075 -53.265 166.305 ;
        RECT -41.145 166.075 -39.645 166.305 ;
        RECT -37.605 166.155 -36.605 166.385 ;
        RECT -54.765 165.585 -53.265 165.815 ;
        RECT -41.145 165.585 -39.645 165.815 ;
        RECT -57.805 165.175 -56.805 165.405 ;
        RECT -54.765 165.095 -53.265 165.325 ;
        RECT -41.145 165.095 -39.645 165.325 ;
        RECT -37.605 165.175 -36.605 165.405 ;
        RECT -54.765 164.530 -53.265 164.760 ;
        RECT -41.145 164.530 -39.645 164.760 ;
        RECT -54.765 164.040 -53.265 164.270 ;
        RECT -41.145 164.040 -39.645 164.270 ;
        RECT -54.765 163.550 -53.265 163.780 ;
        RECT -41.145 163.550 -39.645 163.780 ;
        RECT -57.805 161.485 -56.805 161.715 ;
        RECT -54.265 161.485 -53.265 161.715 ;
        RECT -41.145 161.485 -40.145 161.715 ;
        RECT -37.605 161.485 -36.605 161.715 ;
        RECT -55.775 161.045 -55.510 161.465 ;
        RECT -38.900 161.045 -38.635 161.465 ;
        RECT -55.775 160.760 -52.980 161.045 ;
        RECT -57.890 158.795 -56.890 159.025 ;
        RECT -55.990 158.795 -55.490 159.025 ;
        RECT -57.890 157.815 -56.890 158.045 ;
        RECT -55.990 157.815 -55.490 158.045 ;
        RECT -57.890 156.835 -56.890 157.065 ;
        RECT -55.990 156.835 -55.490 157.065 ;
        RECT -53.265 156.735 -52.980 160.760 ;
        RECT -54.695 156.395 -54.395 156.600 ;
        RECT -56.495 156.105 -54.395 156.395 ;
        RECT -56.495 156.095 -55.835 156.105 ;
        RECT -54.695 155.940 -54.395 156.105 ;
        RECT -54.155 156.450 -52.980 156.735 ;
        RECT -41.430 160.760 -38.635 161.045 ;
        RECT -41.430 156.735 -41.145 160.760 ;
        RECT -38.920 158.795 -38.420 159.025 ;
        RECT -37.520 158.795 -36.520 159.025 ;
        RECT -38.920 157.815 -38.420 158.045 ;
        RECT -37.520 157.815 -36.520 158.045 ;
        RECT -40.450 157.300 -40.150 157.650 ;
        RECT -40.450 157.010 -39.715 157.300 ;
        RECT -40.450 156.990 -40.150 157.010 ;
        RECT -41.430 156.450 -40.255 156.735 ;
        RECT -54.155 155.690 -53.870 156.450 ;
        RECT -57.800 155.405 -53.870 155.690 ;
        RECT -40.540 155.690 -40.255 156.450 ;
        RECT -40.005 156.395 -39.715 157.010 ;
        RECT -38.920 156.835 -38.420 157.065 ;
        RECT -37.520 156.835 -36.520 157.065 ;
        RECT -40.005 156.105 -37.915 156.395 ;
        RECT -38.575 156.095 -37.915 156.105 ;
        RECT -53.690 155.540 -51.790 155.580 ;
        RECT -57.890 154.385 -56.890 154.615 ;
        RECT -57.890 153.405 -56.890 153.635 ;
        RECT -57.890 152.425 -56.890 152.655 ;
        RECT -57.815 151.330 -57.315 151.560 ;
        RECT -56.625 151.545 -56.340 155.405 ;
        RECT -53.695 155.350 -51.790 155.540 ;
        RECT -55.990 154.385 -55.490 154.615 ;
        RECT -55.990 153.405 -55.490 153.635 ;
        RECT -55.990 152.425 -55.490 152.655 ;
        RECT -53.695 151.715 -53.465 155.350 ;
        RECT -52.950 154.870 -52.450 155.100 ;
        RECT -52.090 154.810 -51.790 155.350 ;
        RECT -42.620 155.540 -40.720 155.580 ;
        RECT -42.620 155.350 -40.715 155.540 ;
        RECT -40.540 155.405 -36.610 155.690 ;
        RECT -50.875 154.870 -50.375 155.100 ;
        RECT -44.035 154.870 -43.535 155.100 ;
        RECT -42.620 154.810 -42.320 155.350 ;
        RECT -41.960 154.870 -41.460 155.100 ;
        RECT -52.950 154.380 -52.450 154.610 ;
        RECT -50.875 154.380 -50.375 154.610 ;
        RECT -44.035 154.380 -43.535 154.610 ;
        RECT -41.960 154.380 -41.460 154.610 ;
        RECT -52.950 153.890 -52.450 154.120 ;
        RECT -50.875 153.890 -50.375 154.120 ;
        RECT -44.035 153.890 -43.535 154.120 ;
        RECT -41.960 153.890 -41.460 154.120 ;
        RECT -52.950 153.400 -52.450 153.630 ;
        RECT -50.875 153.400 -50.375 153.630 ;
        RECT -44.035 153.400 -43.535 153.630 ;
        RECT -41.960 153.400 -41.460 153.630 ;
        RECT -52.950 152.910 -52.450 153.140 ;
        RECT -50.875 152.910 -50.375 153.140 ;
        RECT -44.035 152.910 -43.535 153.140 ;
        RECT -41.960 152.910 -41.460 153.140 ;
        RECT -52.950 152.420 -52.450 152.650 ;
        RECT -50.875 152.420 -50.375 152.650 ;
        RECT -44.035 152.420 -43.535 152.650 ;
        RECT -41.960 152.420 -41.460 152.650 ;
        RECT -52.950 151.930 -52.450 152.160 ;
        RECT -57.815 150.840 -57.315 151.070 ;
        RECT -56.675 150.700 -56.305 151.545 ;
        RECT -55.740 151.330 -55.240 151.560 ;
        RECT -54.755 151.485 -53.465 151.715 ;
        RECT -55.740 151.055 -55.240 151.070 ;
        RECT -54.755 151.055 -54.525 151.485 ;
        RECT -52.950 151.440 -52.450 151.670 ;
        RECT -51.885 151.455 -51.515 152.300 ;
        RECT -50.875 151.930 -50.375 152.160 ;
        RECT -44.035 151.930 -43.535 152.160 ;
        RECT -55.740 150.845 -54.525 151.055 ;
        RECT -55.740 150.840 -55.240 150.845 ;
        RECT -57.815 150.350 -57.315 150.580 ;
        RECT -55.740 150.350 -55.240 150.580 ;
        RECT -57.815 149.860 -57.315 150.090 ;
        RECT -55.740 150.075 -55.240 150.090 ;
        RECT -54.755 150.075 -54.525 150.845 ;
        RECT -52.700 150.345 -52.200 150.575 ;
        RECT -55.740 149.865 -54.525 150.075 ;
        RECT -55.740 149.860 -55.240 149.865 ;
        RECT -57.815 149.370 -57.315 149.600 ;
        RECT -55.740 149.370 -55.240 149.600 ;
        RECT -57.815 148.880 -57.315 149.110 ;
        RECT -55.740 149.100 -55.240 149.110 ;
        RECT -54.755 149.100 -54.525 149.865 ;
        RECT -52.700 149.365 -52.200 149.595 ;
        RECT -55.740 148.890 -54.525 149.100 ;
        RECT -55.740 148.880 -55.240 148.890 ;
        RECT -57.815 148.390 -57.315 148.620 ;
        RECT -55.740 148.390 -55.240 148.620 ;
        RECT -54.755 148.145 -54.525 148.890 ;
        RECT -52.700 148.385 -52.200 148.615 ;
        RECT -57.815 147.900 -57.315 148.130 ;
        RECT -55.740 147.915 -54.525 148.145 ;
        RECT -55.740 147.900 -55.240 147.915 ;
        RECT -51.850 147.595 -51.565 151.455 ;
        RECT -50.875 151.440 -50.375 151.670 ;
        RECT -44.035 151.440 -43.535 151.670 ;
        RECT -42.895 151.455 -42.525 152.300 ;
        RECT -41.960 151.930 -41.460 152.160 ;
        RECT -40.945 151.715 -40.715 155.350 ;
        RECT -38.920 154.385 -38.420 154.615 ;
        RECT -38.920 153.405 -38.420 153.635 ;
        RECT -38.920 152.425 -38.420 152.655 ;
        RECT -51.300 150.345 -50.300 150.575 ;
        RECT -44.110 150.345 -43.110 150.575 ;
        RECT -51.300 149.365 -50.300 149.595 ;
        RECT -44.110 149.365 -43.110 149.595 ;
        RECT -51.300 148.385 -50.300 148.615 ;
        RECT -44.110 148.385 -43.110 148.615 ;
        RECT -42.845 147.595 -42.560 151.455 ;
        RECT -41.960 151.440 -41.460 151.670 ;
        RECT -40.945 151.485 -39.655 151.715 ;
        RECT -39.885 151.055 -39.655 151.485 ;
        RECT -39.170 151.330 -38.670 151.560 ;
        RECT -38.070 151.545 -37.785 155.405 ;
        RECT -37.520 154.385 -36.520 154.615 ;
        RECT -37.520 153.405 -36.520 153.635 ;
        RECT -37.520 152.425 -36.520 152.655 ;
        RECT -39.170 151.055 -38.670 151.070 ;
        RECT -39.885 150.845 -38.670 151.055 ;
        RECT -42.210 150.345 -41.710 150.575 ;
        RECT -39.885 150.075 -39.655 150.845 ;
        RECT -39.170 150.840 -38.670 150.845 ;
        RECT -38.105 150.700 -37.735 151.545 ;
        RECT -37.095 151.330 -36.595 151.560 ;
        RECT -37.095 150.840 -36.595 151.070 ;
        RECT -39.170 150.350 -38.670 150.580 ;
        RECT -37.095 150.350 -36.595 150.580 ;
        RECT -39.170 150.075 -38.670 150.090 ;
        RECT -39.885 149.865 -38.670 150.075 ;
        RECT -42.210 149.365 -41.710 149.595 ;
        RECT -39.885 149.100 -39.655 149.865 ;
        RECT -39.170 149.860 -38.670 149.865 ;
        RECT -37.095 149.860 -36.595 150.090 ;
        RECT -39.170 149.370 -38.670 149.600 ;
        RECT -37.095 149.370 -36.595 149.600 ;
        RECT -39.170 149.100 -38.670 149.110 ;
        RECT -39.885 148.890 -38.670 149.100 ;
        RECT -42.210 148.385 -41.710 148.615 ;
        RECT -39.885 148.145 -39.655 148.890 ;
        RECT -39.170 148.880 -38.670 148.890 ;
        RECT -37.095 148.880 -36.595 149.110 ;
        RECT -39.170 148.390 -38.670 148.620 ;
        RECT -37.095 148.390 -36.595 148.620 ;
        RECT -39.885 147.915 -38.670 148.145 ;
        RECT -39.170 147.900 -38.670 147.915 ;
        RECT -37.095 147.900 -36.595 148.130 ;
        RECT -51.850 147.310 -50.390 147.595 ;
        RECT -44.020 147.310 -42.560 147.595 ;
        RECT -40.445 147.365 -40.145 147.580 ;
        RECT -42.265 147.065 -40.145 147.365 ;
        RECT -40.445 146.920 -40.145 147.065 ;
        RECT -52.700 146.160 -52.200 146.390 ;
        RECT -51.300 146.160 -50.300 146.390 ;
        RECT -44.110 146.160 -43.110 146.390 ;
        RECT -42.210 146.160 -41.710 146.390 ;
        RECT -57.890 145.670 -56.890 145.900 ;
        RECT -55.990 145.670 -55.490 145.900 ;
        RECT -38.920 145.670 -38.420 145.900 ;
        RECT -37.520 145.670 -36.520 145.900 ;
        RECT -52.700 145.180 -52.200 145.410 ;
        RECT -51.300 145.180 -50.300 145.410 ;
        RECT -44.110 145.180 -43.110 145.410 ;
        RECT -42.210 145.180 -41.710 145.410 ;
        RECT -57.890 144.690 -56.890 144.920 ;
        RECT -55.990 144.690 -55.490 144.920 ;
        RECT -38.920 144.690 -38.420 144.920 ;
        RECT -37.520 144.690 -36.520 144.920 ;
        RECT -52.700 144.200 -52.200 144.430 ;
        RECT -51.300 144.200 -50.300 144.430 ;
        RECT -44.110 144.200 -43.110 144.430 ;
        RECT -42.210 144.200 -41.710 144.430 ;
        RECT -57.890 143.710 -56.890 143.940 ;
        RECT -55.990 143.710 -55.490 143.940 ;
        RECT -51.975 143.315 -51.675 143.730 ;
        RECT -42.735 143.315 -42.435 143.730 ;
        RECT -38.920 143.710 -38.420 143.940 ;
        RECT -37.520 143.710 -36.520 143.940 ;
        RECT -55.940 143.310 -51.645 143.315 ;
        RECT -56.375 143.015 -51.645 143.310 ;
        RECT -42.765 143.310 -38.470 143.315 ;
        RECT -42.765 143.015 -38.035 143.310 ;
        RECT -56.375 143.010 -55.715 143.015 ;
        RECT -38.695 143.010 -38.035 143.015 ;
        RECT -40.450 142.735 -40.150 142.875 ;
        RECT -40.450 142.435 -37.910 142.735 ;
        RECT -40.450 142.190 -40.150 142.435 ;
        RECT -57.800 141.905 -56.340 142.190 ;
        RECT -52.080 142.045 -51.780 142.050 ;
        RECT -42.630 142.045 -42.330 142.050 ;
        RECT -57.890 140.885 -56.890 141.115 ;
        RECT -57.890 139.905 -56.890 140.135 ;
        RECT -57.890 138.925 -56.890 139.155 ;
        RECT -57.815 137.830 -57.315 138.060 ;
        RECT -56.625 138.045 -56.340 141.905 ;
        RECT -54.745 141.840 -51.775 142.045 ;
        RECT -42.635 141.840 -39.665 142.045 ;
        RECT -55.990 140.885 -55.490 141.115 ;
        RECT -55.990 139.905 -55.490 140.135 ;
        RECT -55.990 138.925 -55.490 139.155 ;
        RECT -57.815 137.340 -57.315 137.570 ;
        RECT -56.675 137.200 -56.305 138.045 ;
        RECT -55.740 137.830 -55.240 138.060 ;
        RECT -54.745 137.590 -54.505 141.840 ;
        RECT -52.950 141.370 -52.450 141.600 ;
        RECT -52.080 141.365 -51.780 141.840 ;
        RECT -50.875 141.370 -50.375 141.600 ;
        RECT -44.035 141.370 -43.535 141.600 ;
        RECT -42.630 141.365 -42.330 141.840 ;
        RECT -41.960 141.370 -41.460 141.600 ;
        RECT -52.950 140.880 -52.450 141.110 ;
        RECT -50.875 140.880 -50.375 141.110 ;
        RECT -44.035 140.880 -43.535 141.110 ;
        RECT -41.960 140.880 -41.460 141.110 ;
        RECT -52.950 140.390 -52.450 140.620 ;
        RECT -50.875 140.390 -50.375 140.620 ;
        RECT -44.035 140.390 -43.535 140.620 ;
        RECT -41.960 140.390 -41.460 140.620 ;
        RECT -52.950 139.900 -52.450 140.130 ;
        RECT -50.875 139.900 -50.375 140.130 ;
        RECT -44.035 139.900 -43.535 140.130 ;
        RECT -41.960 139.900 -41.460 140.130 ;
        RECT -52.950 139.410 -52.450 139.640 ;
        RECT -50.875 139.410 -50.375 139.640 ;
        RECT -44.035 139.410 -43.535 139.640 ;
        RECT -41.960 139.410 -41.460 139.640 ;
        RECT -52.950 138.920 -52.450 139.150 ;
        RECT -50.875 138.920 -50.375 139.150 ;
        RECT -44.035 138.920 -43.535 139.150 ;
        RECT -41.960 138.920 -41.460 139.150 ;
        RECT -52.950 138.430 -52.450 138.660 ;
        RECT -52.950 137.940 -52.450 138.170 ;
        RECT -51.885 137.955 -51.515 138.800 ;
        RECT -50.875 138.430 -50.375 138.660 ;
        RECT -44.035 138.430 -43.535 138.660 ;
        RECT -55.335 137.570 -54.505 137.590 ;
        RECT -55.740 137.340 -54.505 137.570 ;
        RECT -55.335 137.285 -54.505 137.340 ;
        RECT -57.815 136.850 -57.315 137.080 ;
        RECT -55.740 136.850 -55.240 137.080 ;
        RECT -54.745 136.635 -54.505 137.285 ;
        RECT -52.700 136.845 -52.200 137.075 ;
        RECT -55.345 136.590 -54.505 136.635 ;
        RECT -57.815 136.360 -57.315 136.590 ;
        RECT -55.740 136.360 -54.505 136.590 ;
        RECT -55.345 136.330 -54.505 136.360 ;
        RECT -57.815 135.870 -57.315 136.100 ;
        RECT -55.740 135.870 -55.240 136.100 ;
        RECT -54.745 135.655 -54.505 136.330 ;
        RECT -52.700 135.865 -52.200 136.095 ;
        RECT -55.335 135.610 -54.505 135.655 ;
        RECT -57.815 135.380 -57.315 135.610 ;
        RECT -55.740 135.380 -54.505 135.610 ;
        RECT -55.335 135.350 -54.505 135.380 ;
        RECT -57.815 134.890 -57.315 135.120 ;
        RECT -55.740 134.890 -55.240 135.120 ;
        RECT -54.745 134.630 -54.505 135.350 ;
        RECT -52.700 134.885 -52.200 135.115 ;
        RECT -57.815 134.400 -57.315 134.630 ;
        RECT -55.740 134.400 -54.505 134.630 ;
        RECT -55.515 134.390 -54.505 134.400 ;
        RECT -51.850 134.095 -51.565 137.955 ;
        RECT -50.875 137.940 -50.375 138.170 ;
        RECT -44.035 137.940 -43.535 138.170 ;
        RECT -42.895 137.955 -42.525 138.800 ;
        RECT -41.960 138.430 -41.460 138.660 ;
        RECT -51.300 136.845 -50.300 137.075 ;
        RECT -44.110 136.845 -43.110 137.075 ;
        RECT -51.300 135.865 -50.300 136.095 ;
        RECT -44.110 135.865 -43.110 136.095 ;
        RECT -51.300 134.885 -50.300 135.115 ;
        RECT -44.110 134.885 -43.110 135.115 ;
        RECT -42.845 134.095 -42.560 137.955 ;
        RECT -41.960 137.940 -41.460 138.170 ;
        RECT -39.905 137.590 -39.665 141.840 ;
        RECT -38.070 141.905 -36.610 142.190 ;
        RECT -38.920 140.885 -38.420 141.115 ;
        RECT -38.920 139.905 -38.420 140.135 ;
        RECT -38.920 138.925 -38.420 139.155 ;
        RECT -39.170 137.830 -38.670 138.060 ;
        RECT -38.070 138.045 -37.785 141.905 ;
        RECT -37.520 140.885 -36.520 141.115 ;
        RECT -37.520 139.905 -36.520 140.135 ;
        RECT -37.520 138.925 -36.520 139.155 ;
        RECT -39.905 137.570 -39.075 137.590 ;
        RECT -39.905 137.340 -38.670 137.570 ;
        RECT -39.905 137.285 -39.075 137.340 ;
        RECT -42.210 136.845 -41.710 137.075 ;
        RECT -39.905 136.635 -39.665 137.285 ;
        RECT -38.105 137.200 -37.735 138.045 ;
        RECT -37.095 137.830 -36.595 138.060 ;
        RECT -37.095 137.340 -36.595 137.570 ;
        RECT -39.170 136.850 -38.670 137.080 ;
        RECT -37.095 136.850 -36.595 137.080 ;
        RECT -39.905 136.590 -39.065 136.635 ;
        RECT -39.905 136.360 -38.670 136.590 ;
        RECT -37.095 136.360 -36.595 136.590 ;
        RECT -39.905 136.330 -39.065 136.360 ;
        RECT -42.210 135.865 -41.710 136.095 ;
        RECT -39.905 135.655 -39.665 136.330 ;
        RECT -39.170 135.870 -38.670 136.100 ;
        RECT -37.095 135.870 -36.595 136.100 ;
        RECT -39.905 135.610 -39.075 135.655 ;
        RECT -39.905 135.380 -38.670 135.610 ;
        RECT -37.095 135.380 -36.595 135.610 ;
        RECT -39.905 135.350 -39.075 135.380 ;
        RECT -42.210 134.885 -41.710 135.115 ;
        RECT -39.905 134.630 -39.665 135.350 ;
        RECT -39.170 134.890 -38.670 135.120 ;
        RECT -37.095 134.890 -36.595 135.120 ;
        RECT -39.905 134.400 -38.670 134.630 ;
        RECT -37.095 134.400 -36.595 134.630 ;
        RECT -39.905 134.390 -38.895 134.400 ;
        RECT -54.705 133.805 -54.405 133.985 ;
        RECT -51.850 133.810 -50.390 134.095 ;
        RECT -44.020 133.810 -42.560 134.095 ;
        RECT -54.705 133.505 -52.070 133.805 ;
        RECT -54.705 133.325 -54.405 133.505 ;
        RECT -52.700 132.660 -52.200 132.890 ;
        RECT -51.300 132.660 -50.300 132.890 ;
        RECT -44.110 132.660 -43.110 132.890 ;
        RECT -42.210 132.660 -41.710 132.890 ;
        RECT -57.890 132.170 -56.890 132.400 ;
        RECT -55.990 132.170 -55.490 132.400 ;
        RECT -38.920 132.170 -38.420 132.400 ;
        RECT -37.520 132.170 -36.520 132.400 ;
        RECT -52.700 131.680 -52.200 131.910 ;
        RECT -51.300 131.680 -50.300 131.910 ;
        RECT -44.110 131.680 -43.110 131.910 ;
        RECT -42.210 131.680 -41.710 131.910 ;
        RECT -57.890 131.190 -56.890 131.420 ;
        RECT -55.990 131.190 -55.490 131.420 ;
        RECT -38.920 131.190 -38.420 131.420 ;
        RECT -37.520 131.190 -36.520 131.420 ;
        RECT -52.700 130.700 -52.200 130.930 ;
        RECT -51.300 130.700 -50.300 130.930 ;
        RECT -44.110 130.700 -43.110 130.930 ;
        RECT -42.210 130.700 -41.710 130.930 ;
        RECT -57.890 130.210 -56.890 130.440 ;
        RECT -55.990 130.210 -55.490 130.440 ;
        RECT -38.920 130.210 -38.420 130.440 ;
        RECT -37.520 130.210 -36.520 130.440 ;
        RECT -54.555 129.640 -53.870 129.940 ;
        RECT -40.540 129.640 -39.855 129.940 ;
        RECT -60.025 129.205 -59.760 129.265 ;
        RECT -60.025 128.585 -59.795 129.205 ;
        RECT -54.425 128.785 -54.105 129.640 ;
        RECT -54.580 127.910 -53.010 128.785 ;
        RECT -40.305 127.950 -39.985 129.640 ;
        RECT -34.650 129.265 -34.440 175.710 ;
        RECT -34.240 141.665 -34.030 176.230 ;
        RECT -34.250 140.985 -34.020 141.665 ;
        RECT -33.435 139.650 -33.180 210.415 ;
        RECT -32.685 152.505 -32.430 211.195 ;
        RECT -32.005 164.865 -31.865 212.105 ;
        RECT -31.370 177.240 -31.180 212.815 ;
        RECT -30.655 207.765 -29.930 213.630 ;
        RECT -30.655 193.765 -30.515 207.765 ;
        RECT -27.140 207.705 -27.000 214.410 ;
        RECT -27.140 206.705 -25.240 207.705 ;
        RECT -27.140 203.895 -27.000 206.705 ;
        RECT -27.210 203.200 -26.940 203.895 ;
        RECT -29.390 202.755 -28.390 202.985 ;
        RECT -27.510 202.265 -27.280 202.945 ;
        RECT -29.390 201.210 -28.390 201.440 ;
        RECT -28.230 200.735 -28.000 201.390 ;
        RECT -29.390 200.150 -28.390 200.380 ;
        RECT -29.390 199.660 -28.390 199.890 ;
        RECT -29.390 198.680 -28.390 198.910 ;
        RECT -29.390 198.190 -28.390 198.420 ;
        RECT -29.390 196.870 -28.390 197.100 ;
        RECT -28.200 196.105 -28.060 200.735 ;
        RECT -27.465 198.775 -27.325 202.265 ;
        RECT -27.140 200.820 -27.000 203.200 ;
        RECT -26.360 202.755 -25.360 202.985 ;
        RECT -26.360 201.210 -25.360 201.440 ;
        RECT -27.180 200.125 -26.910 200.820 ;
        RECT -26.360 199.660 -25.360 199.890 ;
        RECT -27.550 198.080 -27.280 198.775 ;
        RECT -26.360 198.680 -25.360 198.910 ;
        RECT -26.360 196.870 -25.360 197.100 ;
        RECT -26.360 196.380 -25.360 196.610 ;
        RECT -28.200 195.965 -27.195 196.105 ;
        RECT -27.335 195.030 -27.195 195.965 ;
        RECT -26.360 195.890 -25.360 196.120 ;
        RECT -26.360 195.290 -25.360 195.520 ;
        RECT -29.390 194.800 -28.390 195.030 ;
        RECT -27.400 194.335 -27.130 195.030 ;
        RECT -26.360 194.800 -25.360 195.030 ;
        RECT -26.360 194.310 -25.360 194.540 ;
        RECT -30.655 193.625 -27.000 193.765 ;
        RECT -30.955 192.945 -30.725 193.140 ;
        RECT -29.245 192.945 -28.565 192.950 ;
        RECT -30.955 192.725 -28.565 192.945 ;
        RECT -30.955 192.460 -30.725 192.725 ;
        RECT -29.245 192.720 -28.565 192.725 ;
        RECT -27.140 188.895 -27.000 193.625 ;
        RECT -27.210 188.200 -26.940 188.895 ;
        RECT -29.390 187.755 -28.390 187.985 ;
        RECT -27.510 187.265 -27.280 187.945 ;
        RECT -29.390 186.210 -28.390 186.440 ;
        RECT -28.230 185.735 -28.000 186.390 ;
        RECT -29.390 185.150 -28.390 185.380 ;
        RECT -29.390 184.660 -28.390 184.890 ;
        RECT -29.390 183.680 -28.390 183.910 ;
        RECT -29.390 183.190 -28.390 183.420 ;
        RECT -29.390 181.870 -28.390 182.100 ;
        RECT -28.200 181.105 -28.060 185.735 ;
        RECT -27.465 183.775 -27.325 187.265 ;
        RECT -27.140 185.820 -27.000 188.200 ;
        RECT -26.360 187.755 -25.360 187.985 ;
        RECT -26.360 186.210 -25.360 186.440 ;
        RECT -27.180 185.125 -26.910 185.820 ;
        RECT -26.360 184.660 -25.360 184.890 ;
        RECT -27.550 183.080 -27.280 183.775 ;
        RECT -26.360 183.680 -25.360 183.910 ;
        RECT -26.360 181.870 -25.360 182.100 ;
        RECT -26.360 181.380 -25.360 181.610 ;
        RECT -28.200 180.965 -27.195 181.105 ;
        RECT -27.335 180.030 -27.195 180.965 ;
        RECT -26.360 180.890 -25.360 181.120 ;
        RECT -26.360 180.290 -25.360 180.520 ;
        RECT -29.390 179.800 -28.390 180.030 ;
        RECT -27.400 179.335 -27.130 180.030 ;
        RECT -26.360 179.800 -25.360 180.030 ;
        RECT -26.360 179.310 -25.360 179.540 ;
        RECT -31.035 178.420 -30.805 178.615 ;
        RECT -29.245 178.420 -28.565 178.425 ;
        RECT -31.035 178.200 -28.565 178.420 ;
        RECT -31.035 177.935 -30.805 178.200 ;
        RECT -29.245 178.195 -28.565 178.200 ;
        RECT -31.370 177.100 -27.000 177.240 ;
        RECT -27.140 176.395 -27.000 177.100 ;
        RECT -27.210 175.700 -26.940 176.395 ;
        RECT -29.390 175.255 -28.390 175.485 ;
        RECT -27.510 174.765 -27.280 175.445 ;
        RECT -29.390 173.710 -28.390 173.940 ;
        RECT -28.230 173.235 -28.000 173.890 ;
        RECT -29.390 172.650 -28.390 172.880 ;
        RECT -29.390 172.160 -28.390 172.390 ;
        RECT -29.390 171.180 -28.390 171.410 ;
        RECT -29.390 170.690 -28.390 170.920 ;
        RECT -29.390 169.370 -28.390 169.600 ;
        RECT -28.200 168.605 -28.060 173.235 ;
        RECT -27.465 171.275 -27.325 174.765 ;
        RECT -27.140 173.320 -27.000 175.700 ;
        RECT -26.360 175.255 -25.360 175.485 ;
        RECT -26.360 173.710 -25.360 173.940 ;
        RECT -27.180 172.625 -26.910 173.320 ;
        RECT -26.360 172.160 -25.360 172.390 ;
        RECT -27.550 170.580 -27.280 171.275 ;
        RECT -26.360 171.180 -25.360 171.410 ;
        RECT -26.360 169.370 -25.360 169.600 ;
        RECT -26.360 168.880 -25.360 169.110 ;
        RECT -28.200 168.465 -27.195 168.605 ;
        RECT -30.720 167.020 -30.490 167.700 ;
        RECT -27.335 167.530 -27.195 168.465 ;
        RECT -26.360 168.390 -25.360 168.620 ;
        RECT -26.360 167.790 -25.360 168.020 ;
        RECT -29.390 167.300 -28.390 167.530 ;
        RECT -30.715 166.335 -30.495 167.020 ;
        RECT -27.400 166.835 -27.130 167.530 ;
        RECT -26.360 167.300 -25.360 167.530 ;
        RECT -26.360 166.810 -25.360 167.040 ;
        RECT -29.245 166.335 -28.565 166.340 ;
        RECT -30.715 166.115 -28.565 166.335 ;
        RECT -29.245 166.110 -28.565 166.115 ;
        RECT -32.005 164.725 -27.000 164.865 ;
        RECT -27.140 163.895 -27.000 164.725 ;
        RECT -27.210 163.200 -26.940 163.895 ;
        RECT -29.390 162.755 -28.390 162.985 ;
        RECT -27.510 162.265 -27.280 162.945 ;
        RECT -29.390 161.210 -28.390 161.440 ;
        RECT -28.230 160.735 -28.000 161.390 ;
        RECT -29.390 160.150 -28.390 160.380 ;
        RECT -29.390 159.660 -28.390 159.890 ;
        RECT -29.390 158.680 -28.390 158.910 ;
        RECT -29.390 158.190 -28.390 158.420 ;
        RECT -29.390 156.870 -28.390 157.100 ;
        RECT -28.200 156.105 -28.060 160.735 ;
        RECT -27.465 158.775 -27.325 162.265 ;
        RECT -27.140 160.820 -27.000 163.200 ;
        RECT -26.360 162.755 -25.360 162.985 ;
        RECT -26.360 161.210 -25.360 161.440 ;
        RECT -27.180 160.125 -26.910 160.820 ;
        RECT -26.360 159.660 -25.360 159.890 ;
        RECT -27.550 158.080 -27.280 158.775 ;
        RECT -26.360 158.680 -25.360 158.910 ;
        RECT -26.360 156.870 -25.360 157.100 ;
        RECT -26.360 156.380 -25.360 156.610 ;
        RECT -28.200 155.965 -27.195 156.105 ;
        RECT -30.655 154.535 -30.425 155.215 ;
        RECT -27.335 155.030 -27.195 155.965 ;
        RECT -26.360 155.890 -25.360 156.120 ;
        RECT -26.360 155.290 -25.360 155.520 ;
        RECT -29.390 154.800 -28.390 155.030 ;
        RECT -30.650 153.935 -30.430 154.535 ;
        RECT -27.400 154.335 -27.130 155.030 ;
        RECT -26.360 154.800 -25.360 155.030 ;
        RECT -26.360 154.310 -25.360 154.540 ;
        RECT -29.245 153.935 -28.565 153.940 ;
        RECT -30.650 153.715 -28.565 153.935 ;
        RECT -30.650 153.710 -30.430 153.715 ;
        RECT -29.245 153.710 -28.565 153.715 ;
        RECT -32.685 152.365 -27.000 152.505 ;
        RECT -27.140 151.395 -27.000 152.365 ;
        RECT -27.210 150.700 -26.940 151.395 ;
        RECT -29.390 150.255 -28.390 150.485 ;
        RECT -27.510 149.765 -27.280 150.445 ;
        RECT -29.390 148.710 -28.390 148.940 ;
        RECT -28.230 148.235 -28.000 148.890 ;
        RECT -29.390 147.650 -28.390 147.880 ;
        RECT -29.390 147.160 -28.390 147.390 ;
        RECT -29.390 146.180 -28.390 146.410 ;
        RECT -29.390 145.690 -28.390 145.920 ;
        RECT -29.390 144.370 -28.390 144.600 ;
        RECT -28.200 143.605 -28.060 148.235 ;
        RECT -27.465 146.275 -27.325 149.765 ;
        RECT -27.140 148.320 -27.000 150.700 ;
        RECT -26.360 150.255 -25.360 150.485 ;
        RECT -26.360 148.710 -25.360 148.940 ;
        RECT -27.180 147.625 -26.910 148.320 ;
        RECT -26.360 147.160 -25.360 147.390 ;
        RECT -27.550 145.580 -27.280 146.275 ;
        RECT -26.360 146.180 -25.360 146.410 ;
        RECT -26.360 144.370 -25.360 144.600 ;
        RECT -26.360 143.880 -25.360 144.110 ;
        RECT -28.200 143.465 -27.195 143.605 ;
        RECT -27.335 142.530 -27.195 143.465 ;
        RECT -26.360 143.390 -25.360 143.620 ;
        RECT -26.360 142.790 -25.360 143.020 ;
        RECT -29.390 142.300 -28.390 142.530 ;
        RECT -27.400 141.835 -27.130 142.530 ;
        RECT -26.360 142.300 -25.360 142.530 ;
        RECT -26.360 141.810 -25.360 142.040 ;
        RECT -32.755 141.195 -32.075 141.200 ;
        RECT -29.225 141.195 -28.545 141.200 ;
        RECT -32.755 140.975 -28.545 141.195 ;
        RECT -32.755 140.970 -32.075 140.975 ;
        RECT -29.225 140.970 -28.545 140.975 ;
        RECT -33.435 139.510 -27.000 139.650 ;
        RECT -31.700 139.150 -27.685 139.290 ;
        RECT -31.700 139.060 -31.020 139.150 ;
        RECT -29.390 137.755 -28.390 137.985 ;
        RECT -27.825 137.330 -27.685 139.150 ;
        RECT -27.140 138.895 -27.000 139.510 ;
        RECT -27.210 138.200 -26.940 138.895 ;
        RECT -27.950 136.635 -27.680 137.330 ;
        RECT -27.510 137.265 -27.280 137.945 ;
        RECT -29.390 136.210 -28.390 136.440 ;
        RECT -28.230 135.735 -28.000 136.390 ;
        RECT -29.390 135.150 -28.390 135.380 ;
        RECT -29.390 134.660 -28.390 134.890 ;
        RECT -33.005 133.945 -32.005 134.175 ;
        RECT -31.105 133.945 -30.605 134.175 ;
        RECT -29.390 133.680 -28.390 133.910 ;
        RECT -33.005 132.965 -32.005 133.195 ;
        RECT -31.105 132.965 -30.605 133.195 ;
        RECT -29.390 133.190 -28.390 133.420 ;
        RECT -33.005 131.985 -32.005 132.215 ;
        RECT -31.105 131.985 -30.605 132.215 ;
        RECT -29.390 131.870 -28.390 132.100 ;
        RECT -28.200 131.105 -28.060 135.735 ;
        RECT -27.835 131.940 -27.695 136.635 ;
        RECT -27.465 133.775 -27.325 137.265 ;
        RECT -27.140 135.820 -27.000 138.200 ;
        RECT -26.360 137.755 -25.360 137.985 ;
        RECT -26.360 136.210 -25.360 136.440 ;
        RECT -27.180 135.125 -26.910 135.820 ;
        RECT -26.360 134.660 -25.360 134.890 ;
        RECT -27.550 133.080 -27.280 133.775 ;
        RECT -26.360 133.680 -25.360 133.910 ;
        RECT -27.920 131.245 -27.650 131.940 ;
        RECT -26.360 131.870 -25.360 132.100 ;
        RECT -26.360 131.380 -25.360 131.610 ;
        RECT -28.200 130.965 -27.195 131.105 ;
        RECT -27.335 130.030 -27.195 130.965 ;
        RECT -26.360 130.890 -25.360 131.120 ;
        RECT -26.360 130.290 -25.360 130.520 ;
        RECT -29.390 129.800 -28.390 130.030 ;
        RECT -27.400 129.335 -27.130 130.030 ;
        RECT -26.360 129.800 -25.360 130.030 ;
        RECT -26.360 129.310 -25.360 129.540 ;
        RECT -34.660 128.585 -34.430 129.265 ;
        RECT -40.300 127.865 -39.985 127.950 ;
        RECT -83.320 127.235 -82.640 127.255 ;
        RECT -70.865 127.235 -69.990 127.335 ;
        RECT -83.320 126.575 -27.630 127.235 ;
        RECT -70.865 126.520 -69.990 126.575 ;
        RECT -52.050 125.390 -49.050 125.620 ;
        RECT -27.380 125.255 -24.380 125.485 ;
        RECT -55.110 124.900 -53.610 125.130 ;
        RECT -30.440 124.765 -28.940 124.995 ;
        RECT -52.050 124.335 -49.050 124.565 ;
        RECT -27.380 124.200 -24.380 124.430 ;
        RECT -52.050 123.845 -49.050 124.075 ;
        RECT -27.380 123.710 -24.380 123.940 ;
        RECT -52.050 123.355 -49.050 123.585 ;
        RECT -27.380 123.220 -24.380 123.450 ;
        RECT -55.110 122.710 -53.610 122.940 ;
        RECT -30.440 122.575 -28.940 122.805 ;
        RECT -52.050 122.295 -49.050 122.525 ;
        RECT -27.380 122.160 -24.380 122.390 ;
        RECT -69.555 121.780 -68.700 121.835 ;
        RECT -69.555 120.900 -36.125 121.780 ;
        RECT -69.555 120.835 -68.700 120.900 ;
        RECT -56.555 119.425 -55.555 119.655 ;
        RECT -54.655 119.425 -54.155 119.655 ;
        RECT -31.920 119.425 -30.920 119.655 ;
        RECT -30.020 119.425 -29.520 119.655 ;
        RECT -56.555 118.445 -55.555 118.675 ;
        RECT -54.655 118.445 -54.155 118.675 ;
        RECT -31.920 118.445 -30.920 118.675 ;
        RECT -30.020 118.445 -29.520 118.675 ;
        RECT -56.555 117.465 -55.555 117.695 ;
        RECT -54.655 117.465 -54.155 117.695 ;
        RECT -31.920 117.465 -30.920 117.695 ;
        RECT -30.020 117.465 -29.520 117.695 ;
        RECT -53.360 117.025 -53.060 117.230 ;
        RECT -28.725 117.025 -28.425 117.230 ;
        RECT -55.160 116.735 -53.060 117.025 ;
        RECT -55.160 116.725 -54.500 116.735 ;
        RECT -53.360 116.570 -53.060 116.735 ;
        RECT -30.525 116.735 -28.425 117.025 ;
        RECT -30.525 116.725 -29.865 116.735 ;
        RECT -28.725 116.570 -28.425 116.735 ;
        RECT -57.180 116.035 -55.005 116.320 ;
        RECT -52.355 116.170 -50.455 116.210 ;
        RECT -57.180 98.215 -56.895 116.035 ;
        RECT -56.555 115.015 -55.555 115.245 ;
        RECT -56.555 114.035 -55.555 114.265 ;
        RECT -56.555 113.055 -55.555 113.285 ;
        RECT -56.480 111.960 -55.980 112.190 ;
        RECT -55.290 112.175 -55.005 116.035 ;
        RECT -52.360 115.980 -50.455 116.170 ;
        RECT -54.655 115.015 -54.155 115.245 ;
        RECT -54.655 114.035 -54.155 114.265 ;
        RECT -54.655 113.055 -54.155 113.285 ;
        RECT -52.360 112.345 -52.130 115.980 ;
        RECT -51.615 115.500 -51.115 115.730 ;
        RECT -50.755 115.440 -50.455 115.980 ;
        RECT -32.545 116.035 -30.370 116.320 ;
        RECT -27.720 116.170 -25.820 116.210 ;
        RECT -49.540 115.500 -49.040 115.730 ;
        RECT -51.615 115.010 -51.115 115.240 ;
        RECT -49.540 115.010 -49.040 115.240 ;
        RECT -51.615 114.520 -51.115 114.750 ;
        RECT -49.540 114.520 -49.040 114.750 ;
        RECT -51.615 114.030 -51.115 114.260 ;
        RECT -49.540 114.030 -49.040 114.260 ;
        RECT -51.615 113.540 -51.115 113.770 ;
        RECT -49.540 113.540 -49.040 113.770 ;
        RECT -51.615 113.050 -51.115 113.280 ;
        RECT -49.540 113.050 -49.040 113.280 ;
        RECT -51.615 112.560 -51.115 112.790 ;
        RECT -56.480 111.470 -55.980 111.700 ;
        RECT -55.340 111.330 -54.970 112.175 ;
        RECT -54.405 111.960 -53.905 112.190 ;
        RECT -53.420 112.115 -52.130 112.345 ;
        RECT -54.405 111.685 -53.905 111.700 ;
        RECT -53.420 111.685 -53.190 112.115 ;
        RECT -51.615 112.070 -51.115 112.300 ;
        RECT -50.550 112.085 -50.180 112.930 ;
        RECT -49.540 112.560 -49.040 112.790 ;
        RECT -54.405 111.475 -53.190 111.685 ;
        RECT -54.405 111.470 -53.905 111.475 ;
        RECT -56.480 110.980 -55.980 111.210 ;
        RECT -54.405 110.980 -53.905 111.210 ;
        RECT -56.480 110.490 -55.980 110.720 ;
        RECT -54.405 110.705 -53.905 110.720 ;
        RECT -53.420 110.705 -53.190 111.475 ;
        RECT -51.365 110.975 -50.865 111.205 ;
        RECT -54.405 110.495 -53.190 110.705 ;
        RECT -54.405 110.490 -53.905 110.495 ;
        RECT -56.480 110.000 -55.980 110.230 ;
        RECT -54.405 110.000 -53.905 110.230 ;
        RECT -56.480 109.510 -55.980 109.740 ;
        RECT -54.405 109.730 -53.905 109.740 ;
        RECT -53.420 109.730 -53.190 110.495 ;
        RECT -51.365 109.995 -50.865 110.225 ;
        RECT -54.405 109.520 -53.190 109.730 ;
        RECT -54.405 109.510 -53.905 109.520 ;
        RECT -56.480 109.020 -55.980 109.250 ;
        RECT -54.405 109.020 -53.905 109.250 ;
        RECT -53.420 108.775 -53.190 109.520 ;
        RECT -51.365 109.015 -50.865 109.245 ;
        RECT -56.480 108.530 -55.980 108.760 ;
        RECT -54.405 108.545 -53.190 108.775 ;
        RECT -54.405 108.530 -53.905 108.545 ;
        RECT -50.515 108.225 -50.230 112.085 ;
        RECT -49.540 112.070 -49.040 112.300 ;
        RECT -49.965 110.975 -48.965 111.205 ;
        RECT -49.965 109.995 -48.965 110.225 ;
        RECT -49.965 109.015 -48.965 109.245 ;
        RECT -37.215 108.295 -36.855 108.465 ;
        RECT -52.930 107.995 -52.630 108.210 ;
        RECT -52.930 107.695 -50.810 107.995 ;
        RECT -50.515 107.940 -49.055 108.225 ;
        RECT -37.215 107.970 -36.115 108.295 ;
        RECT -37.215 107.940 -36.855 107.970 ;
        RECT -52.930 107.550 -52.630 107.695 ;
        RECT -51.365 106.790 -50.865 107.020 ;
        RECT -49.965 106.790 -48.965 107.020 ;
        RECT -44.070 106.685 -43.840 107.680 ;
        RECT -40.510 106.785 -37.510 107.015 ;
        RECT -56.555 106.300 -55.555 106.530 ;
        RECT -54.655 106.300 -54.155 106.530 ;
        RECT -44.070 106.455 -43.060 106.685 ;
        RECT -44.070 106.195 -43.840 106.455 ;
        RECT -51.365 105.810 -50.865 106.040 ;
        RECT -49.965 105.810 -48.965 106.040 ;
        RECT -44.715 105.965 -43.830 106.195 ;
        RECT -44.070 105.705 -43.830 105.965 ;
        RECT -40.510 105.725 -37.510 105.955 ;
        RECT -56.555 105.320 -55.555 105.550 ;
        RECT -54.655 105.320 -54.155 105.550 ;
        RECT -44.070 105.475 -43.060 105.705 ;
        RECT -44.070 105.215 -43.830 105.475 ;
        RECT -40.510 105.235 -37.510 105.465 ;
        RECT -51.365 104.830 -50.865 105.060 ;
        RECT -49.965 104.830 -48.965 105.060 ;
        RECT -44.715 104.985 -43.830 105.215 ;
        RECT -44.070 104.725 -43.840 104.985 ;
        RECT -40.510 104.745 -37.510 104.975 ;
        RECT -56.555 104.340 -55.555 104.570 ;
        RECT -54.655 104.340 -54.155 104.570 ;
        RECT -44.070 104.495 -43.060 104.725 ;
        RECT -50.640 103.945 -50.340 104.360 ;
        RECT -54.605 103.940 -50.310 103.945 ;
        RECT -55.040 103.645 -50.310 103.940 ;
        RECT -40.510 103.690 -37.510 103.920 ;
        RECT -55.040 103.640 -54.380 103.645 ;
        RECT -52.925 103.365 -52.625 103.505 ;
        RECT -55.165 103.065 -52.625 103.365 ;
        RECT -36.440 103.195 -36.115 107.970 ;
        RECT -35.950 106.370 -34.450 106.600 ;
        RECT -35.950 104.180 -34.450 104.410 ;
        RECT -52.925 102.820 -52.625 103.065 ;
        RECT -47.665 102.920 -45.750 103.150 ;
        RECT -56.465 102.535 -55.005 102.820 ;
        RECT -50.745 102.675 -50.445 102.680 ;
        RECT -56.555 101.515 -55.555 101.745 ;
        RECT -56.555 100.535 -55.555 100.765 ;
        RECT -56.555 99.555 -55.555 99.785 ;
        RECT -56.480 98.460 -55.980 98.690 ;
        RECT -55.290 98.675 -55.005 102.535 ;
        RECT -53.410 102.470 -50.440 102.675 ;
        RECT -54.655 101.515 -54.155 101.745 ;
        RECT -54.655 100.535 -54.155 100.765 ;
        RECT -54.655 99.555 -54.155 99.785 ;
        RECT -57.180 98.200 -56.290 98.215 ;
        RECT -57.180 97.970 -55.980 98.200 ;
        RECT -57.180 97.960 -56.290 97.970 ;
        RECT -57.180 97.245 -56.895 97.960 ;
        RECT -55.340 97.830 -54.970 98.675 ;
        RECT -54.405 98.460 -53.905 98.690 ;
        RECT -53.410 98.220 -53.170 102.470 ;
        RECT -51.615 102.000 -51.115 102.230 ;
        RECT -50.745 101.995 -50.445 102.470 ;
        RECT -49.540 102.000 -49.040 102.230 ;
        RECT -47.665 102.170 -47.430 102.920 ;
        RECT -47.250 102.430 -43.065 102.660 ;
        RECT -47.665 101.940 -45.750 102.170 ;
        RECT -51.615 101.510 -51.115 101.740 ;
        RECT -49.540 101.510 -49.040 101.740 ;
        RECT -51.615 101.020 -51.115 101.250 ;
        RECT -49.540 101.020 -49.040 101.250 ;
        RECT -47.665 101.190 -47.430 101.940 ;
        RECT -39.290 101.690 -39.060 102.685 ;
        RECT -44.565 101.450 -43.065 101.680 ;
        RECT -40.070 101.460 -39.060 101.690 ;
        RECT -47.665 100.960 -45.750 101.190 ;
        RECT -47.665 100.955 -47.245 100.960 ;
        RECT -45.085 100.880 -44.795 101.275 ;
        RECT -39.290 101.200 -39.060 101.460 ;
        RECT -51.615 100.530 -51.115 100.760 ;
        RECT -49.540 100.530 -49.040 100.760 ;
        RECT -45.630 100.610 -44.795 100.880 ;
        RECT -39.300 100.970 -38.415 101.200 ;
        RECT -39.300 100.710 -39.060 100.970 ;
        RECT -51.615 100.040 -51.115 100.270 ;
        RECT -49.540 100.040 -49.040 100.270 ;
        RECT -51.615 99.550 -51.115 99.780 ;
        RECT -49.540 99.550 -49.040 99.780 ;
        RECT -45.630 99.510 -45.360 100.610 ;
        RECT -45.085 100.480 -44.795 100.610 ;
        RECT -40.070 100.480 -39.060 100.710 ;
        RECT -39.300 100.220 -39.060 100.480 ;
        RECT -39.300 99.990 -38.415 100.220 ;
        RECT -51.615 99.060 -51.115 99.290 ;
        RECT -51.615 98.570 -51.115 98.800 ;
        RECT -50.550 98.585 -50.180 99.430 ;
        RECT -49.540 99.060 -49.040 99.290 ;
        RECT -47.350 99.240 -45.360 99.510 ;
        RECT -54.000 98.200 -53.170 98.220 ;
        RECT -54.405 97.970 -53.170 98.200 ;
        RECT -54.000 97.915 -53.170 97.970 ;
        RECT -56.480 97.480 -55.980 97.710 ;
        RECT -54.405 97.480 -53.905 97.710 ;
        RECT -53.410 97.265 -53.170 97.915 ;
        RECT -51.365 97.475 -50.865 97.705 ;
        RECT -57.180 97.220 -56.290 97.245 ;
        RECT -54.010 97.220 -53.170 97.265 ;
        RECT -57.180 96.990 -55.980 97.220 ;
        RECT -54.405 96.990 -53.170 97.220 ;
        RECT -57.180 96.245 -56.895 96.990 ;
        RECT -54.010 96.960 -53.170 96.990 ;
        RECT -56.480 96.500 -55.980 96.730 ;
        RECT -54.405 96.500 -53.905 96.730 ;
        RECT -53.410 96.285 -53.170 96.960 ;
        RECT -51.365 96.495 -50.865 96.725 ;
        RECT -57.180 96.240 -56.195 96.245 ;
        RECT -54.000 96.240 -53.170 96.285 ;
        RECT -57.180 96.010 -55.980 96.240 ;
        RECT -54.405 96.010 -53.170 96.240 ;
        RECT -57.180 95.990 -56.195 96.010 ;
        RECT -57.180 95.285 -56.895 95.990 ;
        RECT -54.000 95.980 -53.170 96.010 ;
        RECT -56.480 95.520 -55.980 95.750 ;
        RECT -54.405 95.520 -53.905 95.750 ;
        RECT -57.180 95.260 -56.320 95.285 ;
        RECT -53.410 95.260 -53.170 95.980 ;
        RECT -51.365 95.515 -50.865 95.745 ;
        RECT -57.180 95.035 -55.980 95.260 ;
        RECT -56.480 95.030 -55.980 95.035 ;
        RECT -54.405 95.030 -53.170 95.260 ;
        RECT -54.180 95.020 -53.170 95.030 ;
        RECT -50.515 94.725 -50.230 98.585 ;
        RECT -49.540 98.570 -49.040 98.800 ;
        RECT -49.965 97.475 -48.965 97.705 ;
        RECT -49.965 96.495 -48.965 96.725 ;
        RECT -49.965 95.515 -48.965 95.745 ;
        RECT -53.370 94.435 -53.070 94.615 ;
        RECT -50.515 94.440 -49.055 94.725 ;
        RECT -53.370 94.135 -50.735 94.435 ;
        RECT -53.370 93.955 -53.070 94.135 ;
        RECT -51.365 93.290 -50.865 93.520 ;
        RECT -49.965 93.290 -48.965 93.520 ;
        RECT -56.555 92.800 -55.555 93.030 ;
        RECT -54.655 92.800 -54.155 93.030 ;
        RECT -51.365 92.310 -50.865 92.540 ;
        RECT -49.965 92.310 -48.965 92.540 ;
        RECT -56.555 91.820 -55.555 92.050 ;
        RECT -54.655 91.820 -54.155 92.050 ;
        RECT -51.365 91.330 -50.865 91.560 ;
        RECT -49.965 91.330 -48.965 91.560 ;
        RECT -56.555 90.840 -55.555 91.070 ;
        RECT -54.655 90.840 -54.155 91.070 ;
        RECT -53.220 90.270 -52.535 90.570 ;
        RECT -53.090 88.940 -52.770 90.270 ;
        RECT -47.350 88.940 -47.080 99.240 ;
        RECT -45.220 98.775 -44.990 99.770 ;
        RECT -39.290 99.730 -39.060 99.990 ;
        RECT -40.070 99.500 -39.060 99.730 ;
        RECT -45.220 98.545 -43.710 98.775 ;
        RECT -45.220 98.285 -44.990 98.545 ;
        RECT -46.360 98.055 -44.980 98.285 ;
        RECT -32.545 98.215 -32.260 116.035 ;
        RECT -31.920 115.015 -30.920 115.245 ;
        RECT -31.920 114.035 -30.920 114.265 ;
        RECT -31.920 113.055 -30.920 113.285 ;
        RECT -31.845 111.960 -31.345 112.190 ;
        RECT -30.655 112.175 -30.370 116.035 ;
        RECT -27.725 115.980 -25.820 116.170 ;
        RECT -30.020 115.015 -29.520 115.245 ;
        RECT -30.020 114.035 -29.520 114.265 ;
        RECT -30.020 113.055 -29.520 113.285 ;
        RECT -27.725 112.345 -27.495 115.980 ;
        RECT -26.980 115.500 -26.480 115.730 ;
        RECT -26.120 115.440 -25.820 115.980 ;
        RECT -24.905 115.500 -24.405 115.730 ;
        RECT -26.980 115.010 -26.480 115.240 ;
        RECT -24.905 115.010 -24.405 115.240 ;
        RECT -26.980 114.520 -26.480 114.750 ;
        RECT -24.905 114.520 -24.405 114.750 ;
        RECT -26.980 114.030 -26.480 114.260 ;
        RECT -24.905 114.030 -24.405 114.260 ;
        RECT -26.980 113.540 -26.480 113.770 ;
        RECT -24.905 113.540 -24.405 113.770 ;
        RECT -26.980 113.050 -26.480 113.280 ;
        RECT -24.905 113.050 -24.405 113.280 ;
        RECT -26.980 112.560 -26.480 112.790 ;
        RECT -31.845 111.470 -31.345 111.700 ;
        RECT -30.705 111.330 -30.335 112.175 ;
        RECT -29.770 111.960 -29.270 112.190 ;
        RECT -28.785 112.115 -27.495 112.345 ;
        RECT -29.770 111.685 -29.270 111.700 ;
        RECT -28.785 111.685 -28.555 112.115 ;
        RECT -26.980 112.070 -26.480 112.300 ;
        RECT -25.915 112.085 -25.545 112.930 ;
        RECT -24.905 112.560 -24.405 112.790 ;
        RECT -29.770 111.475 -28.555 111.685 ;
        RECT -29.770 111.470 -29.270 111.475 ;
        RECT -31.845 110.980 -31.345 111.210 ;
        RECT -29.770 110.980 -29.270 111.210 ;
        RECT -31.845 110.490 -31.345 110.720 ;
        RECT -29.770 110.705 -29.270 110.720 ;
        RECT -28.785 110.705 -28.555 111.475 ;
        RECT -26.730 110.975 -26.230 111.205 ;
        RECT -29.770 110.495 -28.555 110.705 ;
        RECT -29.770 110.490 -29.270 110.495 ;
        RECT -31.845 110.000 -31.345 110.230 ;
        RECT -29.770 110.000 -29.270 110.230 ;
        RECT -31.845 109.510 -31.345 109.740 ;
        RECT -29.770 109.730 -29.270 109.740 ;
        RECT -28.785 109.730 -28.555 110.495 ;
        RECT -26.730 109.995 -26.230 110.225 ;
        RECT -29.770 109.520 -28.555 109.730 ;
        RECT -29.770 109.510 -29.270 109.520 ;
        RECT -31.845 109.020 -31.345 109.250 ;
        RECT -29.770 109.020 -29.270 109.250 ;
        RECT -28.785 108.775 -28.555 109.520 ;
        RECT -26.730 109.015 -26.230 109.245 ;
        RECT -31.845 108.530 -31.345 108.760 ;
        RECT -29.770 108.545 -28.555 108.775 ;
        RECT -29.770 108.530 -29.270 108.545 ;
        RECT -25.880 108.225 -25.595 112.085 ;
        RECT -24.905 112.070 -24.405 112.300 ;
        RECT -25.330 110.975 -24.330 111.205 ;
        RECT -25.330 109.995 -24.330 110.225 ;
        RECT -25.330 109.015 -24.330 109.245 ;
        RECT -28.295 107.995 -27.995 108.210 ;
        RECT -28.295 107.695 -26.175 107.995 ;
        RECT -25.880 107.940 -24.420 108.225 ;
        RECT -28.295 107.550 -27.995 107.695 ;
        RECT -26.730 106.790 -26.230 107.020 ;
        RECT -25.330 106.790 -24.330 107.020 ;
        RECT -31.920 106.300 -30.920 106.530 ;
        RECT -30.020 106.300 -29.520 106.530 ;
        RECT -26.730 105.810 -26.230 106.040 ;
        RECT -25.330 105.810 -24.330 106.040 ;
        RECT -31.920 105.320 -30.920 105.550 ;
        RECT -30.020 105.320 -29.520 105.550 ;
        RECT -26.730 104.830 -26.230 105.060 ;
        RECT -25.330 104.830 -24.330 105.060 ;
        RECT -31.920 104.340 -30.920 104.570 ;
        RECT -30.020 104.340 -29.520 104.570 ;
        RECT -26.005 103.945 -25.705 104.360 ;
        RECT -29.970 103.940 -25.675 103.945 ;
        RECT -30.405 103.645 -25.675 103.940 ;
        RECT -30.405 103.640 -29.745 103.645 ;
        RECT -28.290 103.365 -27.990 103.505 ;
        RECT -30.530 103.065 -27.990 103.365 ;
        RECT -28.290 102.820 -27.990 103.065 ;
        RECT -31.830 102.535 -30.370 102.820 ;
        RECT -26.110 102.675 -25.810 102.680 ;
        RECT -31.920 101.515 -30.920 101.745 ;
        RECT -31.920 100.535 -30.920 100.765 ;
        RECT -31.920 99.555 -30.920 99.785 ;
        RECT -31.845 98.460 -31.345 98.690 ;
        RECT -30.655 98.675 -30.370 102.535 ;
        RECT -28.775 102.470 -25.805 102.675 ;
        RECT -30.020 101.515 -29.520 101.745 ;
        RECT -30.020 100.535 -29.520 100.765 ;
        RECT -30.020 99.555 -29.520 99.785 ;
        RECT -32.545 98.200 -31.655 98.215 ;
        RECT -45.220 97.795 -44.980 98.055 ;
        RECT -37.380 97.925 -35.465 98.155 ;
        RECT -45.220 97.565 -43.710 97.795 ;
        RECT -45.220 97.305 -44.980 97.565 ;
        RECT -40.065 97.435 -35.880 97.665 ;
        RECT -46.360 97.075 -44.980 97.305 ;
        RECT -35.700 97.175 -35.465 97.925 ;
        RECT -45.220 96.815 -44.990 97.075 ;
        RECT -37.380 96.945 -35.465 97.175 ;
        RECT -45.220 96.585 -43.710 96.815 ;
        RECT -40.065 96.455 -38.565 96.685 ;
        RECT -35.700 96.195 -35.465 96.945 ;
        RECT -37.380 95.965 -35.465 96.195 ;
        RECT -35.885 95.960 -35.465 95.965 ;
        RECT -32.545 97.970 -31.345 98.200 ;
        RECT -32.545 97.960 -31.655 97.970 ;
        RECT -32.545 97.245 -32.260 97.960 ;
        RECT -30.705 97.830 -30.335 98.675 ;
        RECT -29.770 98.460 -29.270 98.690 ;
        RECT -28.775 98.220 -28.535 102.470 ;
        RECT -26.980 102.000 -26.480 102.230 ;
        RECT -26.110 101.995 -25.810 102.470 ;
        RECT -24.905 102.000 -24.405 102.230 ;
        RECT -26.980 101.510 -26.480 101.740 ;
        RECT -24.905 101.510 -24.405 101.740 ;
        RECT -26.980 101.020 -26.480 101.250 ;
        RECT -24.905 101.020 -24.405 101.250 ;
        RECT -26.980 100.530 -26.480 100.760 ;
        RECT -24.905 100.530 -24.405 100.760 ;
        RECT -26.980 100.040 -26.480 100.270 ;
        RECT -24.905 100.040 -24.405 100.270 ;
        RECT -26.980 99.550 -26.480 99.780 ;
        RECT -24.905 99.550 -24.405 99.780 ;
        RECT -26.980 99.060 -26.480 99.290 ;
        RECT -26.980 98.570 -26.480 98.800 ;
        RECT -25.915 98.585 -25.545 99.430 ;
        RECT -24.905 99.060 -24.405 99.290 ;
        RECT -29.365 98.200 -28.535 98.220 ;
        RECT -29.770 97.970 -28.535 98.200 ;
        RECT -29.365 97.915 -28.535 97.970 ;
        RECT -31.845 97.480 -31.345 97.710 ;
        RECT -29.770 97.480 -29.270 97.710 ;
        RECT -28.775 97.265 -28.535 97.915 ;
        RECT -26.730 97.475 -26.230 97.705 ;
        RECT -32.545 97.220 -31.655 97.245 ;
        RECT -29.375 97.220 -28.535 97.265 ;
        RECT -32.545 96.990 -31.345 97.220 ;
        RECT -29.770 96.990 -28.535 97.220 ;
        RECT -32.545 96.245 -32.260 96.990 ;
        RECT -29.375 96.960 -28.535 96.990 ;
        RECT -31.845 96.500 -31.345 96.730 ;
        RECT -29.770 96.500 -29.270 96.730 ;
        RECT -28.775 96.285 -28.535 96.960 ;
        RECT -26.730 96.495 -26.230 96.725 ;
        RECT -32.545 96.240 -31.560 96.245 ;
        RECT -29.365 96.240 -28.535 96.285 ;
        RECT -32.545 96.010 -31.345 96.240 ;
        RECT -29.770 96.010 -28.535 96.240 ;
        RECT -32.545 95.990 -31.560 96.010 ;
        RECT -32.545 95.285 -32.260 95.990 ;
        RECT -29.365 95.980 -28.535 96.010 ;
        RECT -31.845 95.520 -31.345 95.750 ;
        RECT -29.770 95.520 -29.270 95.750 ;
        RECT -32.545 95.260 -31.685 95.285 ;
        RECT -28.775 95.260 -28.535 95.980 ;
        RECT -26.730 95.515 -26.230 95.745 ;
        RECT -32.545 95.035 -31.345 95.260 ;
        RECT -31.845 95.030 -31.345 95.035 ;
        RECT -29.770 95.030 -28.535 95.260 ;
        RECT -29.545 95.020 -28.535 95.030 ;
        RECT -25.880 94.725 -25.595 98.585 ;
        RECT -24.905 98.570 -24.405 98.800 ;
        RECT -25.330 97.475 -24.330 97.705 ;
        RECT -25.330 96.495 -24.330 96.725 ;
        RECT -25.330 95.515 -24.330 95.745 ;
        RECT -28.735 94.435 -28.435 94.615 ;
        RECT -25.880 94.440 -24.420 94.725 ;
        RECT -38.595 93.270 -37.825 94.200 ;
        RECT -28.735 94.135 -26.100 94.435 ;
        RECT -28.735 93.955 -28.435 94.135 ;
        RECT -26.730 93.290 -26.230 93.520 ;
        RECT -25.330 93.290 -24.330 93.520 ;
        RECT -38.355 89.280 -38.035 93.270 ;
        RECT -31.920 92.800 -30.920 93.030 ;
        RECT -30.020 92.800 -29.520 93.030 ;
        RECT -26.730 92.310 -26.230 92.540 ;
        RECT -25.330 92.310 -24.330 92.540 ;
        RECT -31.920 91.820 -30.920 92.050 ;
        RECT -30.020 91.820 -29.520 92.050 ;
        RECT -26.730 91.330 -26.230 91.560 ;
        RECT -25.330 91.330 -24.330 91.560 ;
        RECT -31.920 90.840 -30.920 91.070 ;
        RECT -30.020 90.840 -29.520 91.070 ;
        RECT -28.585 90.270 -27.900 90.570 ;
        RECT -28.455 89.280 -28.135 90.270 ;
        RECT -38.355 88.960 -28.135 89.280 ;
        RECT -53.090 88.670 -47.080 88.940 ;
        RECT -56.990 85.790 -45.010 86.830 ;
        RECT -57.335 83.350 -56.975 83.520 ;
        RECT -32.335 83.350 -31.975 83.520 ;
        RECT -57.335 83.025 -56.235 83.350 ;
        RECT -57.335 82.995 -56.975 83.025 ;
        RECT -64.190 81.740 -63.960 82.735 ;
        RECT -60.630 81.840 -57.630 82.070 ;
        RECT -64.190 81.510 -63.180 81.740 ;
        RECT -64.190 81.250 -63.960 81.510 ;
        RECT -64.835 81.020 -63.950 81.250 ;
        RECT -64.190 80.760 -63.950 81.020 ;
        RECT -60.630 80.780 -57.630 81.010 ;
        RECT -64.190 80.530 -63.180 80.760 ;
        RECT -64.190 80.270 -63.950 80.530 ;
        RECT -60.630 80.290 -57.630 80.520 ;
        RECT -64.835 80.040 -63.950 80.270 ;
        RECT -64.190 79.780 -63.960 80.040 ;
        RECT -60.630 79.800 -57.630 80.030 ;
        RECT -64.190 79.550 -63.180 79.780 ;
        RECT -60.630 78.745 -57.630 78.975 ;
        RECT -56.560 78.250 -56.235 83.025 ;
        RECT -32.335 83.025 -31.235 83.350 ;
        RECT -32.335 82.995 -31.975 83.025 ;
        RECT -48.430 82.255 -47.105 82.435 ;
        RECT -44.330 82.255 -43.005 82.410 ;
        RECT -56.070 81.425 -54.570 81.655 ;
        RECT -48.430 81.315 -43.005 82.255 ;
        RECT -48.430 81.095 -47.105 81.315 ;
        RECT -44.330 81.070 -43.005 81.315 ;
        RECT -39.190 81.740 -38.960 82.735 ;
        RECT -35.630 81.840 -32.630 82.070 ;
        RECT -39.190 81.510 -38.180 81.740 ;
        RECT -39.190 81.250 -38.960 81.510 ;
        RECT -39.835 81.020 -38.950 81.250 ;
        RECT -39.190 80.760 -38.950 81.020 ;
        RECT -35.630 80.780 -32.630 81.010 ;
        RECT -39.190 80.530 -38.180 80.760 ;
        RECT -39.190 80.270 -38.950 80.530 ;
        RECT -35.630 80.290 -32.630 80.520 ;
        RECT -39.835 80.040 -38.950 80.270 ;
        RECT -39.190 79.780 -38.960 80.040 ;
        RECT -35.630 79.800 -32.630 80.030 ;
        RECT -39.190 79.550 -38.180 79.780 ;
        RECT -56.070 79.235 -54.570 79.465 ;
        RECT -35.630 78.745 -32.630 78.975 ;
        RECT -31.560 78.250 -31.235 83.025 ;
        RECT -31.070 81.425 -29.570 81.655 ;
        RECT -31.070 79.235 -29.570 79.465 ;
        RECT -67.785 77.975 -65.870 78.205 ;
        RECT -42.785 77.975 -40.870 78.205 ;
        RECT -67.785 77.225 -67.550 77.975 ;
        RECT -67.370 77.485 -63.185 77.715 ;
        RECT -67.785 76.995 -65.870 77.225 ;
        RECT -67.785 76.245 -67.550 76.995 ;
        RECT -59.410 76.745 -59.180 77.740 ;
        RECT -64.685 76.505 -63.185 76.735 ;
        RECT -60.190 76.515 -59.180 76.745 ;
        RECT -67.785 76.015 -65.870 76.245 ;
        RECT -67.785 76.010 -67.365 76.015 ;
        RECT -65.205 75.935 -64.915 76.330 ;
        RECT -59.410 76.255 -59.180 76.515 ;
        RECT -42.785 77.225 -42.550 77.975 ;
        RECT -42.370 77.485 -38.185 77.715 ;
        RECT -42.785 76.995 -40.870 77.225 ;
        RECT -65.750 75.665 -64.915 75.935 ;
        RECT -59.420 76.025 -58.535 76.255 ;
        RECT -42.785 76.245 -42.550 76.995 ;
        RECT -34.410 76.745 -34.180 77.740 ;
        RECT -39.685 76.505 -38.185 76.735 ;
        RECT -35.190 76.515 -34.180 76.745 ;
        RECT -59.420 75.765 -59.180 76.025 ;
        RECT -42.785 76.015 -40.870 76.245 ;
        RECT -42.785 76.010 -42.365 76.015 ;
        RECT -40.205 75.935 -39.915 76.330 ;
        RECT -34.410 76.255 -34.180 76.515 ;
        RECT -65.750 74.565 -65.480 75.665 ;
        RECT -65.205 75.535 -64.915 75.665 ;
        RECT -60.190 75.535 -59.180 75.765 ;
        RECT -59.420 75.275 -59.180 75.535 ;
        RECT -40.750 75.665 -39.915 75.935 ;
        RECT -34.420 76.025 -33.535 76.255 ;
        RECT -34.420 75.765 -34.180 76.025 ;
        RECT -59.420 75.045 -58.535 75.275 ;
        RECT -67.470 74.295 -65.480 74.565 ;
        RECT -69.500 69.350 -68.820 69.650 ;
        RECT -67.470 69.350 -67.200 74.295 ;
        RECT -65.340 73.830 -65.110 74.825 ;
        RECT -59.410 74.785 -59.180 75.045 ;
        RECT -60.190 74.555 -59.180 74.785 ;
        RECT -40.750 74.565 -40.480 75.665 ;
        RECT -40.205 75.535 -39.915 75.665 ;
        RECT -35.190 75.535 -34.180 75.765 ;
        RECT -34.420 75.275 -34.180 75.535 ;
        RECT -34.420 75.045 -33.535 75.275 ;
        RECT -42.470 74.295 -40.480 74.565 ;
        RECT -65.340 73.600 -63.830 73.830 ;
        RECT -65.340 73.340 -65.110 73.600 ;
        RECT -66.480 73.110 -65.100 73.340 ;
        RECT -65.340 72.850 -65.100 73.110 ;
        RECT -57.500 72.980 -55.585 73.210 ;
        RECT -65.340 72.620 -63.830 72.850 ;
        RECT -65.340 72.360 -65.100 72.620 ;
        RECT -60.185 72.490 -56.000 72.720 ;
        RECT -66.480 72.130 -65.100 72.360 ;
        RECT -55.820 72.230 -55.585 72.980 ;
        RECT -65.340 71.870 -65.110 72.130 ;
        RECT -57.500 72.000 -55.585 72.230 ;
        RECT -65.340 71.640 -63.830 71.870 ;
        RECT -60.185 71.510 -58.685 71.740 ;
        RECT -55.820 71.250 -55.585 72.000 ;
        RECT -57.500 71.020 -55.585 71.250 ;
        RECT -56.005 71.015 -55.585 71.020 ;
        RECT -65.750 70.730 -65.000 70.860 ;
        RECT -65.750 70.460 -57.710 70.730 ;
        RECT -65.750 70.210 -65.000 70.460 ;
        RECT -57.980 69.745 -57.710 70.460 ;
        RECT -42.470 70.340 -42.200 74.295 ;
        RECT -40.340 73.830 -40.110 74.825 ;
        RECT -34.410 74.785 -34.180 75.045 ;
        RECT -35.190 74.555 -34.180 74.785 ;
        RECT -40.340 73.600 -38.830 73.830 ;
        RECT -40.340 73.340 -40.110 73.600 ;
        RECT -41.480 73.110 -40.100 73.340 ;
        RECT -40.340 72.850 -40.100 73.110 ;
        RECT -32.500 72.980 -30.585 73.210 ;
        RECT -40.340 72.620 -38.830 72.850 ;
        RECT -40.340 72.360 -40.100 72.620 ;
        RECT -35.185 72.490 -31.000 72.720 ;
        RECT -41.480 72.130 -40.100 72.360 ;
        RECT -30.820 72.230 -30.585 72.980 ;
        RECT -40.340 71.870 -40.110 72.130 ;
        RECT -32.500 72.000 -30.585 72.230 ;
        RECT -40.340 71.640 -38.830 71.870 ;
        RECT -35.185 71.510 -33.685 71.740 ;
        RECT -30.820 71.250 -30.585 72.000 ;
        RECT -32.500 71.020 -30.585 71.250 ;
        RECT -31.005 71.015 -30.585 71.020 ;
        RECT -69.500 69.080 -67.200 69.350 ;
        RECT -46.040 69.140 -42.200 70.340 ;
        RECT -40.750 70.730 -40.000 70.860 ;
        RECT -40.750 70.460 -32.710 70.730 ;
        RECT -40.750 70.210 -40.000 70.460 ;
        RECT -32.980 69.745 -32.710 70.460 ;
        RECT -30.005 70.380 -29.715 70.705 ;
        RECT -30.310 69.975 -29.715 70.380 ;
        RECT -42.470 69.080 -42.200 69.140 ;
        RECT -69.500 68.930 -68.820 69.080 ;
        RECT -70.775 68.505 -70.090 68.735 ;
        RECT -58.770 68.505 -58.155 68.615 ;
        RECT -30.310 68.590 -30.135 69.975 ;
        RECT -70.775 68.045 -58.155 68.505 ;
        RECT -35.835 68.415 -30.135 68.590 ;
        RECT -29.880 68.565 -29.650 69.560 ;
        RECT -42.485 68.135 -41.485 68.365 ;
        RECT -38.945 68.135 -37.945 68.365 ;
        RECT -71.265 67.735 -70.975 68.040 ;
        RECT -58.770 68.030 -58.155 68.045 ;
        RECT -65.795 67.735 -65.110 67.825 ;
        RECT -71.265 67.540 -65.110 67.735 ;
        RECT -71.265 67.355 -70.975 67.540 ;
        RECT -65.795 67.535 -65.110 67.540 ;
        RECT -68.240 67.325 -67.555 67.400 ;
        RECT -57.280 67.325 -56.990 67.410 ;
        RECT -68.240 67.150 -56.990 67.325 ;
        RECT -68.240 67.110 -67.555 67.150 ;
        RECT -57.280 66.725 -56.990 67.150 ;
        RECT -56.040 66.535 -54.040 66.765 ;
        RECT -56.040 66.045 -54.040 66.275 ;
        RECT -42.485 66.070 -40.985 66.300 ;
        RECT -56.040 65.555 -54.040 65.785 ;
        RECT -42.485 65.580 -40.985 65.810 ;
        RECT -58.500 64.990 -57.500 65.220 ;
        RECT -42.485 65.090 -40.985 65.320 ;
        RECT -56.040 64.500 -54.040 64.730 ;
        RECT -42.485 64.525 -40.985 64.755 ;
        RECT -38.945 64.445 -37.945 64.675 ;
        RECT -42.485 64.035 -40.985 64.265 ;
        RECT -42.485 63.545 -40.985 63.775 ;
        RECT -38.945 63.465 -37.945 63.695 ;
        RECT -42.480 62.975 -40.980 63.205 ;
        RECT -67.810 62.700 -67.125 62.775 ;
        RECT -57.275 62.700 -56.985 62.755 ;
        RECT -67.810 62.525 -56.985 62.700 ;
        RECT -67.810 62.485 -67.125 62.525 ;
        RECT -57.275 62.070 -56.985 62.525 ;
        RECT -38.945 62.485 -37.945 62.715 ;
        RECT -56.035 62.010 -54.035 62.240 ;
        RECT -42.480 61.995 -40.980 62.225 ;
        RECT -56.035 61.520 -54.035 61.750 ;
        RECT -56.035 61.030 -54.035 61.260 ;
        RECT -40.260 61.110 -39.575 61.355 ;
        RECT -35.835 61.110 -35.660 68.415 ;
        RECT -29.880 68.335 -28.870 68.565 ;
        RECT -29.880 68.075 -29.650 68.335 ;
        RECT -30.525 67.845 -29.640 68.075 ;
        RECT -29.880 67.585 -29.640 67.845 ;
        RECT -29.880 67.355 -28.870 67.585 ;
        RECT -29.880 67.095 -29.640 67.355 ;
        RECT -30.525 66.865 -29.640 67.095 ;
        RECT -29.880 66.605 -29.650 66.865 ;
        RECT -29.880 66.375 -28.870 66.605 ;
        RECT -33.475 64.800 -31.560 65.030 ;
        RECT -33.475 64.050 -33.240 64.800 ;
        RECT -33.060 64.310 -28.875 64.540 ;
        RECT -33.475 63.820 -31.560 64.050 ;
        RECT -33.475 63.070 -33.240 63.820 ;
        RECT -30.375 63.330 -28.875 63.560 ;
        RECT -33.475 62.840 -31.560 63.070 ;
        RECT -33.475 62.835 -33.055 62.840 ;
        RECT 469.655 62.300 475.760 192.475 ;
        RECT -40.260 61.065 -35.660 61.110 ;
        RECT -39.805 60.935 -35.660 61.065 ;
        RECT -40.915 60.780 -40.230 60.870 ;
        RECT -58.495 60.465 -57.495 60.695 ;
        RECT -40.915 60.605 -32.385 60.780 ;
        RECT -40.915 60.580 -40.230 60.605 ;
        RECT -56.035 59.975 -54.035 60.205 ;
        RECT -41.400 59.510 -40.715 59.800 ;
        RECT -67.400 58.830 -64.010 59.280 ;
        RECT -66.445 58.400 -64.945 58.630 ;
        RECT -64.460 58.145 -64.010 58.830 ;
        RECT -39.425 58.855 -39.195 59.850 ;
        RECT -32.560 59.215 -32.385 60.605 ;
        RECT -32.805 58.985 -31.805 59.215 ;
        RECT -29.265 58.985 -28.265 59.215 ;
        RECT -39.425 58.625 -38.415 58.855 ;
        RECT -39.425 58.365 -39.195 58.625 ;
        RECT -59.020 58.145 -58.730 58.320 ;
        RECT -69.480 57.910 -68.480 58.140 ;
        RECT -64.460 57.695 -58.730 58.145 ;
        RECT -40.070 58.135 -39.185 58.365 ;
        RECT -39.425 57.875 -39.185 58.135 ;
        RECT -66.445 57.420 -64.945 57.650 ;
        RECT -59.020 57.635 -58.730 57.695 ;
        RECT -57.390 57.530 -54.390 57.760 ;
        RECT -39.425 57.645 -38.415 57.875 ;
        RECT -39.425 57.385 -39.185 57.645 ;
        RECT -69.480 56.930 -68.480 57.160 ;
        RECT -66.440 56.850 -64.940 57.080 ;
        RECT -57.390 57.040 -54.390 57.270 ;
        RECT -40.070 57.155 -39.185 57.385 ;
        RECT -39.425 56.895 -39.195 57.155 ;
        RECT -32.805 56.920 -31.305 57.150 ;
        RECT -66.440 56.360 -64.940 56.590 ;
        RECT -57.390 56.550 -54.390 56.780 ;
        RECT -39.425 56.665 -38.415 56.895 ;
        RECT -32.805 56.430 -31.305 56.660 ;
        RECT -69.480 55.950 -68.480 56.180 ;
        RECT -66.440 55.870 -64.940 56.100 ;
        RECT -57.390 55.985 -54.390 56.215 ;
        RECT -32.805 55.940 -31.305 56.170 ;
        RECT -66.440 55.305 -64.940 55.535 ;
        RECT -60.210 55.415 -59.210 55.645 ;
        RECT -57.390 55.495 -54.390 55.725 ;
        RECT -32.805 55.375 -31.305 55.605 ;
        RECT -66.440 54.815 -64.940 55.045 ;
        RECT -57.390 55.005 -54.390 55.235 ;
        RECT -43.020 55.090 -41.105 55.320 ;
        RECT -29.265 55.295 -28.265 55.525 ;
        RECT -66.440 54.325 -64.940 54.555 ;
        RECT -60.210 54.435 -59.210 54.665 ;
        RECT -43.020 54.340 -42.785 55.090 ;
        RECT -32.805 54.885 -31.305 55.115 ;
        RECT -42.605 54.600 -38.420 54.830 ;
        RECT -32.805 54.395 -31.305 54.625 ;
        RECT -0.785 54.610 0.435 62.285 ;
        RECT -57.390 53.945 -54.390 54.175 ;
        RECT -43.020 54.110 -41.105 54.340 ;
        RECT -29.265 54.315 -28.265 54.545 ;
        RECT -43.020 53.360 -42.785 54.110 ;
        RECT -39.920 53.620 -38.420 53.850 ;
        RECT -32.800 53.825 -31.300 54.055 ;
        RECT -43.020 53.130 -41.105 53.360 ;
        RECT -29.265 53.335 -28.265 53.565 ;
        RECT -43.020 53.125 -42.600 53.130 ;
        RECT -32.800 52.845 -31.300 53.075 ;
        RECT -71.415 52.480 -70.835 52.805 ;
        RECT -69.480 52.480 -68.480 52.490 ;
        RECT -71.415 52.265 -68.480 52.480 ;
        RECT -71.415 52.015 -70.835 52.265 ;
        RECT -69.480 52.260 -68.480 52.265 ;
        RECT -65.940 52.260 -64.940 52.490 ;
        RECT -0.330 52.365 -0.065 54.610 ;
        RECT 75.410 52.495 92.775 52.510 ;
        RECT 75.345 52.365 92.775 52.495 ;
        RECT -0.330 52.100 92.775 52.365 ;
        RECT 75.345 51.700 92.775 52.100 ;
        RECT 75.345 51.440 92.780 51.700 ;
        RECT 75.345 50.865 75.610 51.440 ;
        RECT 81.520 50.890 81.750 51.440 ;
        RECT 88.430 51.360 92.780 51.440 ;
        RECT 73.925 50.635 74.925 50.865 ;
        RECT 75.345 50.635 76.940 50.865 ;
        RECT 81.495 50.660 83.090 50.890 ;
        RECT 75.345 48.285 75.575 50.635 ;
        RECT 75.940 49.345 76.940 49.575 ;
        RECT 77.940 49.345 78.940 49.575 ;
        RECT 80.090 49.370 81.090 49.600 ;
        RECT 81.495 48.310 81.725 50.660 ;
        RECT 82.090 49.370 83.090 49.600 ;
        RECT 84.090 49.370 85.090 49.600 ;
        RECT 73.925 48.055 74.925 48.285 ;
        RECT 75.345 48.055 76.940 48.285 ;
        RECT 81.495 48.080 83.090 48.310 ;
        RECT 75.345 45.705 75.575 48.055 ;
        RECT 75.940 46.765 76.940 46.995 ;
        RECT 77.940 46.765 78.940 46.995 ;
        RECT 80.090 46.790 81.090 47.020 ;
        RECT 81.495 45.730 81.725 48.080 ;
        RECT 88.430 47.800 349.170 51.360 ;
        RECT 470.650 50.490 474.990 62.300 ;
        RECT 458.780 47.700 474.990 50.490 ;
        RECT 82.090 46.790 83.090 47.020 ;
        RECT 84.090 46.790 85.090 47.020 ;
        RECT 73.925 45.475 74.925 45.705 ;
        RECT 75.345 45.475 76.940 45.705 ;
        RECT 81.495 45.500 83.090 45.730 ;
        RECT 69.490 44.575 73.865 44.595 ;
        RECT 34.830 42.330 36.560 43.780 ;
        RECT 69.490 43.685 73.875 44.575 ;
        RECT -29.225 12.415 -27.695 13.820 ;
        RECT -3.065 13.550 7.285 14.080 ;
        RECT -46.955 7.520 -46.725 9.875 ;
        RECT -45.775 7.520 -45.545 9.875 ;
        RECT -44.595 7.520 -44.365 9.875 ;
        RECT -43.415 7.520 -43.185 9.875 ;
        RECT -42.235 7.520 -42.005 9.875 ;
        RECT -41.055 7.520 -40.825 9.875 ;
        RECT -39.875 7.520 -39.645 9.875 ;
        RECT -38.695 7.520 -38.465 9.875 ;
        RECT -36.865 7.520 -36.635 9.875 ;
        RECT -35.685 7.520 -35.455 9.875 ;
        RECT -34.505 7.520 -34.275 9.875 ;
        RECT -33.325 7.520 -33.095 9.875 ;
        RECT -31.495 7.520 -31.265 9.875 ;
        RECT -30.315 7.520 -30.085 9.875 ;
        RECT -28.710 7.605 -27.905 12.415 ;
        RECT -17.460 9.185 -17.230 10.185 ;
        RECT -16.480 9.185 -16.250 10.185 ;
        RECT -15.500 9.185 -15.270 10.185 ;
        RECT -13.210 9.185 -12.980 10.185 ;
        RECT -12.230 9.185 -12.000 10.185 ;
        RECT -11.250 9.185 -11.020 10.185 ;
        RECT -10.470 9.185 -10.240 10.185 ;
        RECT -9.980 8.965 -9.750 10.185 ;
        RECT -9.490 9.185 -9.260 10.185 ;
        RECT -9.000 8.965 -8.770 10.185 ;
        RECT -8.510 9.185 -8.280 10.185 ;
        RECT -8.020 8.965 -7.790 10.185 ;
        RECT -7.530 9.185 -7.300 10.185 ;
        RECT -7.040 8.965 -6.810 10.185 ;
        RECT -6.550 9.185 -6.320 10.185 ;
        RECT -9.980 8.735 -5.810 8.965 ;
        RECT -17.950 7.785 -17.720 8.285 ;
        RECT -17.460 7.785 -17.230 8.285 ;
        RECT -16.970 7.785 -16.740 8.285 ;
        RECT -16.480 7.785 -16.250 8.285 ;
        RECT -15.990 7.785 -15.760 8.285 ;
        RECT -15.500 7.785 -15.270 8.285 ;
        RECT -14.685 8.105 -14.025 8.325 ;
        RECT -47.530 7.150 -37.805 7.520 ;
        RECT -37.500 7.150 -32.450 7.520 ;
        RECT -32.145 7.150 -30.060 7.520 ;
        RECT -38.660 6.510 -38.430 7.150 ;
        RECT -38.855 6.280 -35.085 6.510 ;
        RECT -33.750 6.450 -33.520 7.150 ;
        RECT -66.585 3.835 -66.355 5.835 ;
        RECT -65.995 3.835 -65.765 5.835 ;
        RECT -65.405 3.835 -65.175 5.835 ;
        RECT -64.815 3.835 -64.585 5.835 ;
        RECT -64.225 3.835 -63.995 5.835 ;
        RECT -63.635 3.835 -63.405 5.835 ;
        RECT -63.045 3.835 -62.815 5.835 ;
        RECT -62.455 3.835 -62.225 5.835 ;
        RECT -61.865 3.835 -61.635 5.835 ;
        RECT -61.275 3.835 -61.045 5.835 ;
        RECT -60.685 3.835 -60.455 5.835 ;
        RECT -60.095 3.835 -59.865 5.835 ;
        RECT -59.505 3.835 -59.275 5.835 ;
        RECT -58.915 3.835 -58.685 5.835 ;
        RECT -58.325 3.835 -58.095 5.835 ;
        RECT -57.735 3.835 -57.505 5.835 ;
        RECT -57.145 3.835 -56.915 5.835 ;
        RECT -56.555 3.835 -56.325 5.835 ;
        RECT -55.965 3.835 -55.735 5.835 ;
        RECT -55.375 3.835 -55.145 5.835 ;
        RECT -54.785 3.835 -54.555 5.835 ;
        RECT -54.195 3.835 -53.965 5.835 ;
        RECT -53.605 3.835 -53.375 5.835 ;
        RECT -53.015 3.835 -52.785 5.835 ;
        RECT -52.425 3.835 -52.195 5.835 ;
        RECT -51.835 3.835 -51.605 5.835 ;
        RECT -51.245 3.835 -51.015 5.835 ;
        RECT -50.655 3.835 -50.425 5.835 ;
        RECT -50.065 3.835 -49.835 5.835 ;
        RECT -49.475 3.835 -49.245 5.835 ;
        RECT -48.885 3.835 -48.655 5.835 ;
        RECT -47.705 3.835 -47.475 5.835 ;
        RECT -46.525 3.835 -46.295 5.835 ;
        RECT -45.345 3.835 -45.115 5.835 ;
        RECT -44.165 3.835 -43.935 5.835 ;
        RECT -42.985 3.835 -42.755 5.835 ;
        RECT -41.805 3.835 -41.575 5.835 ;
        RECT -40.625 3.835 -40.395 5.835 ;
        RECT -39.445 3.835 -39.215 5.835 ;
        RECT -38.855 3.835 -38.625 6.280 ;
        RECT -38.265 3.835 -38.035 5.835 ;
        RECT -37.675 3.835 -37.445 6.280 ;
        RECT -37.085 3.835 -36.855 5.835 ;
        RECT -36.495 3.835 -36.265 6.280 ;
        RECT -35.905 3.835 -35.675 5.835 ;
        RECT -35.315 3.835 -35.085 6.280 ;
        RECT -34.135 6.220 -32.725 6.450 ;
        RECT -34.725 3.835 -34.495 5.835 ;
        RECT -34.135 3.835 -33.905 6.220 ;
        RECT -33.545 3.835 -33.315 5.835 ;
        RECT -32.955 3.835 -32.725 6.220 ;
        RECT -32.365 3.835 -32.135 5.835 ;
        RECT -31.775 3.835 -31.545 7.150 ;
        RECT -28.870 7.075 -27.870 7.605 ;
        RECT -21.060 7.490 -20.495 7.675 ;
        RECT -14.245 7.605 -14.025 8.105 ;
        RECT -13.700 7.785 -13.470 8.285 ;
        RECT -13.210 7.785 -12.980 8.285 ;
        RECT -12.720 7.785 -12.490 8.285 ;
        RECT -12.230 7.785 -12.000 8.285 ;
        RECT -11.740 7.785 -11.510 8.285 ;
        RECT -11.250 7.785 -11.020 8.285 ;
        RECT -10.470 7.605 -10.240 8.455 ;
        RECT -17.860 7.490 -15.300 7.510 ;
        RECT -21.060 7.305 -15.300 7.490 ;
        RECT -17.860 7.245 -15.300 7.305 ;
        RECT -14.245 7.385 -10.235 7.605 ;
        RECT -9.980 7.455 -9.750 8.735 ;
        RECT -9.490 7.455 -9.260 8.455 ;
        RECT -9.000 7.455 -8.770 8.735 ;
        RECT -8.510 7.455 -8.280 8.455 ;
        RECT -8.020 7.455 -7.790 8.735 ;
        RECT -7.530 7.455 -7.300 8.455 ;
        RECT -7.040 7.455 -6.810 8.735 ;
        RECT -6.550 7.455 -6.320 8.455 ;
        RECT -6.040 7.875 -5.810 8.735 ;
        RECT -3.065 7.875 -2.280 13.550 ;
        RECT 3.690 12.005 4.875 12.485 ;
        RECT 4.350 10.695 4.875 12.005 ;
        RECT 5.105 12.025 6.285 12.505 ;
        RECT 5.105 10.725 5.560 12.025 ;
        RECT 6.755 10.695 7.285 13.550 ;
        RECT 9.115 12.025 10.060 12.505 ;
        RECT 9.605 11.190 10.060 12.025 ;
        RECT 9.260 10.800 11.425 11.190 ;
        RECT 3.095 10.005 3.325 10.425 ;
        RECT 4.325 9.575 4.555 10.550 ;
        RECT 4.915 9.950 5.145 10.550 ;
        RECT 5.505 9.950 5.735 10.550 ;
        RECT 6.535 9.950 6.765 10.550 ;
        RECT 6.975 9.950 7.205 10.550 ;
        RECT 7.985 9.975 8.215 10.575 ;
        RECT 8.425 10.405 8.655 10.575 ;
        RECT 9.115 10.405 9.345 10.610 ;
        RECT 8.425 10.050 9.345 10.405 ;
        RECT 8.425 9.975 8.655 10.050 ;
        RECT 4.325 9.345 5.005 9.575 ;
        RECT 3.095 8.845 3.325 9.105 ;
        RECT -14.245 7.075 -14.025 7.385 ;
        RECT -28.870 6.855 -14.025 7.075 ;
        RECT -6.040 7.115 -2.280 7.875 ;
        RECT 2.055 8.460 3.325 8.845 ;
        RECT -28.870 6.760 -27.870 6.855 ;
        RECT -31.185 3.835 -30.955 5.835 ;
        RECT -13.700 5.710 -13.470 6.210 ;
        RECT -13.210 5.710 -12.980 6.210 ;
        RECT -12.720 5.710 -12.490 6.210 ;
        RECT -12.230 5.710 -12.000 6.210 ;
        RECT -11.740 5.710 -11.510 6.210 ;
        RECT -11.250 5.710 -11.020 6.210 ;
        RECT -9.980 5.260 -9.750 6.540 ;
        RECT -9.000 5.260 -8.770 6.540 ;
        RECT -8.020 5.260 -7.790 6.540 ;
        RECT -7.040 5.260 -6.810 6.540 ;
        RECT -6.040 5.260 -5.810 7.115 ;
        RECT -9.980 5.030 -5.810 5.260 ;
        RECT -13.210 3.810 -12.980 4.810 ;
        RECT -12.230 3.810 -12.000 4.810 ;
        RECT -11.250 3.810 -11.020 4.810 ;
        RECT -9.980 3.810 -9.750 5.030 ;
        RECT -9.000 3.810 -8.770 5.030 ;
        RECT -8.020 3.810 -7.790 5.030 ;
        RECT -7.040 3.810 -6.810 5.030 ;
        RECT -66.750 2.740 -30.400 3.605 ;
        RECT -63.795 -0.675 -61.360 2.740 ;
        RECT -55.995 -0.675 -53.560 2.740 ;
        RECT -50.030 -0.675 -47.595 2.740 ;
        RECT -44.115 -0.675 -41.680 2.740 ;
        RECT -39.045 -0.675 -36.610 2.740 ;
        RECT 2.055 1.540 2.440 8.460 ;
        RECT 3.095 8.265 3.325 8.460 ;
        RECT 4.775 8.125 5.005 9.345 ;
        RECT 7.495 9.270 7.950 9.665 ;
        RECT 8.190 9.495 8.665 9.625 ;
        RECT 9.115 9.525 9.345 10.050 ;
        RECT 10.295 10.010 10.525 10.610 ;
        RECT 11.475 10.010 11.705 10.610 ;
        RECT 12.910 10.005 13.140 10.425 ;
        RECT 14.455 10.005 14.685 10.425 ;
        RECT 23.035 10.065 23.265 11.065 ;
        RECT 24.015 10.065 24.245 11.065 ;
        RECT 24.995 10.065 25.225 11.065 ;
        RECT 27.285 10.065 27.515 11.065 ;
        RECT 28.265 10.065 28.495 11.065 ;
        RECT 29.245 10.065 29.475 11.065 ;
        RECT 30.025 10.065 30.255 11.065 ;
        RECT 30.515 9.845 30.745 11.065 ;
        RECT 31.005 10.065 31.235 11.065 ;
        RECT 31.495 9.845 31.725 11.065 ;
        RECT 31.985 10.065 32.215 11.065 ;
        RECT 32.475 9.845 32.705 11.065 ;
        RECT 32.965 10.065 33.195 11.065 ;
        RECT 33.455 9.845 33.685 11.065 ;
        RECT 33.945 10.065 34.175 11.065 ;
        RECT 35.400 10.395 36.145 42.330 ;
        RECT 36.445 40.085 38.175 41.535 ;
        RECT 30.515 9.615 34.685 9.845 ;
        RECT 8.190 9.285 8.970 9.495 ;
        RECT 9.115 9.295 9.970 9.525 ;
        RECT 5.655 8.495 5.885 9.095 ;
        RECT 6.535 8.495 6.765 9.095 ;
        RECT 5.585 8.125 5.945 8.275 ;
        RECT 6.470 8.125 6.830 8.270 ;
        RECT 7.540 8.195 7.770 9.095 ;
        RECT 7.980 8.195 8.210 9.095 ;
        RECT 4.775 7.895 6.830 8.125 ;
        RECT 5.585 7.870 5.945 7.895 ;
        RECT 5.600 7.855 5.930 7.870 ;
        RECT 6.470 7.865 6.830 7.895 ;
        RECT 6.485 7.850 6.815 7.865 ;
        RECT 8.800 7.265 8.970 9.285 ;
        RECT 9.740 8.195 9.970 9.295 ;
        RECT 12.910 8.265 13.140 9.105 ;
        RECT 14.455 8.265 14.685 9.105 ;
        RECT 23.035 8.665 23.265 9.165 ;
        RECT 24.015 8.665 24.245 9.165 ;
        RECT 24.995 8.665 25.225 9.165 ;
        RECT 25.810 8.985 26.470 9.205 ;
        RECT 26.250 8.485 26.470 8.985 ;
        RECT 27.285 8.665 27.515 9.165 ;
        RECT 28.265 8.665 28.495 9.165 ;
        RECT 29.245 8.665 29.475 9.165 ;
        RECT 30.025 8.485 30.255 9.335 ;
        RECT 26.250 8.265 30.260 8.485 ;
        RECT 30.515 8.335 30.745 9.615 ;
        RECT 31.005 8.335 31.235 9.335 ;
        RECT 31.495 8.335 31.725 9.615 ;
        RECT 31.985 8.335 32.215 9.335 ;
        RECT 32.475 8.335 32.705 9.615 ;
        RECT 32.965 8.335 33.195 9.335 ;
        RECT 33.455 8.335 33.685 9.615 ;
        RECT 33.945 8.335 34.175 9.335 ;
        RECT 34.455 8.350 34.685 9.615 ;
        RECT 35.270 9.225 36.515 10.395 ;
        RECT 36.705 8.400 37.300 40.085 ;
        RECT 44.980 33.480 45.210 37.480 ;
        RECT 53.560 33.480 53.790 37.480 ;
        RECT 60.790 33.480 61.020 37.480 ;
        RECT 45.160 28.215 45.390 32.215 ;
        RECT 53.740 28.215 53.970 32.215 ;
        RECT 69.490 29.820 70.400 43.685 ;
        RECT 72.735 43.680 73.875 43.685 ;
        RECT 75.395 34.850 75.625 45.475 ;
        RECT 78.630 44.240 80.585 44.470 ;
        RECT 81.130 43.025 81.980 43.715 ;
        RECT 74.985 33.780 76.055 34.850 ;
        RECT 81.250 33.115 81.940 43.025 ;
        RECT 81.135 32.220 82.030 33.115 ;
        RECT 96.005 33.100 98.215 35.425 ;
        RECT 114.695 33.330 116.515 35.580 ;
        RECT 69.330 28.515 70.650 29.820 ;
        RECT 62.320 23.215 62.550 27.215 ;
        RECT 93.955 26.080 95.840 27.865 ;
        RECT 38.650 8.930 38.880 11.285 ;
        RECT 39.830 8.930 40.060 11.285 ;
        RECT 41.660 8.930 41.890 11.285 ;
        RECT 42.840 8.930 43.070 11.285 ;
        RECT 44.020 8.930 44.250 11.285 ;
        RECT 45.200 8.930 45.430 11.285 ;
        RECT 47.030 8.930 47.260 11.285 ;
        RECT 48.210 8.930 48.440 11.285 ;
        RECT 49.390 8.930 49.620 11.285 ;
        RECT 50.570 8.930 50.800 11.285 ;
        RECT 51.750 8.930 51.980 11.285 ;
        RECT 52.930 8.930 53.160 11.285 ;
        RECT 54.110 8.930 54.340 11.285 ;
        RECT 55.290 8.930 55.520 11.285 ;
        RECT 38.625 8.560 40.710 8.930 ;
        RECT 41.015 8.560 46.065 8.930 ;
        RECT 46.370 8.560 56.095 8.930 ;
        RECT 36.685 8.350 37.350 8.400 ;
        RECT 19.950 7.955 20.530 8.190 ;
        RECT 26.250 7.955 26.470 8.265 ;
        RECT 19.950 7.735 26.470 7.955 ;
        RECT 34.455 8.120 37.350 8.350 ;
        RECT 19.950 7.495 20.530 7.735 ;
        RECT 7.540 7.035 8.970 7.265 ;
        RECT 5.600 6.440 5.930 6.455 ;
        RECT 6.485 6.445 6.815 6.460 ;
        RECT 5.585 6.415 5.945 6.440 ;
        RECT 6.470 6.415 6.830 6.445 ;
        RECT 4.775 6.185 6.830 6.415 ;
        RECT 3.095 5.205 3.325 6.045 ;
        RECT 4.775 4.965 5.005 6.185 ;
        RECT 5.585 6.035 5.945 6.185 ;
        RECT 6.470 6.040 6.830 6.185 ;
        RECT 5.655 5.215 5.885 5.815 ;
        RECT 6.535 5.215 6.765 5.815 ;
        RECT 7.540 5.215 7.770 7.035 ;
        RECT 27.285 6.590 27.515 7.090 ;
        RECT 28.265 6.590 28.495 7.090 ;
        RECT 29.245 6.590 29.475 7.090 ;
        RECT 30.515 6.140 30.745 7.420 ;
        RECT 31.495 6.140 31.725 7.420 ;
        RECT 32.475 6.140 32.705 7.420 ;
        RECT 33.455 6.140 33.685 7.420 ;
        RECT 34.455 6.140 34.685 8.120 ;
        RECT 36.685 7.810 37.350 8.120 ;
        RECT 35.305 6.775 36.350 7.770 ;
        RECT 7.980 5.215 8.210 6.115 ;
        RECT 4.325 4.735 5.005 4.965 ;
        RECT 3.095 3.885 3.325 4.305 ;
        RECT 4.325 3.760 4.555 4.735 ;
        RECT 8.190 4.685 8.665 5.025 ;
        RECT 9.740 5.015 9.970 6.115 ;
        RECT 12.910 5.205 13.140 6.045 ;
        RECT 14.455 5.205 14.685 6.045 ;
        RECT 30.515 5.910 34.685 6.140 ;
        RECT 9.115 4.785 9.970 5.015 ;
        RECT 17.815 4.865 18.625 5.195 ;
        RECT 4.915 3.760 5.145 4.360 ;
        RECT 5.505 3.760 5.735 4.360 ;
        RECT 6.535 3.760 6.765 4.360 ;
        RECT 6.975 3.760 7.205 4.360 ;
        RECT 7.985 3.735 8.215 4.335 ;
        RECT 8.425 4.260 8.655 4.335 ;
        RECT 9.115 4.260 9.345 4.785 ;
        RECT 17.815 4.645 19.060 4.865 ;
        RECT 27.285 4.690 27.515 5.690 ;
        RECT 28.265 4.690 28.495 5.690 ;
        RECT 29.245 4.690 29.475 5.690 ;
        RECT 30.515 4.690 30.745 5.910 ;
        RECT 31.495 4.690 31.725 5.910 ;
        RECT 32.475 4.690 32.705 5.910 ;
        RECT 33.455 4.690 33.685 5.910 ;
        RECT 17.815 4.425 18.625 4.645 ;
        RECT 8.425 3.905 9.345 4.260 ;
        RECT 8.425 3.735 8.655 3.905 ;
        RECT 9.115 3.700 9.345 3.905 ;
        RECT 10.295 3.700 10.525 4.300 ;
        RECT 11.475 3.700 11.705 4.300 ;
        RECT 12.910 3.885 13.140 4.305 ;
        RECT 14.455 3.885 14.685 4.305 ;
        RECT 4.350 2.305 4.875 3.615 ;
        RECT 3.690 1.825 4.875 2.305 ;
        RECT 5.105 2.285 5.560 3.585 ;
        RECT 5.105 1.810 6.285 2.285 ;
        RECT 5.100 1.805 6.285 1.810 ;
        RECT 5.100 1.540 5.560 1.805 ;
        RECT 2.055 1.155 5.560 1.540 ;
        RECT 6.755 0.530 7.285 3.615 ;
        RECT 9.260 3.120 11.425 3.510 ;
        RECT 9.605 2.285 10.060 3.120 ;
        RECT 9.115 1.805 10.060 2.285 ;
        RECT -12.605 0.000 7.285 0.530 ;
        RECT -65.985 -2.265 -35.815 -0.675 ;
        RECT -30.295 -1.890 -27.535 -1.380 ;
        RECT -127.765 -5.250 -125.825 -3.270 ;
        RECT -134.535 -55.765 -129.915 -54.900 ;
        RECT -139.045 -58.525 -129.915 -55.765 ;
        RECT -139.045 -214.280 -136.285 -58.525 ;
        RECT -134.535 -59.520 -129.915 -58.525 ;
        RECT -127.505 -70.540 -126.095 -5.250 ;
        RECT -64.325 -54.695 -59.620 -2.265 ;
        RECT -121.240 -59.400 -59.615 -54.695 ;
        RECT -129.655 -74.380 -124.350 -70.540 ;
        RECT -127.505 -113.895 -126.095 -74.380 ;
        RECT -64.325 -74.845 -59.620 -59.400 ;
        RECT -53.070 -74.845 -48.365 -2.265 ;
        RECT -44.675 -74.845 -39.970 -2.265 ;
        RECT -29.880 -4.785 -29.000 -3.920 ;
        RECT -27.720 -4.365 -27.535 -1.890 ;
        RECT -24.800 -2.675 -24.570 -1.675 ;
        RECT -23.820 -2.675 -23.590 -1.675 ;
        RECT -22.840 -2.675 -22.610 -1.675 ;
        RECT -20.550 -2.675 -20.320 -1.675 ;
        RECT -19.570 -2.675 -19.340 -1.675 ;
        RECT -18.590 -2.675 -18.360 -1.675 ;
        RECT -17.810 -2.675 -17.580 -1.675 ;
        RECT -17.320 -2.895 -17.090 -1.675 ;
        RECT -16.830 -2.675 -16.600 -1.675 ;
        RECT -16.340 -2.895 -16.110 -1.675 ;
        RECT -15.850 -2.675 -15.620 -1.675 ;
        RECT -15.360 -2.895 -15.130 -1.675 ;
        RECT -14.870 -2.675 -14.640 -1.675 ;
        RECT -14.380 -2.895 -14.150 -1.675 ;
        RECT -13.890 -2.675 -13.660 -1.675 ;
        RECT -17.320 -3.125 -13.150 -2.895 ;
        RECT -25.290 -4.075 -25.060 -3.575 ;
        RECT -24.800 -4.075 -24.570 -3.575 ;
        RECT -24.310 -4.075 -24.080 -3.575 ;
        RECT -23.820 -4.075 -23.590 -3.575 ;
        RECT -23.330 -4.075 -23.100 -3.575 ;
        RECT -22.840 -4.075 -22.610 -3.575 ;
        RECT -22.025 -3.755 -21.365 -3.535 ;
        RECT -21.585 -4.255 -21.365 -3.755 ;
        RECT -21.040 -4.075 -20.810 -3.575 ;
        RECT -20.550 -4.075 -20.320 -3.575 ;
        RECT -20.060 -4.075 -19.830 -3.575 ;
        RECT -19.570 -4.075 -19.340 -3.575 ;
        RECT -19.080 -4.075 -18.850 -3.575 ;
        RECT -18.590 -4.075 -18.360 -3.575 ;
        RECT -17.810 -4.255 -17.580 -3.405 ;
        RECT -25.280 -4.365 -22.665 -4.305 ;
        RECT -27.720 -4.550 -22.665 -4.365 ;
        RECT -25.280 -4.610 -22.665 -4.550 ;
        RECT -21.585 -4.475 -17.575 -4.255 ;
        RECT -17.320 -4.405 -17.090 -3.125 ;
        RECT -16.830 -4.405 -16.600 -3.405 ;
        RECT -16.340 -4.405 -16.110 -3.125 ;
        RECT -15.850 -4.405 -15.620 -3.405 ;
        RECT -15.360 -4.405 -15.130 -3.125 ;
        RECT -14.870 -4.405 -14.640 -3.405 ;
        RECT -14.380 -4.405 -14.150 -3.125 ;
        RECT -13.890 -4.405 -13.660 -3.405 ;
        RECT -13.380 -3.895 -13.150 -3.125 ;
        RECT -12.605 -3.325 -12.075 0.000 ;
        RECT -12.605 -3.895 -12.110 -3.325 ;
        RECT -21.585 -4.785 -21.365 -4.475 ;
        RECT -29.880 -5.005 -21.365 -4.785 ;
        RECT -13.380 -4.620 -12.110 -3.895 ;
        RECT -29.880 -5.025 -29.000 -5.005 ;
        RECT -20.925 -5.250 -20.310 -4.945 ;
        RECT -21.585 -5.470 -17.575 -5.250 ;
        RECT -21.585 -5.970 -21.365 -5.470 ;
        RECT -26.245 -6.190 -21.365 -5.970 ;
        RECT -21.040 -6.150 -20.810 -5.650 ;
        RECT -20.550 -6.150 -20.320 -5.650 ;
        RECT -20.060 -6.150 -19.830 -5.650 ;
        RECT -19.570 -6.150 -19.340 -5.650 ;
        RECT -19.080 -6.150 -18.850 -5.650 ;
        RECT -18.590 -6.150 -18.360 -5.650 ;
        RECT -17.810 -6.320 -17.580 -5.470 ;
        RECT -17.320 -6.600 -17.090 -5.320 ;
        RECT -16.830 -6.320 -16.600 -5.320 ;
        RECT -16.340 -6.600 -16.110 -5.320 ;
        RECT -15.850 -6.320 -15.620 -5.320 ;
        RECT -15.360 -6.600 -15.130 -5.320 ;
        RECT -14.870 -6.320 -14.640 -5.320 ;
        RECT -14.380 -6.600 -14.150 -5.320 ;
        RECT -13.890 -6.320 -13.660 -5.320 ;
        RECT -13.380 -6.600 -13.150 -4.620 ;
        RECT 18.840 -5.495 19.060 4.645 ;
        RECT 23.110 -3.385 23.340 -2.385 ;
        RECT 24.090 -3.385 24.320 -2.385 ;
        RECT 25.070 -3.385 25.300 -2.385 ;
        RECT 27.360 -3.385 27.590 -2.385 ;
        RECT 28.340 -3.385 28.570 -2.385 ;
        RECT 29.320 -3.385 29.550 -2.385 ;
        RECT 30.100 -3.385 30.330 -2.385 ;
        RECT 30.590 -3.605 30.820 -2.385 ;
        RECT 31.080 -3.385 31.310 -2.385 ;
        RECT 31.570 -3.605 31.800 -2.385 ;
        RECT 32.060 -3.385 32.290 -2.385 ;
        RECT 32.550 -3.605 32.780 -2.385 ;
        RECT 33.040 -3.385 33.270 -2.385 ;
        RECT 33.530 -3.605 33.760 -2.385 ;
        RECT 34.020 -3.385 34.250 -2.385 ;
        RECT 30.590 -3.835 34.760 -3.605 ;
        RECT 23.110 -4.785 23.340 -4.285 ;
        RECT 24.090 -4.785 24.320 -4.285 ;
        RECT 25.070 -4.785 25.300 -4.285 ;
        RECT 25.885 -4.465 26.545 -4.245 ;
        RECT 26.325 -4.965 26.545 -4.465 ;
        RECT 27.360 -4.785 27.590 -4.285 ;
        RECT 28.340 -4.785 28.570 -4.285 ;
        RECT 29.320 -4.785 29.550 -4.285 ;
        RECT 30.100 -4.965 30.330 -4.115 ;
        RECT 26.325 -5.185 30.335 -4.965 ;
        RECT 30.590 -5.115 30.820 -3.835 ;
        RECT 31.080 -5.115 31.310 -4.115 ;
        RECT 31.570 -5.115 31.800 -3.835 ;
        RECT 32.060 -5.115 32.290 -4.115 ;
        RECT 32.550 -5.115 32.780 -3.835 ;
        RECT 33.040 -5.115 33.270 -4.115 ;
        RECT 33.530 -5.115 33.760 -3.835 ;
        RECT 34.020 -5.115 34.250 -4.115 ;
        RECT 34.530 -5.100 34.760 -3.835 ;
        RECT 35.655 -5.100 36.150 6.775 ;
        RECT 40.110 5.245 40.340 8.560 ;
        RECT 42.085 7.860 42.315 8.560 ;
        RECT 46.995 7.920 47.225 8.560 ;
        RECT 41.290 7.630 42.700 7.860 ;
        RECT 41.290 5.245 41.520 7.630 ;
        RECT 42.470 5.245 42.700 7.630 ;
        RECT 43.650 7.690 47.420 7.920 ;
        RECT 43.650 5.245 43.880 7.690 ;
        RECT 44.830 5.245 45.060 7.690 ;
        RECT 46.010 5.245 46.240 7.690 ;
        RECT 47.190 5.245 47.420 7.690 ;
        RECT 38.445 -4.850 38.675 -2.495 ;
        RECT 39.625 -4.850 39.855 -2.495 ;
        RECT 41.455 -4.850 41.685 -2.495 ;
        RECT 42.635 -4.850 42.865 -2.495 ;
        RECT 43.815 -4.850 44.045 -2.495 ;
        RECT 44.995 -4.850 45.225 -2.495 ;
        RECT 46.825 -4.850 47.055 -2.495 ;
        RECT 48.005 -4.850 48.235 -2.495 ;
        RECT 49.185 -4.850 49.415 -2.495 ;
        RECT 50.365 -4.850 50.595 -2.495 ;
        RECT 51.545 -4.850 51.775 -2.495 ;
        RECT 52.725 -4.850 52.955 -2.495 ;
        RECT 53.905 -4.850 54.135 -2.495 ;
        RECT 55.085 -4.850 55.315 -2.495 ;
        RECT 94.305 -2.970 95.765 26.080 ;
        RECT 96.705 13.780 97.350 33.100 ;
        RECT 99.430 15.890 99.660 16.890 ;
        RECT 100.410 15.890 100.640 16.890 ;
        RECT 101.390 15.890 101.620 16.890 ;
        RECT 103.680 15.890 103.910 16.890 ;
        RECT 104.660 15.890 104.890 16.890 ;
        RECT 105.640 15.890 105.870 16.890 ;
        RECT 106.420 15.890 106.650 16.890 ;
        RECT 106.910 15.670 107.140 16.890 ;
        RECT 107.400 15.890 107.630 16.890 ;
        RECT 107.890 15.670 108.120 16.890 ;
        RECT 108.380 15.890 108.610 16.890 ;
        RECT 108.870 15.670 109.100 16.890 ;
        RECT 109.360 15.890 109.590 16.890 ;
        RECT 109.850 15.670 110.080 16.890 ;
        RECT 110.340 15.890 110.570 16.890 ;
        RECT 106.910 15.440 111.080 15.670 ;
        RECT 99.430 14.490 99.660 14.990 ;
        RECT 100.410 14.490 100.640 14.990 ;
        RECT 101.390 14.490 101.620 14.990 ;
        RECT 102.205 14.810 102.865 15.030 ;
        RECT 102.645 14.310 102.865 14.810 ;
        RECT 103.680 14.490 103.910 14.990 ;
        RECT 104.660 14.490 104.890 14.990 ;
        RECT 105.640 14.490 105.870 14.990 ;
        RECT 106.420 14.310 106.650 15.160 ;
        RECT 102.645 14.090 106.655 14.310 ;
        RECT 106.910 14.160 107.140 15.440 ;
        RECT 107.400 14.160 107.630 15.160 ;
        RECT 107.890 14.160 108.120 15.440 ;
        RECT 108.380 14.160 108.610 15.160 ;
        RECT 108.870 14.160 109.100 15.440 ;
        RECT 109.360 14.160 109.590 15.160 ;
        RECT 109.850 14.160 110.080 15.440 ;
        RECT 110.340 14.160 110.570 15.160 ;
        RECT 110.850 14.375 111.080 15.440 ;
        RECT 111.580 14.375 112.770 14.500 ;
        RECT 102.645 13.780 102.865 14.090 ;
        RECT 96.705 13.560 102.865 13.780 ;
        RECT 110.850 13.725 112.770 14.375 ;
        RECT 96.705 13.500 97.350 13.560 ;
        RECT 103.680 12.415 103.910 12.915 ;
        RECT 104.660 12.415 104.890 12.915 ;
        RECT 105.640 12.415 105.870 12.915 ;
        RECT 106.910 11.965 107.140 13.245 ;
        RECT 107.890 11.965 108.120 13.245 ;
        RECT 108.870 11.965 109.100 13.245 ;
        RECT 109.850 11.965 110.080 13.245 ;
        RECT 110.850 11.965 111.080 13.725 ;
        RECT 111.580 13.555 112.770 13.725 ;
        RECT 106.910 11.735 111.080 11.965 ;
        RECT 103.680 10.515 103.910 11.515 ;
        RECT 104.660 10.515 104.890 11.515 ;
        RECT 105.640 10.515 105.870 11.515 ;
        RECT 106.910 10.515 107.140 11.735 ;
        RECT 107.890 10.515 108.120 11.735 ;
        RECT 108.870 10.515 109.100 11.735 ;
        RECT 109.850 10.515 110.080 11.735 ;
        RECT 100.290 -0.860 100.520 0.140 ;
        RECT 101.270 -0.860 101.500 0.140 ;
        RECT 102.250 -0.860 102.480 0.140 ;
        RECT 104.540 -0.860 104.770 0.140 ;
        RECT 105.520 -0.860 105.750 0.140 ;
        RECT 106.500 -0.860 106.730 0.140 ;
        RECT 107.280 -0.860 107.510 0.140 ;
        RECT 107.770 -1.080 108.000 0.140 ;
        RECT 108.260 -0.860 108.490 0.140 ;
        RECT 108.750 -1.080 108.980 0.140 ;
        RECT 109.240 -0.860 109.470 0.140 ;
        RECT 109.730 -1.080 109.960 0.140 ;
        RECT 110.220 -0.860 110.450 0.140 ;
        RECT 110.710 -1.080 110.940 0.140 ;
        RECT 111.200 -0.860 111.430 0.140 ;
        RECT 107.770 -1.310 111.940 -1.080 ;
        RECT 100.290 -2.260 100.520 -1.760 ;
        RECT 101.270 -2.260 101.500 -1.760 ;
        RECT 102.250 -2.260 102.480 -1.760 ;
        RECT 103.065 -1.940 103.725 -1.720 ;
        RECT 103.505 -2.440 103.725 -1.940 ;
        RECT 104.540 -2.260 104.770 -1.760 ;
        RECT 105.520 -2.260 105.750 -1.760 ;
        RECT 106.500 -2.260 106.730 -1.760 ;
        RECT 107.280 -2.440 107.510 -1.590 ;
        RECT 103.505 -2.660 107.515 -2.440 ;
        RECT 107.770 -2.590 108.000 -1.310 ;
        RECT 108.260 -2.590 108.490 -1.590 ;
        RECT 108.750 -2.590 108.980 -1.310 ;
        RECT 109.240 -2.590 109.470 -1.590 ;
        RECT 109.730 -2.590 109.960 -1.310 ;
        RECT 110.220 -2.590 110.450 -1.590 ;
        RECT 110.710 -2.590 110.940 -1.310 ;
        RECT 111.200 -2.590 111.430 -1.590 ;
        RECT 111.710 -1.725 111.940 -1.310 ;
        RECT 111.710 -1.765 112.565 -1.725 ;
        RECT 115.230 -1.765 116.085 33.330 ;
        RECT 131.620 15.085 192.950 15.765 ;
        RECT 125.305 11.475 126.665 11.860 ;
        RECT 129.735 11.475 130.750 11.785 ;
        RECT 125.305 10.620 130.750 11.475 ;
        RECT 125.305 10.425 126.665 10.620 ;
        RECT 129.735 10.460 130.750 10.620 ;
        RECT 131.620 5.470 132.300 15.085 ;
        RECT 138.005 12.855 160.555 13.260 ;
        RECT 138.005 11.390 138.410 12.855 ;
        RECT 136.360 11.130 138.410 11.390 ;
        RECT 138.955 11.130 139.760 11.200 ;
        RECT 136.360 10.855 139.760 11.130 ;
        RECT 145.955 10.895 146.345 10.975 ;
        RECT 136.360 10.725 138.260 10.855 ;
        RECT 138.955 10.805 139.760 10.855 ;
        RECT 145.375 10.765 146.345 10.895 ;
        RECT 140.080 10.620 146.345 10.765 ;
        RECT 140.080 7.025 140.270 10.620 ;
        RECT 140.515 9.285 140.745 10.285 ;
        RECT 142.095 9.285 142.325 10.620 ;
        RECT 143.675 9.285 143.905 10.285 ;
        RECT 144.325 9.310 144.555 10.620 ;
        RECT 152.410 10.480 152.640 12.480 ;
        RECT 153.990 10.480 154.220 12.480 ;
        RECT 160.150 11.165 160.555 12.855 ;
        RECT 160.150 10.765 164.045 11.165 ;
        RECT 170.230 10.860 170.620 10.940 ;
        RECT 160.150 10.760 163.400 10.765 ;
        RECT 169.650 10.730 170.620 10.860 ;
        RECT 164.355 10.585 170.620 10.730 ;
        RECT 176.085 10.590 176.315 12.590 ;
        RECT 177.665 10.590 177.895 12.590 ;
        RECT 145.905 9.310 146.135 10.310 ;
        RECT 140.515 7.025 140.745 8.340 ;
        RECT 142.095 7.340 142.325 8.340 ;
        RECT 143.675 7.025 143.905 8.340 ;
        RECT 144.325 7.340 144.555 8.340 ;
        RECT 145.905 7.035 146.135 8.340 ;
        RECT 152.410 7.200 152.640 9.200 ;
        RECT 153.990 7.200 154.220 9.200 ;
        RECT 155.570 7.200 155.800 9.200 ;
        RECT 157.150 7.200 157.380 9.200 ;
        RECT 146.300 7.035 147.075 7.110 ;
        RECT 145.905 7.025 147.075 7.035 ;
        RECT 140.080 6.840 147.075 7.025 ;
        RECT 140.080 6.480 146.080 6.840 ;
        RECT 146.300 6.780 147.075 6.840 ;
        RECT 164.355 6.990 164.545 10.585 ;
        RECT 164.790 9.250 165.020 10.250 ;
        RECT 166.370 9.250 166.600 10.585 ;
        RECT 167.950 9.250 168.180 10.250 ;
        RECT 168.600 9.275 168.830 10.585 ;
        RECT 184.690 10.375 184.920 12.375 ;
        RECT 186.270 10.375 186.500 12.375 ;
        RECT 170.180 9.275 170.410 10.275 ;
        RECT 192.270 10.065 192.950 15.085 ;
        RECT 199.725 15.015 221.010 15.300 ;
        RECT 196.390 13.675 196.620 14.675 ;
        RECT 197.370 13.675 197.600 14.675 ;
        RECT 198.350 13.675 198.580 14.675 ;
        RECT 199.725 13.410 200.010 15.015 ;
        RECT 200.800 13.675 201.030 14.675 ;
        RECT 201.780 13.675 202.010 14.675 ;
        RECT 202.760 13.675 202.990 14.675 ;
        RECT 203.855 14.100 204.085 14.600 ;
        RECT 204.345 14.100 204.575 14.600 ;
        RECT 204.835 14.100 205.065 14.600 ;
        RECT 205.325 14.100 205.555 14.600 ;
        RECT 205.815 14.100 206.045 14.600 ;
        RECT 206.305 14.100 206.535 14.600 ;
        RECT 206.795 14.100 207.025 14.600 ;
        RECT 207.285 14.100 207.515 14.600 ;
        RECT 209.515 13.675 209.745 14.675 ;
        RECT 210.495 13.675 210.725 14.675 ;
        RECT 211.475 13.675 211.705 14.675 ;
        RECT 203.870 13.410 204.715 13.460 ;
        RECT 196.390 12.275 196.620 12.775 ;
        RECT 197.370 12.275 197.600 12.775 ;
        RECT 198.350 12.275 198.580 12.775 ;
        RECT 199.020 12.620 199.320 13.280 ;
        RECT 199.725 13.125 204.715 13.410 ;
        RECT 213.225 13.410 213.510 14.585 ;
        RECT 214.300 13.675 214.530 14.675 ;
        RECT 215.280 13.675 215.510 14.675 ;
        RECT 216.260 13.675 216.490 14.675 ;
        RECT 217.355 14.100 217.585 14.600 ;
        RECT 217.830 14.410 218.085 15.015 ;
        RECT 217.845 14.100 218.075 14.410 ;
        RECT 218.335 14.100 218.565 14.600 ;
        RECT 218.800 14.410 219.055 15.015 ;
        RECT 218.825 14.100 219.055 14.410 ;
        RECT 219.315 14.100 219.545 14.600 ;
        RECT 219.800 14.315 220.055 15.015 ;
        RECT 220.760 14.600 221.010 15.015 ;
        RECT 219.805 14.100 220.035 14.315 ;
        RECT 220.295 14.100 220.525 14.600 ;
        RECT 220.760 14.440 221.015 14.600 ;
        RECT 220.785 14.100 221.015 14.440 ;
        RECT 223.015 13.675 223.245 14.675 ;
        RECT 223.995 13.675 224.225 14.675 ;
        RECT 224.975 13.675 225.205 14.675 ;
        RECT 217.370 13.410 218.215 13.460 ;
        RECT 203.870 13.090 204.715 13.125 ;
        RECT 199.020 11.480 199.310 12.620 ;
        RECT 200.800 12.275 201.030 12.775 ;
        RECT 201.780 12.275 202.010 12.775 ;
        RECT 202.760 12.275 202.990 12.775 ;
        RECT 203.855 12.025 204.085 12.525 ;
        RECT 204.345 12.025 204.575 12.525 ;
        RECT 204.835 12.025 205.065 12.525 ;
        RECT 205.325 12.025 205.555 12.525 ;
        RECT 205.815 12.025 206.045 12.525 ;
        RECT 206.305 12.025 206.535 12.525 ;
        RECT 206.795 12.025 207.025 12.525 ;
        RECT 207.270 12.025 207.515 12.525 ;
        RECT 209.515 12.275 209.745 12.775 ;
        RECT 210.495 12.275 210.725 12.775 ;
        RECT 211.475 12.275 211.705 12.775 ;
        RECT 212.105 12.725 212.405 13.160 ;
        RECT 212.100 12.500 212.405 12.725 ;
        RECT 204.360 11.540 204.570 12.025 ;
        RECT 205.340 11.540 205.550 12.025 ;
        RECT 206.315 11.540 206.525 12.025 ;
        RECT 207.270 11.540 207.500 12.025 ;
        RECT 198.815 11.180 199.475 11.480 ;
        RECT 203.700 11.310 207.500 11.540 ;
        RECT 203.700 10.480 203.930 11.310 ;
        RECT 207.835 10.750 208.495 11.050 ;
        RECT 199.875 10.475 203.930 10.480 ;
        RECT 199.835 10.250 203.930 10.475 ;
        RECT 164.790 6.990 165.020 8.305 ;
        RECT 166.370 7.305 166.600 8.305 ;
        RECT 167.950 6.990 168.180 8.305 ;
        RECT 168.600 7.305 168.830 8.305 ;
        RECT 170.180 7.000 170.410 8.305 ;
        RECT 176.085 7.310 176.315 9.310 ;
        RECT 177.665 7.310 177.895 9.310 ;
        RECT 179.245 7.310 179.475 9.310 ;
        RECT 180.825 7.310 181.055 9.310 ;
        RECT 184.690 7.095 184.920 9.095 ;
        RECT 186.270 7.095 186.500 9.095 ;
        RECT 187.850 7.095 188.080 9.095 ;
        RECT 189.430 7.095 189.660 9.095 ;
        RECT 192.145 8.775 193.105 10.065 ;
        RECT 199.835 8.875 200.065 10.250 ;
        RECT 200.315 9.235 200.545 9.735 ;
        RECT 200.805 9.235 201.035 9.735 ;
        RECT 201.295 9.235 201.525 9.735 ;
        RECT 201.785 9.235 202.015 9.735 ;
        RECT 202.275 9.235 202.505 9.735 ;
        RECT 202.765 9.235 202.995 9.735 ;
        RECT 203.255 9.235 203.485 9.735 ;
        RECT 203.745 9.235 203.975 9.735 ;
        RECT 204.840 8.985 205.070 9.485 ;
        RECT 205.820 8.985 206.050 9.485 ;
        RECT 206.800 8.985 207.030 9.485 ;
        RECT 208.050 8.930 208.350 10.750 ;
        RECT 209.025 8.985 209.255 9.485 ;
        RECT 210.005 8.985 210.235 9.485 ;
        RECT 210.985 8.985 211.215 9.485 ;
        RECT 199.835 8.575 200.605 8.875 ;
        RECT 212.100 8.760 212.400 12.500 ;
        RECT 212.680 11.045 212.980 13.285 ;
        RECT 213.225 13.125 218.215 13.410 ;
        RECT 217.370 13.090 218.215 13.125 ;
        RECT 255.040 12.815 255.270 15.170 ;
        RECT 256.220 12.815 256.450 15.170 ;
        RECT 258.050 12.815 258.280 15.170 ;
        RECT 259.230 12.815 259.460 15.170 ;
        RECT 260.410 12.815 260.640 15.170 ;
        RECT 261.590 12.815 261.820 15.170 ;
        RECT 263.420 12.815 263.650 15.170 ;
        RECT 264.600 12.815 264.830 15.170 ;
        RECT 265.780 12.815 266.010 15.170 ;
        RECT 266.960 12.815 267.190 15.170 ;
        RECT 268.140 12.815 268.370 15.170 ;
        RECT 269.320 12.815 269.550 15.170 ;
        RECT 270.500 12.815 270.730 15.170 ;
        RECT 271.680 12.815 271.910 15.170 ;
        RECT 214.300 12.275 214.530 12.775 ;
        RECT 215.280 12.275 215.510 12.775 ;
        RECT 216.260 12.275 216.490 12.775 ;
        RECT 217.355 12.025 217.585 12.525 ;
        RECT 217.845 12.120 218.075 12.525 ;
        RECT 217.825 11.530 218.130 12.120 ;
        RECT 218.335 12.025 218.565 12.525 ;
        RECT 218.825 12.130 219.055 12.525 ;
        RECT 218.780 11.530 219.085 12.130 ;
        RECT 219.315 12.025 219.545 12.525 ;
        RECT 219.805 12.120 220.035 12.525 ;
        RECT 219.760 11.530 220.065 12.120 ;
        RECT 220.295 12.025 220.525 12.525 ;
        RECT 220.785 12.300 221.015 12.525 ;
        RECT 220.785 11.530 221.025 12.300 ;
        RECT 223.015 12.275 223.245 12.775 ;
        RECT 223.995 12.275 224.225 12.775 ;
        RECT 224.975 12.275 225.205 12.775 ;
        RECT 255.015 12.445 257.100 12.815 ;
        RECT 257.405 12.445 262.455 12.815 ;
        RECT 262.760 12.445 272.485 12.815 ;
        RECT 213.370 11.290 221.025 11.530 ;
        RECT 212.540 10.745 213.225 11.045 ;
        RECT 213.370 8.865 213.575 11.290 ;
        RECT 221.430 11.190 222.090 11.490 ;
        RECT 225.475 11.210 225.775 11.340 ;
        RECT 213.815 9.235 214.045 9.735 ;
        RECT 214.305 9.235 214.535 9.735 ;
        RECT 214.795 9.235 215.025 9.735 ;
        RECT 215.285 9.235 215.515 9.735 ;
        RECT 215.775 9.235 216.005 9.735 ;
        RECT 216.265 9.235 216.495 9.735 ;
        RECT 216.755 9.235 216.985 9.735 ;
        RECT 217.245 9.235 217.475 9.735 ;
        RECT 218.340 8.985 218.570 9.485 ;
        RECT 219.320 8.985 219.550 9.485 ;
        RECT 220.300 8.985 220.530 9.485 ;
        RECT 203.115 8.635 203.960 8.670 ;
        RECT 203.115 8.350 208.105 8.635 ;
        RECT 211.685 8.460 212.400 8.760 ;
        RECT 213.365 8.565 214.050 8.865 ;
        RECT 221.610 8.855 221.910 11.190 ;
        RECT 225.475 10.890 227.245 11.210 ;
        RECT 252.550 11.075 253.745 12.335 ;
        RECT 225.475 10.655 225.775 10.890 ;
        RECT 226.925 10.605 227.245 10.890 ;
        RECT 226.755 9.675 227.485 10.605 ;
        RECT 222.525 8.985 222.755 9.485 ;
        RECT 223.505 8.985 223.735 9.485 ;
        RECT 224.485 8.985 224.715 9.485 ;
        RECT 226.925 9.245 227.245 9.675 ;
        RECT 228.355 9.435 228.585 9.935 ;
        RECT 229.335 9.435 229.565 9.935 ;
        RECT 230.315 9.435 230.545 9.935 ;
        RECT 233.185 9.585 234.805 9.985 ;
        RECT 239.480 9.585 241.080 9.960 ;
        RECT 252.710 9.585 253.605 11.075 ;
        RECT 233.185 9.420 241.080 9.585 ;
        RECT 226.925 8.875 227.525 9.245 ;
        RECT 216.615 8.635 217.460 8.670 ;
        RECT 213.370 8.560 213.575 8.565 ;
        RECT 212.100 8.430 212.400 8.460 ;
        RECT 203.115 8.300 203.960 8.350 ;
        RECT 200.315 7.160 200.545 7.660 ;
        RECT 200.805 7.160 201.035 7.660 ;
        RECT 201.295 7.160 201.525 7.660 ;
        RECT 201.785 7.160 202.015 7.660 ;
        RECT 202.275 7.160 202.505 7.660 ;
        RECT 202.765 7.160 202.995 7.660 ;
        RECT 203.255 7.160 203.485 7.660 ;
        RECT 203.745 7.160 203.975 7.660 ;
        RECT 204.840 7.085 205.070 8.085 ;
        RECT 205.820 7.085 206.050 8.085 ;
        RECT 206.800 7.085 207.030 8.085 ;
        RECT 207.820 7.175 208.105 8.350 ;
        RECT 216.615 8.350 221.605 8.635 ;
        RECT 216.615 8.300 217.460 8.350 ;
        RECT 209.025 7.085 209.255 8.085 ;
        RECT 210.005 7.085 210.235 8.085 ;
        RECT 210.985 7.085 211.215 8.085 ;
        RECT 213.815 7.160 214.045 7.660 ;
        RECT 214.305 7.160 214.535 7.660 ;
        RECT 214.795 7.160 215.025 7.660 ;
        RECT 215.285 7.160 215.515 7.660 ;
        RECT 215.775 7.160 216.005 7.660 ;
        RECT 216.265 7.160 216.495 7.660 ;
        RECT 216.755 7.160 216.985 7.660 ;
        RECT 217.245 7.160 217.475 7.660 ;
        RECT 218.340 7.085 218.570 8.085 ;
        RECT 219.320 7.085 219.550 8.085 ;
        RECT 220.300 7.085 220.530 8.085 ;
        RECT 221.320 7.175 221.605 8.350 ;
        RECT 222.525 7.085 222.755 8.085 ;
        RECT 223.505 7.085 223.735 8.085 ;
        RECT 224.485 7.085 224.715 8.085 ;
        RECT 170.575 7.000 171.350 7.075 ;
        RECT 170.180 6.990 171.350 7.000 ;
        RECT 164.355 6.805 171.350 6.990 ;
        RECT 131.390 4.180 132.350 5.470 ;
        RECT 135.660 4.930 137.250 5.030 ;
        RECT 138.275 4.930 138.635 5.175 ;
        RECT 135.660 4.605 138.635 4.930 ;
        RECT 140.450 4.695 140.680 5.695 ;
        RECT 135.660 4.530 137.250 4.605 ;
        RECT 138.275 4.330 138.635 4.605 ;
        RECT 131.205 1.440 132.165 2.730 ;
        RECT 140.450 2.445 140.680 3.445 ;
        RECT 141.240 1.850 141.470 5.695 ;
        RECT 142.030 4.695 142.260 6.480 ;
        RECT 142.030 2.445 142.260 3.445 ;
        RECT 142.820 1.850 143.050 5.695 ;
        RECT 143.610 4.695 143.840 5.695 ;
        RECT 144.200 4.695 144.430 6.480 ;
        RECT 145.620 6.130 147.230 6.480 ;
        RECT 164.355 6.445 170.355 6.805 ;
        RECT 170.575 6.745 171.350 6.805 ;
        RECT 226.925 6.570 227.295 8.875 ;
        RECT 233.185 8.690 246.280 9.420 ;
        RECT 256.500 9.130 256.730 12.445 ;
        RECT 258.475 11.745 258.705 12.445 ;
        RECT 263.385 11.805 263.615 12.445 ;
        RECT 257.680 11.515 259.090 11.745 ;
        RECT 257.680 9.130 257.910 11.515 ;
        RECT 258.860 9.130 259.090 11.515 ;
        RECT 260.040 11.575 263.810 11.805 ;
        RECT 260.040 9.130 260.270 11.575 ;
        RECT 261.220 9.130 261.450 11.575 ;
        RECT 262.400 9.130 262.630 11.575 ;
        RECT 263.580 9.130 263.810 11.575 ;
        RECT 228.355 7.535 228.585 8.535 ;
        RECT 229.335 7.535 229.565 8.535 ;
        RECT 230.315 7.535 230.545 8.535 ;
        RECT 233.185 8.430 234.805 8.690 ;
        RECT 239.480 8.525 246.280 8.690 ;
        RECT 239.480 8.180 241.080 8.525 ;
        RECT 231.805 6.570 232.535 6.785 ;
        RECT 143.610 2.445 143.840 3.445 ;
        RECT 144.200 2.445 144.430 3.445 ;
        RECT 144.990 1.850 145.220 5.695 ;
        RECT 146.855 3.605 147.230 6.130 ;
        RECT 159.935 4.895 161.525 4.995 ;
        RECT 162.550 4.895 162.910 5.140 ;
        RECT 159.935 4.570 162.910 4.895 ;
        RECT 164.725 4.660 164.955 5.660 ;
        RECT 159.935 4.495 161.525 4.570 ;
        RECT 162.550 4.295 162.910 4.570 ;
        RECT 152.410 2.200 152.640 4.200 ;
        RECT 153.990 2.200 154.220 4.200 ;
        RECT 155.570 2.200 155.800 4.200 ;
        RECT 157.150 2.200 157.380 4.200 ;
        RECT 164.725 2.410 164.955 3.410 ;
        RECT 140.310 1.620 145.280 1.850 ;
        RECT 165.515 1.815 165.745 5.660 ;
        RECT 166.305 4.660 166.535 6.445 ;
        RECT 166.305 2.410 166.535 3.410 ;
        RECT 167.095 1.815 167.325 5.660 ;
        RECT 167.885 4.660 168.115 5.660 ;
        RECT 168.475 4.660 168.705 6.445 ;
        RECT 169.895 6.095 171.505 6.445 ;
        RECT 226.925 6.200 232.535 6.570 ;
        RECT 167.885 2.410 168.115 3.410 ;
        RECT 168.475 2.410 168.705 3.410 ;
        RECT 169.265 1.815 169.495 5.660 ;
        RECT 171.130 3.570 171.505 6.095 ;
        RECT 176.085 2.315 176.315 4.315 ;
        RECT 177.665 2.315 177.895 4.315 ;
        RECT 179.245 2.315 179.475 4.315 ;
        RECT 180.825 2.315 181.055 4.315 ;
        RECT 184.690 2.530 184.920 4.530 ;
        RECT 186.270 2.530 186.500 4.530 ;
        RECT 187.850 2.530 188.080 4.530 ;
        RECT 189.430 2.530 189.660 4.530 ;
        RECT 111.710 -2.620 116.085 -1.765 ;
        RECT 103.505 -2.970 103.725 -2.660 ;
        RECT 94.305 -3.190 103.725 -2.970 ;
        RECT 111.710 -2.805 112.565 -2.620 ;
        RECT 104.540 -4.335 104.770 -3.835 ;
        RECT 105.520 -4.335 105.750 -3.835 ;
        RECT 106.500 -4.335 106.730 -3.835 ;
        RECT 107.770 -4.785 108.000 -3.505 ;
        RECT 108.750 -4.785 108.980 -3.505 ;
        RECT 109.730 -4.785 109.960 -3.505 ;
        RECT 110.710 -4.785 110.940 -3.505 ;
        RECT 111.710 -4.785 111.940 -2.805 ;
        RECT 131.395 -3.100 132.075 1.440 ;
        RECT 141.235 1.220 141.465 1.620 ;
        RECT 142.820 1.220 143.050 1.620 ;
        RECT 144.975 1.220 145.205 1.620 ;
        RECT 164.585 1.585 169.555 1.815 ;
        RECT 139.000 1.075 147.175 1.220 ;
        RECT 165.510 1.185 165.740 1.585 ;
        RECT 167.095 1.185 167.325 1.585 ;
        RECT 169.250 1.185 169.480 1.585 ;
        RECT 192.255 1.535 193.215 2.825 ;
        RECT 139.015 -0.105 139.245 1.075 ;
        RECT 140.595 -0.105 140.825 1.075 ;
        RECT 141.235 1.055 141.465 1.075 ;
        RECT 142.175 -0.105 142.405 1.075 ;
        RECT 143.755 -0.105 143.985 1.075 ;
        RECT 145.335 -0.105 145.565 1.075 ;
        RECT 146.915 -0.105 147.145 1.075 ;
        RECT 163.275 1.040 171.450 1.185 ;
        RECT 152.410 -1.080 152.640 0.920 ;
        RECT 153.990 -1.080 154.220 0.920 ;
        RECT 163.290 -0.140 163.520 1.040 ;
        RECT 164.870 -0.140 165.100 1.040 ;
        RECT 165.510 1.020 165.740 1.040 ;
        RECT 166.450 -0.140 166.680 1.040 ;
        RECT 168.030 -0.140 168.260 1.040 ;
        RECT 169.610 -0.140 169.840 1.040 ;
        RECT 171.190 -0.140 171.420 1.040 ;
        RECT 176.085 -0.965 176.315 1.035 ;
        RECT 177.665 -0.965 177.895 1.035 ;
        RECT 184.690 -0.750 184.920 1.250 ;
        RECT 186.270 -0.750 186.500 1.250 ;
        RECT 192.405 -3.100 193.085 1.535 ;
        RECT 131.395 -3.780 193.085 -3.100 ;
        RECT 231.135 -3.160 231.505 6.200 ;
        RECT 231.805 5.855 232.535 6.200 ;
        RECT 238.790 -3.160 239.765 -2.860 ;
        RECT 231.135 -3.530 239.765 -3.160 ;
        RECT 238.790 -3.760 239.765 -3.530 ;
        RECT 26.325 -5.495 26.545 -5.185 ;
        RECT 18.840 -5.715 26.545 -5.495 ;
        RECT 34.530 -5.330 37.060 -5.100 ;
        RECT 38.420 -5.220 40.505 -4.850 ;
        RECT 40.810 -5.220 45.860 -4.850 ;
        RECT 46.165 -5.220 55.890 -4.850 ;
        RECT 107.770 -5.015 111.940 -4.785 ;
        RECT -17.320 -6.830 -13.150 -6.600 ;
        RECT -20.550 -8.050 -20.320 -7.050 ;
        RECT -19.570 -8.050 -19.340 -7.050 ;
        RECT -18.590 -8.050 -18.360 -7.050 ;
        RECT -17.810 -8.050 -17.580 -7.050 ;
        RECT -17.320 -8.050 -17.090 -6.830 ;
        RECT -16.830 -8.050 -16.600 -7.050 ;
        RECT -16.340 -8.050 -16.110 -6.830 ;
        RECT -15.850 -8.050 -15.620 -7.050 ;
        RECT -15.360 -8.050 -15.130 -6.830 ;
        RECT -14.870 -8.050 -14.640 -7.050 ;
        RECT -14.380 -8.050 -14.150 -6.830 ;
        RECT 27.360 -6.860 27.590 -6.360 ;
        RECT 28.340 -6.860 28.570 -6.360 ;
        RECT 29.320 -6.860 29.550 -6.360 ;
        RECT -13.890 -8.050 -13.660 -7.050 ;
        RECT 30.590 -7.310 30.820 -6.030 ;
        RECT 31.570 -7.310 31.800 -6.030 ;
        RECT 32.550 -7.310 32.780 -6.030 ;
        RECT 33.530 -7.310 33.760 -6.030 ;
        RECT 34.530 -7.310 34.760 -5.330 ;
        RECT 36.670 -5.465 37.060 -5.330 ;
        RECT 36.670 -6.035 37.215 -5.465 ;
        RECT 30.590 -7.540 34.760 -7.310 ;
        RECT 27.360 -8.760 27.590 -7.760 ;
        RECT 28.340 -8.760 28.570 -7.760 ;
        RECT 29.320 -8.760 29.550 -7.760 ;
        RECT 30.590 -8.760 30.820 -7.540 ;
        RECT 31.570 -8.760 31.800 -7.540 ;
        RECT 32.550 -8.760 32.780 -7.540 ;
        RECT 33.530 -8.760 33.760 -7.540 ;
        RECT 39.905 -8.535 40.135 -5.220 ;
        RECT 41.880 -5.920 42.110 -5.220 ;
        RECT 46.790 -5.860 47.020 -5.220 ;
        RECT 41.085 -6.150 42.495 -5.920 ;
        RECT 41.085 -8.535 41.315 -6.150 ;
        RECT 42.265 -8.535 42.495 -6.150 ;
        RECT 43.445 -6.090 47.215 -5.860 ;
        RECT 43.445 -8.535 43.675 -6.090 ;
        RECT 44.625 -8.535 44.855 -6.090 ;
        RECT 45.805 -8.535 46.035 -6.090 ;
        RECT 46.985 -8.535 47.215 -6.090 ;
        RECT 104.540 -6.235 104.770 -5.235 ;
        RECT 105.520 -6.235 105.750 -5.235 ;
        RECT 106.500 -6.235 106.730 -5.235 ;
        RECT 107.770 -6.235 108.000 -5.015 ;
        RECT 108.750 -6.235 108.980 -5.015 ;
        RECT 109.730 -6.235 109.960 -5.015 ;
        RECT 110.710 -6.235 110.940 -5.015 ;
        RECT 245.385 -16.855 246.280 8.525 ;
        RECT 254.025 -1.740 254.255 0.615 ;
        RECT 255.205 -1.740 255.435 0.615 ;
        RECT 257.035 -1.740 257.265 0.615 ;
        RECT 258.215 -1.740 258.445 0.615 ;
        RECT 259.395 -1.740 259.625 0.615 ;
        RECT 260.575 -1.740 260.805 0.615 ;
        RECT 262.405 -1.740 262.635 0.615 ;
        RECT 263.585 -1.740 263.815 0.615 ;
        RECT 264.765 -1.740 264.995 0.615 ;
        RECT 265.945 -1.740 266.175 0.615 ;
        RECT 267.125 -1.740 267.355 0.615 ;
        RECT 268.305 -1.740 268.535 0.615 ;
        RECT 269.485 -1.740 269.715 0.615 ;
        RECT 270.665 -1.740 270.895 0.615 ;
        RECT 254.000 -2.110 256.085 -1.740 ;
        RECT 256.390 -2.110 261.440 -1.740 ;
        RECT 261.745 -2.110 271.470 -1.740 ;
        RECT 255.485 -5.425 255.715 -2.110 ;
        RECT 257.460 -2.810 257.690 -2.110 ;
        RECT 262.370 -2.750 262.600 -2.110 ;
        RECT 256.665 -3.040 258.075 -2.810 ;
        RECT 256.665 -5.425 256.895 -3.040 ;
        RECT 257.845 -5.425 258.075 -3.040 ;
        RECT 259.025 -2.980 262.795 -2.750 ;
        RECT 259.025 -5.425 259.255 -2.980 ;
        RECT 260.205 -5.425 260.435 -2.980 ;
        RECT 261.385 -5.425 261.615 -2.980 ;
        RECT 262.565 -5.425 262.795 -2.980 ;
        RECT 244.830 -18.485 246.385 -16.855 ;
        RECT 254.025 -16.975 254.255 -14.620 ;
        RECT 255.205 -16.975 255.435 -14.620 ;
        RECT 257.035 -16.975 257.265 -14.620 ;
        RECT 258.215 -16.975 258.445 -14.620 ;
        RECT 259.395 -16.975 259.625 -14.620 ;
        RECT 260.575 -16.975 260.805 -14.620 ;
        RECT 262.405 -16.975 262.635 -14.620 ;
        RECT 263.585 -16.975 263.815 -14.620 ;
        RECT 264.765 -16.975 264.995 -14.620 ;
        RECT 265.945 -16.975 266.175 -14.620 ;
        RECT 267.125 -16.975 267.355 -14.620 ;
        RECT 268.305 -16.975 268.535 -14.620 ;
        RECT 269.485 -16.975 269.715 -14.620 ;
        RECT 270.665 -16.975 270.895 -14.620 ;
        RECT 271.905 -16.975 272.135 -14.620 ;
        RECT 273.085 -16.975 273.315 -14.620 ;
        RECT 274.265 -16.975 274.495 -14.620 ;
        RECT 275.445 -16.975 275.675 -14.620 ;
        RECT 276.625 -16.975 276.855 -14.620 ;
        RECT 277.805 -16.975 278.035 -14.620 ;
        RECT 278.985 -16.975 279.215 -14.620 ;
        RECT 280.165 -16.975 280.395 -14.620 ;
        RECT 281.345 -16.975 281.575 -14.620 ;
        RECT 282.525 -16.975 282.755 -14.620 ;
        RECT 283.705 -16.975 283.935 -14.620 ;
        RECT 284.885 -16.975 285.115 -14.620 ;
        RECT 286.065 -16.975 286.295 -14.620 ;
        RECT 287.245 -16.975 287.475 -14.620 ;
        RECT 288.425 -16.975 288.655 -14.620 ;
        RECT 289.605 -16.975 289.835 -14.620 ;
        RECT 290.785 -16.975 291.015 -14.620 ;
        RECT 312.425 -15.190 312.655 -14.190 ;
        RECT 313.405 -15.190 313.635 -14.190 ;
        RECT 314.385 -15.190 314.615 -14.190 ;
        RECT 316.675 -15.190 316.905 -14.190 ;
        RECT 317.655 -15.190 317.885 -14.190 ;
        RECT 318.635 -15.190 318.865 -14.190 ;
        RECT 319.415 -15.190 319.645 -14.190 ;
        RECT 319.905 -15.410 320.135 -14.190 ;
        RECT 320.395 -15.190 320.625 -14.190 ;
        RECT 320.885 -15.410 321.115 -14.190 ;
        RECT 321.375 -15.190 321.605 -14.190 ;
        RECT 321.865 -15.410 322.095 -14.190 ;
        RECT 322.355 -15.190 322.585 -14.190 ;
        RECT 322.845 -15.410 323.075 -14.190 ;
        RECT 323.335 -15.190 323.565 -14.190 ;
        RECT 319.905 -15.640 324.075 -15.410 ;
        RECT 312.425 -16.590 312.655 -16.090 ;
        RECT 313.405 -16.590 313.635 -16.090 ;
        RECT 314.385 -16.590 314.615 -16.090 ;
        RECT 315.200 -16.270 315.860 -16.050 ;
        RECT 315.640 -16.770 315.860 -16.270 ;
        RECT 316.675 -16.590 316.905 -16.090 ;
        RECT 317.655 -16.590 317.885 -16.090 ;
        RECT 318.635 -16.590 318.865 -16.090 ;
        RECT 319.415 -16.770 319.645 -15.920 ;
        RECT 254.000 -17.345 256.085 -16.975 ;
        RECT 256.390 -17.345 261.440 -16.975 ;
        RECT 261.745 -17.345 271.470 -16.975 ;
        RECT 271.775 -17.345 291.160 -16.975 ;
        RECT 315.640 -16.990 319.650 -16.770 ;
        RECT 319.905 -16.920 320.135 -15.640 ;
        RECT 320.395 -16.920 320.625 -15.920 ;
        RECT 320.885 -16.920 321.115 -15.640 ;
        RECT 321.375 -16.920 321.605 -15.920 ;
        RECT 321.865 -16.920 322.095 -15.640 ;
        RECT 322.355 -16.920 322.585 -15.920 ;
        RECT 322.845 -16.920 323.075 -15.640 ;
        RECT 323.335 -16.920 323.565 -15.920 ;
        RECT 323.845 -16.905 324.075 -15.640 ;
        RECT 325.935 -16.905 326.650 -16.685 ;
        RECT 309.365 -17.300 310.335 -17.035 ;
        RECT 315.640 -17.300 315.860 -16.990 ;
        RECT 255.485 -20.660 255.715 -17.345 ;
        RECT 257.460 -18.045 257.690 -17.345 ;
        RECT 262.370 -17.985 262.600 -17.345 ;
        RECT 272.005 -17.925 272.235 -17.345 ;
        RECT 309.365 -17.520 315.860 -17.300 ;
        RECT 323.845 -17.135 326.650 -16.905 ;
        RECT 309.365 -17.580 310.335 -17.520 ;
        RECT 256.665 -18.275 258.075 -18.045 ;
        RECT 256.665 -20.660 256.895 -18.275 ;
        RECT 257.845 -20.660 258.075 -18.275 ;
        RECT 259.025 -18.215 262.795 -17.985 ;
        RECT 259.025 -20.660 259.255 -18.215 ;
        RECT 260.205 -20.660 260.435 -18.215 ;
        RECT 261.385 -20.660 261.615 -18.215 ;
        RECT 262.565 -20.660 262.795 -18.215 ;
        RECT 263.745 -18.155 272.235 -17.925 ;
        RECT 263.745 -20.660 263.975 -18.155 ;
        RECT 264.925 -20.660 265.155 -18.155 ;
        RECT 266.105 -20.660 266.335 -18.155 ;
        RECT 267.285 -20.660 267.515 -18.155 ;
        RECT 268.465 -20.660 268.695 -18.155 ;
        RECT 269.645 -20.660 269.875 -18.155 ;
        RECT 270.825 -20.660 271.055 -18.155 ;
        RECT 272.005 -20.660 272.235 -18.155 ;
        RECT 316.675 -18.665 316.905 -18.165 ;
        RECT 317.655 -18.665 317.885 -18.165 ;
        RECT 318.635 -18.665 318.865 -18.165 ;
        RECT 319.905 -19.115 320.135 -17.835 ;
        RECT 320.885 -19.115 321.115 -17.835 ;
        RECT 321.865 -19.115 322.095 -17.835 ;
        RECT 322.845 -19.115 323.075 -17.835 ;
        RECT 323.845 -19.115 324.075 -17.135 ;
        RECT 325.935 -17.340 326.650 -17.135 ;
        RECT 438.925 -17.905 441.050 -15.945 ;
        RECT 319.905 -19.345 324.075 -19.115 ;
        RECT 316.675 -20.565 316.905 -19.565 ;
        RECT 317.655 -20.565 317.885 -19.565 ;
        RECT 318.635 -20.565 318.865 -19.565 ;
        RECT 319.905 -20.565 320.135 -19.345 ;
        RECT 320.885 -20.565 321.115 -19.345 ;
        RECT 321.865 -20.565 322.095 -19.345 ;
        RECT 322.845 -20.565 323.075 -19.345 ;
        RECT -64.370 -76.190 -39.350 -74.845 ;
        RECT -64.325 -76.200 -59.620 -76.190 ;
        RECT -74.785 -78.640 -74.555 -76.640 ;
        RECT -74.195 -78.640 -73.965 -76.640 ;
        RECT -73.605 -78.640 -73.375 -76.640 ;
        RECT -73.015 -78.640 -72.785 -76.640 ;
        RECT -72.425 -78.640 -72.195 -76.640 ;
        RECT -71.835 -78.640 -71.605 -76.640 ;
        RECT -71.245 -78.640 -71.015 -76.640 ;
        RECT -70.655 -78.640 -70.425 -76.640 ;
        RECT -70.065 -78.640 -69.835 -76.640 ;
        RECT -69.475 -78.640 -69.245 -76.640 ;
        RECT -68.885 -78.640 -68.655 -76.640 ;
        RECT -68.295 -78.640 -68.065 -76.640 ;
        RECT -67.705 -78.640 -67.475 -76.640 ;
        RECT -67.115 -78.640 -66.885 -76.640 ;
        RECT -66.525 -78.640 -66.295 -76.640 ;
        RECT -65.935 -78.640 -65.705 -76.640 ;
        RECT -65.345 -78.640 -65.115 -76.640 ;
        RECT -64.755 -78.640 -64.525 -76.640 ;
        RECT -64.165 -78.640 -63.935 -76.640 ;
        RECT -63.575 -78.640 -63.345 -76.640 ;
        RECT -62.985 -78.640 -62.755 -76.640 ;
        RECT -62.395 -78.640 -62.165 -76.640 ;
        RECT -61.805 -78.640 -61.575 -76.640 ;
        RECT -61.215 -78.640 -60.985 -76.640 ;
        RECT -60.625 -78.640 -60.395 -76.640 ;
        RECT -60.035 -78.640 -59.805 -76.640 ;
        RECT -59.445 -78.640 -59.215 -76.640 ;
        RECT -58.855 -78.640 -58.625 -76.640 ;
        RECT -58.265 -78.640 -58.035 -76.640 ;
        RECT -57.675 -78.640 -57.445 -76.640 ;
        RECT -57.085 -78.640 -56.855 -76.640 ;
        RECT -55.905 -78.640 -55.675 -76.640 ;
        RECT -54.725 -78.640 -54.495 -76.640 ;
        RECT -53.545 -78.640 -53.315 -76.640 ;
        RECT -52.365 -78.640 -52.135 -76.640 ;
        RECT -51.185 -78.640 -50.955 -76.640 ;
        RECT -50.005 -78.640 -49.775 -76.640 ;
        RECT -48.825 -78.640 -48.595 -76.640 ;
        RECT -47.645 -78.640 -47.415 -76.640 ;
        RECT -47.055 -79.085 -46.825 -76.640 ;
        RECT -46.465 -78.640 -46.235 -76.640 ;
        RECT -45.875 -79.085 -45.645 -76.640 ;
        RECT -45.285 -78.640 -45.055 -76.640 ;
        RECT -44.695 -79.085 -44.465 -76.640 ;
        RECT -44.105 -78.640 -43.875 -76.640 ;
        RECT -43.515 -79.085 -43.285 -76.640 ;
        RECT -42.925 -78.640 -42.695 -76.640 ;
        RECT -47.055 -79.315 -43.285 -79.085 ;
        RECT -42.335 -79.025 -42.105 -76.640 ;
        RECT -41.745 -78.640 -41.515 -76.640 ;
        RECT -41.155 -79.025 -40.925 -76.640 ;
        RECT -40.565 -78.640 -40.335 -76.640 ;
        RECT -42.335 -79.255 -40.925 -79.025 ;
        RECT -46.860 -79.955 -46.630 -79.315 ;
        RECT -41.950 -79.955 -41.720 -79.255 ;
        RECT -39.975 -79.955 -39.745 -76.640 ;
        RECT -39.385 -78.640 -39.155 -76.640 ;
        RECT 60.375 -77.225 438.480 -75.805 ;
        RECT -55.730 -80.325 -46.005 -79.955 ;
        RECT -45.700 -80.325 -40.650 -79.955 ;
        RECT -40.345 -80.325 -38.260 -79.955 ;
        RECT -55.155 -82.680 -54.925 -80.325 ;
        RECT -53.975 -82.680 -53.745 -80.325 ;
        RECT -52.795 -82.680 -52.565 -80.325 ;
        RECT -51.615 -82.680 -51.385 -80.325 ;
        RECT -50.435 -82.680 -50.205 -80.325 ;
        RECT -49.255 -82.680 -49.025 -80.325 ;
        RECT -48.075 -82.680 -47.845 -80.325 ;
        RECT -46.895 -82.680 -46.665 -80.325 ;
        RECT -45.065 -82.680 -44.835 -80.325 ;
        RECT -43.885 -82.680 -43.655 -80.325 ;
        RECT -42.705 -82.680 -42.475 -80.325 ;
        RECT -41.525 -82.680 -41.295 -80.325 ;
        RECT -39.695 -82.680 -39.465 -80.325 ;
        RECT -38.515 -82.680 -38.285 -80.325 ;
        RECT -83.020 -90.675 39.020 -89.725 ;
        RECT -113.230 -96.920 -113.000 -95.920 ;
        RECT -112.250 -96.920 -112.020 -95.920 ;
        RECT -111.270 -96.920 -111.040 -95.920 ;
        RECT -107.580 -96.920 -107.350 -95.920 ;
        RECT -83.020 -96.120 -82.070 -90.675 ;
        RECT -75.235 -92.985 -75.005 -91.985 ;
        RECT -74.255 -92.985 -74.025 -91.985 ;
        RECT -73.275 -92.985 -73.045 -91.985 ;
        RECT -72.125 -93.250 -71.840 -92.075 ;
        RECT -71.050 -92.985 -70.820 -91.985 ;
        RECT -70.070 -92.985 -69.840 -91.985 ;
        RECT -69.090 -92.985 -68.860 -91.985 ;
        RECT -67.995 -92.560 -67.765 -92.060 ;
        RECT -67.505 -92.560 -67.275 -92.060 ;
        RECT -67.015 -92.560 -66.785 -92.060 ;
        RECT -66.525 -92.560 -66.295 -92.060 ;
        RECT -66.035 -92.560 -65.805 -92.060 ;
        RECT -65.545 -92.560 -65.315 -92.060 ;
        RECT -65.055 -92.560 -64.825 -92.060 ;
        RECT -64.565 -92.560 -64.335 -92.060 ;
        RECT -61.735 -92.985 -61.505 -91.985 ;
        RECT -60.755 -92.985 -60.525 -91.985 ;
        RECT -59.775 -92.985 -59.545 -91.985 ;
        RECT -67.980 -93.250 -67.135 -93.200 ;
        RECT -72.125 -93.535 -67.135 -93.250 ;
        RECT -58.625 -93.250 -58.340 -92.075 ;
        RECT -57.550 -92.985 -57.320 -91.985 ;
        RECT -56.570 -92.985 -56.340 -91.985 ;
        RECT -55.590 -92.985 -55.360 -91.985 ;
        RECT -54.495 -92.560 -54.265 -92.060 ;
        RECT -54.005 -92.560 -53.775 -92.060 ;
        RECT -53.515 -92.560 -53.285 -92.060 ;
        RECT -53.025 -92.560 -52.795 -92.060 ;
        RECT -52.535 -92.560 -52.305 -92.060 ;
        RECT -52.045 -92.560 -51.815 -92.060 ;
        RECT -51.555 -92.560 -51.325 -92.060 ;
        RECT -51.065 -92.560 -50.835 -92.060 ;
        RECT -54.480 -93.250 -53.635 -93.200 ;
        RECT -62.920 -93.360 -62.620 -93.330 ;
        RECT -64.095 -93.465 -63.890 -93.460 ;
        RECT -67.980 -93.570 -67.135 -93.535 ;
        RECT -75.725 -94.385 -75.495 -93.885 ;
        RECT -75.235 -94.385 -75.005 -93.885 ;
        RECT -74.745 -94.385 -74.515 -93.885 ;
        RECT -74.255 -94.385 -74.025 -93.885 ;
        RECT -73.765 -94.385 -73.535 -93.885 ;
        RECT -73.275 -94.385 -73.045 -93.885 ;
        RECT -74.555 -95.500 -73.870 -95.200 ;
        RECT -76.295 -95.790 -75.995 -95.555 ;
        RECT -77.605 -96.110 -75.995 -95.790 ;
        RECT -103.235 -98.030 -103.005 -96.530 ;
        RECT -113.720 -100.455 -113.490 -98.955 ;
        RECT -113.230 -100.455 -113.000 -98.955 ;
        RECT -112.740 -100.455 -112.510 -98.955 ;
        RECT -112.170 -100.460 -111.940 -98.960 ;
        RECT -111.680 -100.460 -111.450 -98.960 ;
        RECT -111.190 -100.460 -110.960 -98.960 ;
        RECT -110.625 -100.460 -110.395 -98.960 ;
        RECT -110.135 -100.460 -109.905 -98.960 ;
        RECT -109.645 -100.460 -109.415 -98.960 ;
        RECT -108.070 -100.460 -107.840 -99.460 ;
        RECT -107.580 -100.040 -107.350 -99.460 ;
        RECT -107.580 -100.215 -105.785 -100.040 ;
        RECT -107.580 -100.460 -107.350 -100.215 ;
        RECT -120.160 -103.055 -119.655 -102.780 ;
        RECT -120.920 -103.995 -119.655 -103.055 ;
        RECT -120.920 -104.210 -119.720 -103.995 ;
        RECT -128.320 -117.020 -125.195 -113.895 ;
        RECT -120.920 -148.835 -120.240 -104.210 ;
        RECT -112.945 -107.575 -112.715 -106.075 ;
        RECT -113.435 -110.255 -113.205 -108.760 ;
        RECT -113.440 -110.440 -113.205 -110.255 ;
        RECT -112.945 -110.260 -112.715 -108.760 ;
        RECT -112.455 -110.440 -112.225 -108.760 ;
        RECT -111.965 -110.260 -111.735 -106.075 ;
        RECT -109.900 -106.850 -109.670 -106.070 ;
        RECT -108.920 -106.840 -108.690 -106.070 ;
        RECT -109.410 -106.850 -108.200 -106.840 ;
        RECT -107.940 -106.850 -107.710 -106.070 ;
        RECT -109.900 -107.080 -106.715 -106.850 ;
        RECT -109.900 -107.725 -109.670 -107.225 ;
        RECT -109.410 -107.725 -109.180 -107.080 ;
        RECT -108.920 -107.725 -108.690 -107.225 ;
        RECT -108.430 -107.725 -108.200 -107.080 ;
        RECT -105.960 -107.885 -105.785 -100.215 ;
        RECT -103.725 -100.710 -103.495 -99.215 ;
        RECT -103.730 -100.895 -103.495 -100.710 ;
        RECT -103.235 -100.715 -103.005 -99.215 ;
        RECT -102.745 -100.895 -102.515 -99.215 ;
        RECT -102.255 -100.715 -102.025 -96.530 ;
        RECT -100.190 -97.305 -99.960 -96.525 ;
        RECT -99.210 -97.295 -98.980 -96.525 ;
        RECT -99.700 -97.305 -98.490 -97.295 ;
        RECT -98.230 -97.305 -98.000 -96.525 ;
        RECT -84.925 -96.685 -81.540 -96.120 ;
        RECT -100.190 -97.535 -97.005 -97.305 ;
        RECT -100.190 -98.180 -99.960 -97.680 ;
        RECT -99.700 -98.180 -99.470 -97.535 ;
        RECT -99.210 -98.180 -98.980 -97.680 ;
        RECT -98.720 -98.180 -98.490 -97.535 ;
        RECT -96.590 -97.660 -95.860 -97.370 ;
        RECT -96.590 -97.790 -96.185 -97.660 ;
        RECT -98.150 -97.965 -96.185 -97.790 ;
        RECT -101.765 -100.895 -101.535 -99.215 ;
        RECT -103.730 -101.130 -101.535 -100.895 ;
        RECT -98.150 -103.315 -97.975 -97.965 ;
        RECT -95.550 -98.475 -93.355 -98.240 ;
        RECT -95.550 -98.660 -95.315 -98.475 ;
        RECT -95.545 -100.155 -95.315 -98.660 ;
        RECT -95.055 -100.155 -94.825 -98.655 ;
        RECT -94.565 -100.155 -94.335 -98.475 ;
        RECT -96.820 -100.635 -95.835 -100.365 ;
        RECT -105.630 -103.490 -97.975 -103.315 ;
        RECT -105.630 -107.230 -105.455 -103.490 ;
        RECT -104.080 -106.600 -103.850 -105.600 ;
        RECT -103.100 -106.600 -102.870 -105.600 ;
        RECT -102.120 -106.600 -101.890 -105.600 ;
        RECT -98.430 -106.600 -98.200 -105.600 ;
        RECT -105.630 -107.460 -105.210 -107.230 ;
        RECT -111.475 -110.440 -111.245 -108.760 ;
        RECT -107.055 -109.055 -106.765 -108.370 ;
        RECT -105.985 -108.570 -105.695 -107.885 ;
        RECT -105.500 -107.915 -105.210 -107.460 ;
        RECT -96.105 -107.655 -95.835 -100.635 ;
        RECT -95.055 -102.840 -94.825 -101.340 ;
        RECT -94.075 -102.840 -93.845 -98.655 ;
        RECT -93.585 -100.155 -93.355 -98.475 ;
        RECT -87.820 -98.725 -87.590 -97.225 ;
        RECT -87.330 -98.725 -87.100 -97.225 ;
        RECT -86.840 -98.725 -86.610 -97.225 ;
        RECT -85.630 -98.725 -85.400 -97.225 ;
        RECT -85.140 -98.725 -84.910 -97.225 ;
        RECT -88.315 -99.215 -83.215 -98.890 ;
        RECT -83.540 -99.630 -83.215 -99.215 ;
        RECT -83.570 -99.990 -83.045 -99.630 ;
        RECT -92.010 -101.690 -91.780 -101.190 ;
        RECT -91.520 -101.835 -91.290 -101.190 ;
        RECT -91.030 -101.690 -90.800 -101.190 ;
        RECT -90.540 -101.835 -90.310 -101.190 ;
        RECT -92.010 -102.065 -88.825 -101.835 ;
        RECT -92.010 -102.845 -91.780 -102.065 ;
        RECT -91.520 -102.075 -90.310 -102.065 ;
        RECT -91.030 -102.845 -90.800 -102.075 ;
        RECT -90.050 -102.845 -89.820 -102.065 ;
        RECT -87.820 -103.285 -87.590 -100.285 ;
        RECT -86.765 -103.285 -86.535 -100.285 ;
        RECT -86.275 -103.285 -86.045 -100.285 ;
        RECT -85.785 -103.285 -85.555 -100.285 ;
        RECT -84.725 -103.285 -84.495 -100.285 ;
        RECT -96.355 -108.405 -95.705 -107.655 ;
        RECT -94.925 -107.765 -94.695 -106.485 ;
        RECT -93.945 -107.755 -93.715 -106.485 ;
        RECT -94.435 -107.765 -93.225 -107.755 ;
        RECT -92.965 -107.765 -92.735 -106.485 ;
        RECT -90.060 -107.340 -89.830 -105.840 ;
        RECT -94.925 -107.995 -91.740 -107.765 ;
        RECT -91.030 -107.860 -90.235 -107.570 ;
        RECT -104.570 -110.135 -104.340 -108.635 ;
        RECT -104.080 -110.135 -103.850 -108.635 ;
        RECT -103.590 -110.135 -103.360 -108.635 ;
        RECT -103.020 -110.140 -102.790 -108.640 ;
        RECT -102.530 -110.140 -102.300 -108.640 ;
        RECT -102.040 -110.140 -101.810 -108.640 ;
        RECT -101.475 -110.140 -101.245 -108.640 ;
        RECT -100.985 -110.140 -100.755 -108.640 ;
        RECT -100.495 -110.140 -100.265 -108.640 ;
        RECT -94.925 -109.135 -94.695 -108.135 ;
        RECT -94.435 -109.135 -94.205 -107.995 ;
        RECT -93.945 -109.135 -93.715 -108.135 ;
        RECT -93.455 -109.135 -93.225 -107.995 ;
        RECT -90.900 -108.135 -90.630 -107.860 ;
        RECT -92.270 -108.405 -90.630 -108.135 ;
        RECT -98.920 -110.140 -98.690 -109.140 ;
        RECT -98.430 -110.140 -98.200 -109.140 ;
        RECT -92.270 -109.855 -92.000 -108.405 ;
        RECT -97.485 -110.125 -92.000 -109.855 ;
        RECT -90.550 -110.020 -90.320 -108.525 ;
        RECT -113.440 -110.675 -111.245 -110.440 ;
        RECT -97.425 -113.695 -96.225 -110.125 ;
        RECT -90.555 -110.205 -90.320 -110.020 ;
        RECT -90.060 -110.025 -89.830 -108.525 ;
        RECT -89.570 -110.205 -89.340 -108.525 ;
        RECT -89.080 -110.025 -88.850 -105.840 ;
        RECT -87.015 -106.615 -86.785 -105.835 ;
        RECT -86.035 -106.605 -85.805 -105.835 ;
        RECT -86.525 -106.615 -85.315 -106.605 ;
        RECT -85.055 -106.615 -84.825 -105.835 ;
        RECT -87.015 -106.845 -83.830 -106.615 ;
        RECT -87.015 -107.490 -86.785 -106.990 ;
        RECT -86.525 -107.490 -86.295 -106.845 ;
        RECT -86.035 -107.490 -85.805 -106.990 ;
        RECT -85.545 -107.490 -85.315 -106.845 ;
        RECT -82.105 -107.665 -81.540 -96.685 ;
        RECT -77.605 -105.690 -77.285 -96.110 ;
        RECT -76.295 -96.240 -75.995 -96.110 ;
        RECT -74.480 -96.590 -74.005 -95.500 ;
        RECT -72.430 -96.090 -72.130 -93.755 ;
        RECT -64.570 -93.765 -63.885 -93.465 ;
        RECT -62.920 -93.660 -62.205 -93.360 ;
        RECT -58.625 -93.535 -53.635 -93.250 ;
        RECT -54.480 -93.570 -53.635 -93.535 ;
        RECT -71.540 -94.385 -71.310 -93.885 ;
        RECT -71.050 -94.385 -70.820 -93.885 ;
        RECT -70.560 -94.385 -70.330 -93.885 ;
        RECT -70.070 -94.385 -69.840 -93.885 ;
        RECT -69.580 -94.385 -69.350 -93.885 ;
        RECT -69.090 -94.385 -68.860 -93.885 ;
        RECT -67.995 -94.635 -67.765 -94.135 ;
        RECT -67.505 -94.635 -67.275 -94.135 ;
        RECT -67.015 -94.635 -66.785 -94.135 ;
        RECT -66.525 -94.635 -66.295 -94.135 ;
        RECT -66.035 -94.635 -65.805 -94.135 ;
        RECT -65.545 -94.635 -65.315 -94.135 ;
        RECT -65.055 -94.635 -64.825 -94.135 ;
        RECT -64.565 -94.635 -64.335 -94.135 ;
        RECT -72.610 -96.390 -71.950 -96.090 ;
        RECT -64.095 -96.190 -63.890 -93.765 ;
        RECT -63.745 -95.945 -63.060 -95.645 ;
        RECT -71.545 -96.430 -63.890 -96.190 ;
        RECT -74.600 -96.890 -73.940 -96.590 ;
        RECT -75.725 -97.675 -75.495 -97.175 ;
        RECT -75.235 -97.675 -75.005 -97.175 ;
        RECT -74.745 -97.675 -74.515 -97.175 ;
        RECT -74.255 -97.675 -74.025 -97.175 ;
        RECT -73.765 -97.675 -73.535 -97.175 ;
        RECT -73.275 -97.675 -73.045 -97.175 ;
        RECT -71.545 -97.200 -71.305 -96.430 ;
        RECT -71.535 -97.425 -71.305 -97.200 ;
        RECT -71.045 -97.425 -70.815 -96.925 ;
        RECT -70.585 -97.020 -70.280 -96.430 ;
        RECT -70.555 -97.425 -70.325 -97.020 ;
        RECT -70.065 -97.425 -69.835 -96.925 ;
        RECT -69.605 -97.030 -69.300 -96.430 ;
        RECT -69.575 -97.425 -69.345 -97.030 ;
        RECT -69.085 -97.425 -68.855 -96.925 ;
        RECT -68.650 -97.020 -68.345 -96.430 ;
        RECT -68.595 -97.425 -68.365 -97.020 ;
        RECT -68.105 -97.425 -67.875 -96.925 ;
        RECT -67.010 -97.675 -66.780 -97.175 ;
        RECT -66.520 -97.675 -66.290 -97.175 ;
        RECT -66.030 -97.675 -65.800 -97.175 ;
        RECT -65.540 -97.675 -65.310 -97.175 ;
        RECT -65.050 -97.675 -64.820 -97.175 ;
        RECT -64.560 -97.675 -64.330 -97.175 ;
        RECT -68.735 -98.025 -67.890 -97.990 ;
        RECT -68.735 -98.310 -63.745 -98.025 ;
        RECT -63.500 -98.185 -63.200 -95.945 ;
        RECT -62.920 -97.400 -62.620 -93.660 ;
        RECT -51.125 -93.775 -50.355 -93.475 ;
        RECT -62.225 -94.385 -61.995 -93.885 ;
        RECT -61.735 -94.385 -61.505 -93.885 ;
        RECT -61.245 -94.385 -61.015 -93.885 ;
        RECT -60.755 -94.385 -60.525 -93.885 ;
        RECT -60.265 -94.385 -60.035 -93.885 ;
        RECT -59.775 -94.385 -59.545 -93.885 ;
        RECT -61.570 -95.530 -60.885 -95.230 ;
        RECT -61.515 -96.570 -61.040 -95.530 ;
        RECT -58.870 -95.650 -58.570 -93.830 ;
        RECT -58.040 -94.385 -57.810 -93.885 ;
        RECT -57.550 -94.385 -57.320 -93.885 ;
        RECT -57.060 -94.385 -56.830 -93.885 ;
        RECT -56.570 -94.385 -56.340 -93.885 ;
        RECT -56.080 -94.385 -55.850 -93.885 ;
        RECT -55.590 -94.385 -55.360 -93.885 ;
        RECT -54.495 -94.635 -54.265 -94.135 ;
        RECT -54.005 -94.635 -53.775 -94.135 ;
        RECT -53.515 -94.635 -53.285 -94.135 ;
        RECT -53.025 -94.635 -52.795 -94.135 ;
        RECT -52.535 -94.635 -52.305 -94.135 ;
        RECT -52.045 -94.635 -51.815 -94.135 ;
        RECT -51.555 -94.635 -51.325 -94.135 ;
        RECT -51.065 -94.635 -50.835 -94.135 ;
        RECT -50.585 -95.150 -50.355 -93.775 ;
        RECT -54.450 -95.375 -50.355 -95.150 ;
        RECT -54.450 -95.380 -50.395 -95.375 ;
        RECT -59.015 -95.950 -58.355 -95.650 ;
        RECT -54.450 -96.210 -54.220 -95.380 ;
        RECT -48.380 -95.530 -47.720 -95.230 ;
        RECT -48.295 -95.855 -47.820 -95.530 ;
        RECT -45.620 -95.855 -45.145 -90.675 ;
        RECT -44.405 -95.035 -44.175 -92.035 ;
        RECT -43.345 -95.035 -43.115 -92.035 ;
        RECT -42.855 -95.035 -42.625 -92.035 ;
        RECT -42.365 -95.035 -42.135 -92.035 ;
        RECT -41.310 -95.035 -41.080 -92.035 ;
        RECT -37.255 -94.015 -37.025 -93.015 ;
        RECT -36.765 -94.015 -36.535 -93.015 ;
        RECT -36.275 -94.015 -36.045 -93.015 ;
        RECT -35.675 -94.015 -35.445 -93.015 ;
        RECT -35.185 -94.015 -34.955 -93.015 ;
        RECT -34.695 -94.015 -34.465 -93.015 ;
        RECT -32.885 -94.015 -32.655 -93.015 ;
        RECT -31.905 -94.015 -31.675 -93.015 ;
        RECT -30.355 -94.015 -30.125 -93.015 ;
        RECT -28.810 -94.015 -28.580 -93.015 ;
        RECT -24.755 -94.015 -24.525 -93.015 ;
        RECT -24.265 -94.015 -24.035 -93.015 ;
        RECT -23.775 -94.015 -23.545 -93.015 ;
        RECT -23.175 -94.015 -22.945 -93.015 ;
        RECT -22.685 -94.015 -22.455 -93.015 ;
        RECT -22.195 -94.015 -21.965 -93.015 ;
        RECT -20.385 -94.015 -20.155 -93.015 ;
        RECT -19.405 -94.015 -19.175 -93.015 ;
        RECT -17.855 -94.015 -17.625 -93.015 ;
        RECT -16.310 -94.015 -16.080 -93.015 ;
        RECT -12.255 -94.015 -12.025 -93.015 ;
        RECT -11.765 -94.015 -11.535 -93.015 ;
        RECT -11.275 -94.015 -11.045 -93.015 ;
        RECT -10.675 -94.015 -10.445 -93.015 ;
        RECT -10.185 -94.015 -9.955 -93.015 ;
        RECT -9.695 -94.015 -9.465 -93.015 ;
        RECT -7.885 -94.015 -7.655 -93.015 ;
        RECT -6.905 -94.015 -6.675 -93.015 ;
        RECT -5.355 -94.015 -5.125 -93.015 ;
        RECT -3.810 -94.015 -3.580 -93.015 ;
        RECT 0.245 -94.015 0.475 -93.015 ;
        RECT 0.735 -94.015 0.965 -93.015 ;
        RECT 1.225 -94.015 1.455 -93.015 ;
        RECT 1.825 -94.015 2.055 -93.015 ;
        RECT 2.315 -94.015 2.545 -93.015 ;
        RECT 2.805 -94.015 3.035 -93.015 ;
        RECT 4.615 -94.015 4.845 -93.015 ;
        RECT 5.595 -94.015 5.825 -93.015 ;
        RECT 7.145 -94.015 7.375 -93.015 ;
        RECT 8.690 -94.015 8.920 -93.015 ;
        RECT 12.745 -94.015 12.975 -93.015 ;
        RECT 13.235 -94.015 13.465 -93.015 ;
        RECT 13.725 -94.015 13.955 -93.015 ;
        RECT 14.325 -94.015 14.555 -93.015 ;
        RECT 14.815 -94.015 15.045 -93.015 ;
        RECT 15.305 -94.015 15.535 -93.015 ;
        RECT 17.115 -94.015 17.345 -93.015 ;
        RECT 18.095 -94.015 18.325 -93.015 ;
        RECT 19.645 -94.015 19.875 -93.015 ;
        RECT 21.190 -94.015 21.420 -93.015 ;
        RECT 27.745 -94.015 27.975 -93.015 ;
        RECT 28.235 -94.015 28.465 -93.015 ;
        RECT 28.725 -94.015 28.955 -93.015 ;
        RECT 29.325 -94.015 29.555 -93.015 ;
        RECT 29.815 -94.015 30.045 -93.015 ;
        RECT 30.305 -94.015 30.535 -93.015 ;
        RECT 32.115 -94.015 32.345 -93.015 ;
        RECT 33.095 -94.015 33.325 -93.015 ;
        RECT 34.645 -94.015 34.875 -93.015 ;
        RECT 36.190 -94.015 36.420 -93.015 ;
        RECT -31.440 -94.655 -30.745 -94.565 ;
        RECT -28.365 -94.655 -27.670 -94.595 ;
        RECT -18.940 -94.655 -18.245 -94.565 ;
        RECT -15.865 -94.655 -15.170 -94.595 ;
        RECT -6.440 -94.655 -5.745 -94.565 ;
        RECT -3.365 -94.655 -2.670 -94.595 ;
        RECT 6.060 -94.655 6.755 -94.565 ;
        RECT 9.135 -94.655 9.830 -94.595 ;
        RECT 18.560 -94.655 19.255 -94.565 ;
        RECT 21.635 -94.655 22.330 -94.595 ;
        RECT 33.560 -94.655 34.255 -94.565 ;
        RECT 36.635 -94.655 37.330 -94.595 ;
        RECT 40.140 -94.655 41.140 -92.895 ;
        RECT -37.230 -94.850 -36.535 -94.785 ;
        RECT -31.440 -94.795 -26.915 -94.655 ;
        RECT -31.440 -94.835 -30.745 -94.795 ;
        RECT -37.230 -94.990 -35.460 -94.850 ;
        RECT -28.365 -94.865 -27.670 -94.795 ;
        RECT -37.230 -95.055 -36.535 -94.990 ;
        RECT -58.020 -96.440 -54.220 -96.210 ;
        RECT -49.995 -96.380 -49.335 -96.080 ;
        RECT -48.295 -96.330 -45.145 -95.855 ;
        RECT -61.605 -96.870 -60.920 -96.570 ;
        RECT -58.020 -96.925 -57.790 -96.440 ;
        RECT -57.045 -96.925 -56.835 -96.440 ;
        RECT -56.070 -96.925 -55.860 -96.440 ;
        RECT -55.090 -96.925 -54.880 -96.440 ;
        RECT -62.925 -97.625 -62.620 -97.400 ;
        RECT -62.925 -98.060 -62.625 -97.625 ;
        RECT -62.225 -97.675 -61.995 -97.175 ;
        RECT -61.735 -97.675 -61.505 -97.175 ;
        RECT -61.245 -97.675 -61.015 -97.175 ;
        RECT -60.755 -97.675 -60.525 -97.175 ;
        RECT -60.265 -97.675 -60.035 -97.175 ;
        RECT -59.775 -97.675 -59.545 -97.175 ;
        RECT -58.035 -97.425 -57.790 -96.925 ;
        RECT -57.545 -97.425 -57.315 -96.925 ;
        RECT -57.055 -97.425 -56.825 -96.925 ;
        RECT -56.565 -97.425 -56.335 -96.925 ;
        RECT -56.075 -97.425 -55.845 -96.925 ;
        RECT -55.585 -97.425 -55.355 -96.925 ;
        RECT -55.095 -97.425 -54.865 -96.925 ;
        RECT -54.605 -97.425 -54.375 -96.925 ;
        RECT -53.510 -97.675 -53.280 -97.175 ;
        RECT -53.020 -97.675 -52.790 -97.175 ;
        RECT -52.530 -97.675 -52.300 -97.175 ;
        RECT -52.040 -97.675 -51.810 -97.175 ;
        RECT -51.550 -97.675 -51.320 -97.175 ;
        RECT -51.060 -97.675 -50.830 -97.175 ;
        RECT -49.830 -97.520 -49.540 -96.380 ;
        RECT -48.295 -96.575 -47.820 -96.330 ;
        RECT -48.470 -96.875 -47.785 -96.575 ;
        RECT -55.235 -98.025 -54.390 -97.990 ;
        RECT -68.735 -98.360 -67.890 -98.310 ;
        RECT -75.725 -99.575 -75.495 -98.575 ;
        RECT -74.745 -99.575 -74.515 -98.575 ;
        RECT -73.765 -99.575 -73.535 -98.575 ;
        RECT -71.535 -99.340 -71.305 -99.000 ;
        RECT -71.535 -99.500 -71.280 -99.340 ;
        RECT -71.045 -99.500 -70.815 -99.000 ;
        RECT -70.555 -99.215 -70.325 -99.000 ;
        RECT -71.530 -99.915 -71.280 -99.500 ;
        RECT -70.575 -99.915 -70.320 -99.215 ;
        RECT -70.065 -99.500 -69.835 -99.000 ;
        RECT -69.575 -99.310 -69.345 -99.000 ;
        RECT -69.575 -99.915 -69.320 -99.310 ;
        RECT -69.085 -99.500 -68.855 -99.000 ;
        RECT -68.595 -99.310 -68.365 -99.000 ;
        RECT -68.605 -99.915 -68.350 -99.310 ;
        RECT -68.105 -99.500 -67.875 -99.000 ;
        RECT -67.010 -99.575 -66.780 -98.575 ;
        RECT -66.030 -99.575 -65.800 -98.575 ;
        RECT -65.050 -99.575 -64.820 -98.575 ;
        RECT -64.030 -99.485 -63.745 -98.310 ;
        RECT -55.235 -98.310 -50.245 -98.025 ;
        RECT -49.840 -98.180 -49.540 -97.520 ;
        RECT -49.100 -97.675 -48.870 -97.175 ;
        RECT -48.610 -97.675 -48.380 -97.175 ;
        RECT -48.120 -97.675 -47.890 -97.175 ;
        RECT -47.630 -97.675 -47.400 -97.175 ;
        RECT -47.140 -97.675 -46.910 -97.175 ;
        RECT -46.650 -97.675 -46.420 -97.175 ;
        RECT -55.235 -98.360 -54.390 -98.310 ;
        RECT -62.225 -99.575 -61.995 -98.575 ;
        RECT -61.245 -99.575 -61.015 -98.575 ;
        RECT -60.265 -99.575 -60.035 -98.575 ;
        RECT -58.035 -99.500 -57.805 -99.000 ;
        RECT -57.545 -99.500 -57.315 -99.000 ;
        RECT -57.055 -99.500 -56.825 -99.000 ;
        RECT -56.565 -99.500 -56.335 -99.000 ;
        RECT -56.075 -99.500 -55.845 -99.000 ;
        RECT -55.585 -99.500 -55.355 -99.000 ;
        RECT -55.095 -99.500 -54.865 -99.000 ;
        RECT -54.605 -99.500 -54.375 -99.000 ;
        RECT -53.510 -99.575 -53.280 -98.575 ;
        RECT -52.530 -99.575 -52.300 -98.575 ;
        RECT -51.550 -99.575 -51.320 -98.575 ;
        RECT -50.530 -99.915 -50.245 -98.310 ;
        RECT -49.100 -99.575 -48.870 -98.575 ;
        RECT -48.120 -99.575 -47.890 -98.575 ;
        RECT -47.140 -99.575 -46.910 -98.575 ;
        RECT -71.530 -100.200 -50.245 -99.915 ;
        RECT -45.620 -101.000 -45.145 -96.330 ;
        RECT -43.990 -98.095 -43.760 -96.595 ;
        RECT -43.500 -98.095 -43.270 -96.595 ;
        RECT -42.290 -98.095 -42.060 -96.595 ;
        RECT -41.800 -98.095 -41.570 -96.595 ;
        RECT -41.310 -98.095 -41.080 -96.595 ;
        RECT -59.980 -101.565 -45.140 -101.000 ;
        RECT -70.605 -103.355 -68.410 -103.120 ;
        RECT -70.605 -103.540 -70.370 -103.355 ;
        RECT -70.600 -105.035 -70.370 -103.540 ;
        RECT -70.110 -105.035 -69.880 -103.535 ;
        RECT -69.620 -105.035 -69.390 -103.355 ;
        RECT -73.295 -105.690 -72.365 -105.480 ;
        RECT -77.605 -106.010 -72.365 -105.690 ;
        RECT -73.295 -106.250 -72.365 -106.010 ;
        RECT -85.080 -108.230 -81.540 -107.665 ;
        RECT -70.110 -107.720 -69.880 -106.220 ;
        RECT -69.130 -107.720 -68.900 -103.535 ;
        RECT -68.640 -105.035 -68.410 -103.355 ;
        RECT -62.875 -103.605 -62.645 -102.105 ;
        RECT -62.385 -103.605 -62.155 -102.105 ;
        RECT -61.895 -103.605 -61.665 -102.105 ;
        RECT -60.685 -103.605 -60.455 -102.105 ;
        RECT -60.195 -103.605 -59.965 -102.105 ;
        RECT -63.370 -104.095 -58.270 -103.770 ;
        RECT -58.595 -104.510 -58.270 -104.095 ;
        RECT -58.625 -104.870 -58.100 -104.510 ;
        RECT -67.065 -106.570 -66.835 -106.070 ;
        RECT -66.575 -106.715 -66.345 -106.070 ;
        RECT -66.085 -106.570 -65.855 -106.070 ;
        RECT -65.595 -106.715 -65.365 -106.070 ;
        RECT -67.065 -106.945 -63.880 -106.715 ;
        RECT -67.065 -107.725 -66.835 -106.945 ;
        RECT -66.575 -106.955 -65.365 -106.945 ;
        RECT -66.085 -107.725 -65.855 -106.955 ;
        RECT -65.105 -107.725 -64.875 -106.945 ;
        RECT -62.875 -108.165 -62.645 -105.165 ;
        RECT -61.820 -108.165 -61.590 -105.165 ;
        RECT -61.330 -108.165 -61.100 -105.165 ;
        RECT -60.840 -108.165 -60.610 -105.165 ;
        RECT -59.780 -108.165 -59.550 -105.165 ;
        RECT -88.590 -110.205 -88.360 -108.525 ;
        RECT -90.555 -110.440 -88.360 -110.205 ;
        RECT -85.495 -111.985 -84.155 -110.660 ;
        RECT -85.250 -114.760 -84.310 -111.985 ;
        RECT -85.470 -116.085 -84.130 -114.760 ;
        RECT -82.105 -121.120 -81.540 -108.230 ;
        RECT -69.980 -112.645 -69.750 -111.365 ;
        RECT -69.000 -112.635 -68.770 -111.365 ;
        RECT -69.490 -112.645 -68.280 -112.635 ;
        RECT -68.020 -112.645 -67.790 -111.365 ;
        RECT -65.115 -112.220 -64.885 -110.720 ;
        RECT -84.925 -121.685 -81.540 -121.120 ;
        RECT -112.620 -125.045 -112.390 -122.045 ;
        RECT -111.560 -125.045 -111.330 -122.045 ;
        RECT -111.070 -125.045 -110.840 -122.045 ;
        RECT -110.580 -125.045 -110.350 -122.045 ;
        RECT -110.015 -125.045 -109.785 -122.045 ;
        RECT -109.525 -125.045 -109.295 -122.045 ;
        RECT -109.035 -125.045 -108.805 -122.045 ;
        RECT -106.590 -123.690 -106.360 -121.690 ;
        RECT -105.535 -123.690 -105.305 -121.690 ;
        RECT -105.045 -123.690 -104.815 -121.690 ;
        RECT -104.555 -123.690 -104.325 -121.690 ;
        RECT -102.065 -123.695 -101.835 -121.695 ;
        RECT -101.010 -123.695 -100.780 -121.695 ;
        RECT -100.520 -123.695 -100.290 -121.695 ;
        RECT -100.030 -123.695 -99.800 -121.695 ;
        RECT -95.550 -123.475 -93.355 -123.240 ;
        RECT -95.550 -123.660 -95.315 -123.475 ;
        RECT -104.495 -124.930 -103.810 -124.640 ;
        RECT -106.590 -126.150 -106.360 -125.150 ;
        RECT -106.100 -126.150 -105.870 -125.150 ;
        RECT -105.610 -126.150 -105.380 -125.150 ;
        RECT -108.930 -126.675 -108.245 -126.385 ;
        RECT -112.620 -127.865 -112.390 -126.865 ;
        RECT -112.130 -127.865 -111.900 -126.865 ;
        RECT -111.640 -127.865 -111.410 -126.865 ;
        RECT -111.150 -127.865 -110.920 -126.865 ;
        RECT -113.290 -129.095 -109.270 -128.345 ;
        RECT -113.230 -131.155 -112.795 -129.095 ;
        RECT -112.330 -131.155 -111.895 -129.095 ;
        RECT -111.465 -131.155 -111.030 -129.095 ;
        RECT -110.545 -131.155 -110.110 -129.095 ;
        RECT -109.920 -131.155 -109.485 -129.095 ;
        RECT -114.355 -131.730 -109.440 -131.155 ;
        RECT -108.870 -131.665 -108.420 -126.675 ;
        RECT -108.870 -132.115 -107.285 -131.665 ;
        RECT -114.305 -133.595 -114.075 -132.595 ;
        RECT -113.815 -133.595 -113.585 -132.595 ;
        RECT -112.240 -134.095 -112.010 -132.595 ;
        RECT -111.750 -134.095 -111.520 -132.595 ;
        RECT -111.260 -134.095 -111.030 -132.595 ;
        RECT -110.695 -134.095 -110.465 -132.595 ;
        RECT -110.205 -134.095 -109.975 -132.595 ;
        RECT -109.715 -134.095 -109.485 -132.595 ;
        RECT -109.145 -134.100 -108.915 -132.600 ;
        RECT -108.655 -134.100 -108.425 -132.600 ;
        RECT -108.165 -134.100 -107.935 -132.600 ;
        RECT -107.735 -135.055 -107.285 -132.115 ;
        RECT -104.040 -134.780 -103.865 -124.930 ;
        RECT -99.840 -124.935 -99.155 -124.645 ;
        RECT -102.065 -126.155 -101.835 -125.155 ;
        RECT -101.575 -126.155 -101.345 -125.155 ;
        RECT -101.085 -126.155 -100.855 -125.155 ;
        RECT -104.080 -135.465 -103.790 -134.780 ;
        RECT -99.415 -135.210 -99.240 -124.935 ;
        RECT -95.545 -125.155 -95.315 -123.660 ;
        RECT -95.055 -125.155 -94.825 -123.655 ;
        RECT -94.565 -125.155 -94.335 -123.475 ;
        RECT -96.820 -125.635 -95.835 -125.365 ;
        RECT -98.535 -126.425 -97.950 -125.810 ;
        RECT -99.030 -133.450 -98.740 -132.765 ;
        RECT -99.455 -135.895 -99.165 -135.210 ;
        RECT -114.305 -137.135 -114.075 -136.135 ;
        RECT -110.615 -137.135 -110.385 -136.135 ;
        RECT -109.635 -137.135 -109.405 -136.135 ;
        RECT -108.655 -137.135 -108.425 -136.135 ;
        RECT -114.300 -138.490 -114.085 -137.135 ;
        RECT -114.550 -139.070 -113.760 -138.490 ;
        RECT -99.025 -138.630 -98.830 -133.450 ;
        RECT -98.520 -137.745 -98.060 -126.425 ;
        RECT -96.105 -132.655 -95.835 -125.635 ;
        RECT -95.055 -127.840 -94.825 -126.340 ;
        RECT -94.075 -127.840 -93.845 -123.655 ;
        RECT -93.585 -125.155 -93.355 -123.475 ;
        RECT -87.820 -123.725 -87.590 -122.225 ;
        RECT -87.330 -123.725 -87.100 -122.225 ;
        RECT -86.840 -123.725 -86.610 -122.225 ;
        RECT -85.630 -123.725 -85.400 -122.225 ;
        RECT -85.140 -123.725 -84.910 -122.225 ;
        RECT -88.315 -124.215 -83.215 -123.890 ;
        RECT -83.540 -124.630 -83.215 -124.215 ;
        RECT -83.570 -124.990 -83.045 -124.630 ;
        RECT -92.010 -126.690 -91.780 -126.190 ;
        RECT -91.520 -126.835 -91.290 -126.190 ;
        RECT -91.030 -126.690 -90.800 -126.190 ;
        RECT -90.540 -126.835 -90.310 -126.190 ;
        RECT -92.010 -127.065 -88.825 -126.835 ;
        RECT -92.010 -127.845 -91.780 -127.065 ;
        RECT -91.520 -127.075 -90.310 -127.065 ;
        RECT -91.030 -127.845 -90.800 -127.075 ;
        RECT -90.050 -127.845 -89.820 -127.065 ;
        RECT -87.820 -128.285 -87.590 -125.285 ;
        RECT -86.765 -128.285 -86.535 -125.285 ;
        RECT -86.275 -128.285 -86.045 -125.285 ;
        RECT -85.785 -128.285 -85.555 -125.285 ;
        RECT -84.725 -128.285 -84.495 -125.285 ;
        RECT -96.355 -133.405 -95.705 -132.655 ;
        RECT -94.925 -132.765 -94.695 -131.485 ;
        RECT -93.945 -132.755 -93.715 -131.485 ;
        RECT -94.435 -132.765 -93.225 -132.755 ;
        RECT -92.965 -132.765 -92.735 -131.485 ;
        RECT -90.060 -132.340 -89.830 -130.840 ;
        RECT -94.925 -132.995 -91.740 -132.765 ;
        RECT -91.030 -132.860 -90.235 -132.570 ;
        RECT -94.925 -134.135 -94.695 -133.135 ;
        RECT -94.435 -134.135 -94.205 -132.995 ;
        RECT -93.945 -134.135 -93.715 -133.135 ;
        RECT -93.455 -134.135 -93.225 -132.995 ;
        RECT -90.900 -133.135 -90.630 -132.860 ;
        RECT -92.270 -133.405 -90.630 -133.135 ;
        RECT -92.270 -134.855 -92.000 -133.405 ;
        RECT -97.485 -135.125 -92.000 -134.855 ;
        RECT -90.550 -135.020 -90.320 -133.525 ;
        RECT -97.485 -136.475 -97.215 -135.125 ;
        RECT -90.555 -135.205 -90.320 -135.020 ;
        RECT -90.060 -135.025 -89.830 -133.525 ;
        RECT -89.570 -135.205 -89.340 -133.525 ;
        RECT -89.080 -135.025 -88.850 -130.840 ;
        RECT -87.015 -131.615 -86.785 -130.835 ;
        RECT -86.035 -131.605 -85.805 -130.835 ;
        RECT -86.525 -131.615 -85.315 -131.605 ;
        RECT -85.055 -131.615 -84.825 -130.835 ;
        RECT -87.015 -131.845 -83.830 -131.615 ;
        RECT -87.015 -132.490 -86.785 -131.990 ;
        RECT -86.525 -132.490 -86.295 -131.845 ;
        RECT -86.035 -132.490 -85.805 -131.990 ;
        RECT -85.545 -132.490 -85.315 -131.845 ;
        RECT -82.105 -132.665 -81.540 -121.685 ;
        RECT -80.775 -124.645 -79.735 -112.665 ;
        RECT -69.980 -112.875 -66.795 -112.645 ;
        RECT -66.085 -112.740 -65.290 -112.450 ;
        RECT -69.980 -114.015 -69.750 -113.015 ;
        RECT -69.490 -114.015 -69.260 -112.875 ;
        RECT -69.000 -114.015 -68.770 -113.015 ;
        RECT -68.510 -114.015 -68.280 -112.875 ;
        RECT -65.955 -113.015 -65.685 -112.740 ;
        RECT -67.325 -113.285 -65.685 -113.015 ;
        RECT -67.325 -114.735 -67.055 -113.285 ;
        RECT -77.895 -115.005 -67.055 -114.735 ;
        RECT -65.605 -114.900 -65.375 -113.405 ;
        RECT -77.895 -120.425 -77.625 -115.005 ;
        RECT -65.610 -115.085 -65.375 -114.900 ;
        RECT -65.115 -114.905 -64.885 -113.405 ;
        RECT -64.625 -115.085 -64.395 -113.405 ;
        RECT -64.135 -114.905 -63.905 -110.720 ;
        RECT -62.070 -111.495 -61.840 -110.715 ;
        RECT -61.090 -111.485 -60.860 -110.715 ;
        RECT -61.580 -111.495 -60.370 -111.485 ;
        RECT -60.110 -111.495 -59.880 -110.715 ;
        RECT -62.070 -111.725 -58.885 -111.495 ;
        RECT -62.070 -112.370 -61.840 -111.870 ;
        RECT -61.580 -112.370 -61.350 -111.725 ;
        RECT -61.090 -112.370 -60.860 -111.870 ;
        RECT -60.600 -112.370 -60.370 -111.725 ;
        RECT -57.160 -112.545 -56.595 -101.565 ;
        RECT -60.135 -113.110 -56.595 -112.545 ;
        RECT -63.645 -115.085 -63.415 -113.405 ;
        RECT -65.610 -115.320 -63.415 -115.085 ;
        RECT -75.235 -117.620 -75.005 -116.620 ;
        RECT -74.255 -117.620 -74.025 -116.620 ;
        RECT -73.275 -117.620 -73.045 -116.620 ;
        RECT -72.125 -117.885 -71.840 -116.710 ;
        RECT -71.050 -117.620 -70.820 -116.620 ;
        RECT -70.070 -117.620 -69.840 -116.620 ;
        RECT -69.090 -117.620 -68.860 -116.620 ;
        RECT -67.995 -117.195 -67.765 -116.695 ;
        RECT -67.505 -117.195 -67.275 -116.695 ;
        RECT -67.015 -117.195 -66.785 -116.695 ;
        RECT -66.525 -117.195 -66.295 -116.695 ;
        RECT -66.035 -117.195 -65.805 -116.695 ;
        RECT -65.545 -117.195 -65.315 -116.695 ;
        RECT -65.055 -117.195 -64.825 -116.695 ;
        RECT -64.565 -117.195 -64.335 -116.695 ;
        RECT -61.735 -117.620 -61.505 -116.620 ;
        RECT -60.755 -117.620 -60.525 -116.620 ;
        RECT -59.775 -117.620 -59.545 -116.620 ;
        RECT -67.980 -117.885 -67.135 -117.835 ;
        RECT -72.125 -118.170 -67.135 -117.885 ;
        RECT -58.625 -117.885 -58.340 -116.710 ;
        RECT -57.550 -117.620 -57.320 -116.620 ;
        RECT -56.570 -117.620 -56.340 -116.620 ;
        RECT -55.590 -117.620 -55.360 -116.620 ;
        RECT -54.495 -117.195 -54.265 -116.695 ;
        RECT -54.005 -117.195 -53.775 -116.695 ;
        RECT -53.515 -117.195 -53.285 -116.695 ;
        RECT -53.025 -117.195 -52.795 -116.695 ;
        RECT -52.535 -117.195 -52.305 -116.695 ;
        RECT -52.045 -117.195 -51.815 -116.695 ;
        RECT -51.555 -117.195 -51.325 -116.695 ;
        RECT -51.065 -117.195 -50.835 -116.695 ;
        RECT -54.480 -117.885 -53.635 -117.835 ;
        RECT -62.920 -117.995 -62.620 -117.965 ;
        RECT -64.095 -118.100 -63.890 -118.095 ;
        RECT -67.980 -118.205 -67.135 -118.170 ;
        RECT -75.725 -119.020 -75.495 -118.520 ;
        RECT -75.235 -119.020 -75.005 -118.520 ;
        RECT -74.745 -119.020 -74.515 -118.520 ;
        RECT -74.255 -119.020 -74.025 -118.520 ;
        RECT -73.765 -119.020 -73.535 -118.520 ;
        RECT -73.275 -119.020 -73.045 -118.520 ;
        RECT -74.555 -120.135 -73.870 -119.835 ;
        RECT -76.295 -120.425 -75.995 -120.190 ;
        RECT -77.895 -120.745 -75.995 -120.425 ;
        RECT -76.295 -120.875 -75.995 -120.745 ;
        RECT -74.480 -121.225 -74.005 -120.135 ;
        RECT -72.430 -120.725 -72.130 -118.390 ;
        RECT -64.570 -118.400 -63.885 -118.100 ;
        RECT -62.920 -118.295 -62.205 -117.995 ;
        RECT -58.625 -118.170 -53.635 -117.885 ;
        RECT -54.480 -118.205 -53.635 -118.170 ;
        RECT -71.540 -119.020 -71.310 -118.520 ;
        RECT -71.050 -119.020 -70.820 -118.520 ;
        RECT -70.560 -119.020 -70.330 -118.520 ;
        RECT -70.070 -119.020 -69.840 -118.520 ;
        RECT -69.580 -119.020 -69.350 -118.520 ;
        RECT -69.090 -119.020 -68.860 -118.520 ;
        RECT -67.995 -119.270 -67.765 -118.770 ;
        RECT -67.505 -119.270 -67.275 -118.770 ;
        RECT -67.015 -119.270 -66.785 -118.770 ;
        RECT -66.525 -119.270 -66.295 -118.770 ;
        RECT -66.035 -119.270 -65.805 -118.770 ;
        RECT -65.545 -119.270 -65.315 -118.770 ;
        RECT -65.055 -119.270 -64.825 -118.770 ;
        RECT -64.565 -119.270 -64.335 -118.770 ;
        RECT -72.610 -121.025 -71.950 -120.725 ;
        RECT -64.095 -120.825 -63.890 -118.400 ;
        RECT -63.745 -120.580 -63.060 -120.280 ;
        RECT -71.545 -121.065 -63.890 -120.825 ;
        RECT -74.600 -121.525 -73.940 -121.225 ;
        RECT -75.725 -122.310 -75.495 -121.810 ;
        RECT -75.235 -122.310 -75.005 -121.810 ;
        RECT -74.745 -122.310 -74.515 -121.810 ;
        RECT -74.255 -122.310 -74.025 -121.810 ;
        RECT -73.765 -122.310 -73.535 -121.810 ;
        RECT -73.275 -122.310 -73.045 -121.810 ;
        RECT -71.545 -121.835 -71.305 -121.065 ;
        RECT -71.535 -122.060 -71.305 -121.835 ;
        RECT -71.045 -122.060 -70.815 -121.560 ;
        RECT -70.585 -121.655 -70.280 -121.065 ;
        RECT -70.555 -122.060 -70.325 -121.655 ;
        RECT -70.065 -122.060 -69.835 -121.560 ;
        RECT -69.605 -121.665 -69.300 -121.065 ;
        RECT -69.575 -122.060 -69.345 -121.665 ;
        RECT -69.085 -122.060 -68.855 -121.560 ;
        RECT -68.650 -121.655 -68.345 -121.065 ;
        RECT -68.595 -122.060 -68.365 -121.655 ;
        RECT -68.105 -122.060 -67.875 -121.560 ;
        RECT -67.010 -122.310 -66.780 -121.810 ;
        RECT -66.520 -122.310 -66.290 -121.810 ;
        RECT -66.030 -122.310 -65.800 -121.810 ;
        RECT -65.540 -122.310 -65.310 -121.810 ;
        RECT -65.050 -122.310 -64.820 -121.810 ;
        RECT -64.560 -122.310 -64.330 -121.810 ;
        RECT -68.735 -122.660 -67.890 -122.625 ;
        RECT -68.735 -122.945 -63.745 -122.660 ;
        RECT -63.500 -122.820 -63.200 -120.580 ;
        RECT -62.920 -122.035 -62.620 -118.295 ;
        RECT -51.125 -118.410 -50.355 -118.110 ;
        RECT -62.225 -119.020 -61.995 -118.520 ;
        RECT -61.735 -119.020 -61.505 -118.520 ;
        RECT -61.245 -119.020 -61.015 -118.520 ;
        RECT -60.755 -119.020 -60.525 -118.520 ;
        RECT -60.265 -119.020 -60.035 -118.520 ;
        RECT -59.775 -119.020 -59.545 -118.520 ;
        RECT -61.570 -120.165 -60.885 -119.865 ;
        RECT -61.515 -121.205 -61.040 -120.165 ;
        RECT -58.870 -120.285 -58.570 -118.465 ;
        RECT -58.040 -119.020 -57.810 -118.520 ;
        RECT -57.550 -119.020 -57.320 -118.520 ;
        RECT -57.060 -119.020 -56.830 -118.520 ;
        RECT -56.570 -119.020 -56.340 -118.520 ;
        RECT -56.080 -119.020 -55.850 -118.520 ;
        RECT -55.590 -119.020 -55.360 -118.520 ;
        RECT -54.495 -119.270 -54.265 -118.770 ;
        RECT -54.005 -119.270 -53.775 -118.770 ;
        RECT -53.515 -119.270 -53.285 -118.770 ;
        RECT -53.025 -119.270 -52.795 -118.770 ;
        RECT -52.535 -119.270 -52.305 -118.770 ;
        RECT -52.045 -119.270 -51.815 -118.770 ;
        RECT -51.555 -119.270 -51.325 -118.770 ;
        RECT -51.065 -119.270 -50.835 -118.770 ;
        RECT -50.585 -119.785 -50.355 -118.410 ;
        RECT -54.450 -120.010 -50.355 -119.785 ;
        RECT -48.295 -119.865 -47.820 -101.565 ;
        RECT -54.450 -120.015 -50.395 -120.010 ;
        RECT -59.015 -120.585 -58.355 -120.285 ;
        RECT -54.450 -120.845 -54.220 -120.015 ;
        RECT -48.380 -120.165 -47.720 -119.865 ;
        RECT -58.020 -121.075 -54.220 -120.845 ;
        RECT -49.995 -121.015 -49.335 -120.715 ;
        RECT -61.605 -121.505 -60.920 -121.205 ;
        RECT -58.020 -121.560 -57.790 -121.075 ;
        RECT -57.045 -121.560 -56.835 -121.075 ;
        RECT -56.070 -121.560 -55.860 -121.075 ;
        RECT -55.090 -121.560 -54.880 -121.075 ;
        RECT -62.925 -122.260 -62.620 -122.035 ;
        RECT -62.925 -122.695 -62.625 -122.260 ;
        RECT -62.225 -122.310 -61.995 -121.810 ;
        RECT -61.735 -122.310 -61.505 -121.810 ;
        RECT -61.245 -122.310 -61.015 -121.810 ;
        RECT -60.755 -122.310 -60.525 -121.810 ;
        RECT -60.265 -122.310 -60.035 -121.810 ;
        RECT -59.775 -122.310 -59.545 -121.810 ;
        RECT -58.035 -122.060 -57.790 -121.560 ;
        RECT -57.545 -122.060 -57.315 -121.560 ;
        RECT -57.055 -122.060 -56.825 -121.560 ;
        RECT -56.565 -122.060 -56.335 -121.560 ;
        RECT -56.075 -122.060 -55.845 -121.560 ;
        RECT -55.585 -122.060 -55.355 -121.560 ;
        RECT -55.095 -122.060 -54.865 -121.560 ;
        RECT -54.605 -122.060 -54.375 -121.560 ;
        RECT -53.510 -122.310 -53.280 -121.810 ;
        RECT -53.020 -122.310 -52.790 -121.810 ;
        RECT -52.530 -122.310 -52.300 -121.810 ;
        RECT -52.040 -122.310 -51.810 -121.810 ;
        RECT -51.550 -122.310 -51.320 -121.810 ;
        RECT -51.060 -122.310 -50.830 -121.810 ;
        RECT -49.830 -122.155 -49.540 -121.015 ;
        RECT -48.295 -121.210 -47.820 -120.165 ;
        RECT -48.470 -121.510 -47.785 -121.210 ;
        RECT -55.235 -122.660 -54.390 -122.625 ;
        RECT -68.735 -122.995 -67.890 -122.945 ;
        RECT -75.725 -124.210 -75.495 -123.210 ;
        RECT -74.745 -124.210 -74.515 -123.210 ;
        RECT -73.765 -124.210 -73.535 -123.210 ;
        RECT -71.535 -123.975 -71.305 -123.635 ;
        RECT -71.535 -124.135 -71.280 -123.975 ;
        RECT -71.045 -124.135 -70.815 -123.635 ;
        RECT -70.555 -123.850 -70.325 -123.635 ;
        RECT -71.530 -124.550 -71.280 -124.135 ;
        RECT -70.575 -124.550 -70.320 -123.850 ;
        RECT -70.065 -124.135 -69.835 -123.635 ;
        RECT -69.575 -123.945 -69.345 -123.635 ;
        RECT -69.575 -124.550 -69.320 -123.945 ;
        RECT -69.085 -124.135 -68.855 -123.635 ;
        RECT -68.595 -123.945 -68.365 -123.635 ;
        RECT -68.605 -124.550 -68.350 -123.945 ;
        RECT -68.105 -124.135 -67.875 -123.635 ;
        RECT -67.010 -124.210 -66.780 -123.210 ;
        RECT -66.030 -124.210 -65.800 -123.210 ;
        RECT -65.050 -124.210 -64.820 -123.210 ;
        RECT -64.030 -124.120 -63.745 -122.945 ;
        RECT -55.235 -122.945 -50.245 -122.660 ;
        RECT -49.840 -122.815 -49.540 -122.155 ;
        RECT -49.100 -122.310 -48.870 -121.810 ;
        RECT -48.610 -122.310 -48.380 -121.810 ;
        RECT -48.120 -122.310 -47.890 -121.810 ;
        RECT -47.630 -122.310 -47.400 -121.810 ;
        RECT -47.140 -122.310 -46.910 -121.810 ;
        RECT -46.650 -122.310 -46.420 -121.810 ;
        RECT -55.235 -122.995 -54.390 -122.945 ;
        RECT -62.225 -124.210 -61.995 -123.210 ;
        RECT -61.245 -124.210 -61.015 -123.210 ;
        RECT -60.265 -124.210 -60.035 -123.210 ;
        RECT -58.035 -124.135 -57.805 -123.635 ;
        RECT -57.545 -124.135 -57.315 -123.635 ;
        RECT -57.055 -124.135 -56.825 -123.635 ;
        RECT -56.565 -124.135 -56.335 -123.635 ;
        RECT -56.075 -124.135 -55.845 -123.635 ;
        RECT -55.585 -124.135 -55.355 -123.635 ;
        RECT -55.095 -124.135 -54.865 -123.635 ;
        RECT -54.605 -124.135 -54.375 -123.635 ;
        RECT -53.510 -124.210 -53.280 -123.210 ;
        RECT -52.530 -124.210 -52.300 -123.210 ;
        RECT -51.550 -124.210 -51.320 -123.210 ;
        RECT -50.530 -124.550 -50.245 -122.945 ;
        RECT -49.100 -124.210 -48.870 -123.210 ;
        RECT -48.120 -124.210 -47.890 -123.210 ;
        RECT -47.140 -124.210 -46.910 -123.210 ;
        RECT -71.530 -124.835 -50.245 -124.550 ;
        RECT -85.080 -133.230 -81.540 -132.665 ;
        RECT -88.590 -135.205 -88.360 -133.525 ;
        RECT -90.555 -135.440 -88.360 -135.205 ;
        RECT -45.665 -136.355 -44.785 -103.780 ;
        RECT -44.270 -119.705 -44.040 -116.705 ;
        RECT -43.210 -119.705 -42.980 -116.705 ;
        RECT -42.720 -119.705 -42.490 -116.705 ;
        RECT -42.230 -119.705 -42.000 -116.705 ;
        RECT -41.175 -119.705 -40.945 -116.705 ;
        RECT -43.855 -122.765 -43.625 -121.265 ;
        RECT -43.365 -122.765 -43.135 -121.265 ;
        RECT -42.155 -122.765 -41.925 -121.265 ;
        RECT -41.665 -122.765 -41.435 -121.265 ;
        RECT -41.175 -122.765 -40.945 -121.265 ;
        RECT -97.635 -137.155 -96.915 -136.475 ;
        RECT -45.730 -137.210 -44.730 -136.355 ;
        RECT -39.990 -137.645 -39.330 -95.285 ;
        RECT -35.600 -95.715 -35.460 -94.990 ;
        RECT -33.485 -94.980 -32.790 -94.935 ;
        RECT -29.300 -94.980 -28.620 -94.935 ;
        RECT -33.485 -95.120 -28.620 -94.980 ;
        RECT -33.485 -95.205 -32.790 -95.120 ;
        RECT -29.300 -95.165 -28.620 -95.120 ;
        RECT -35.320 -95.350 -34.625 -95.305 ;
        RECT -29.930 -95.340 -29.235 -95.335 ;
        RECT -29.930 -95.350 -27.275 -95.340 ;
        RECT -35.320 -95.480 -27.275 -95.350 ;
        RECT -35.320 -95.490 -29.235 -95.480 ;
        RECT -35.320 -95.575 -34.625 -95.490 ;
        RECT -29.930 -95.605 -29.235 -95.490 ;
        RECT -30.830 -95.715 -30.175 -95.655 ;
        RECT -35.600 -95.855 -30.175 -95.715 ;
        RECT -30.830 -95.885 -30.175 -95.855 ;
        RECT -37.255 -97.045 -37.025 -96.045 ;
        RECT -36.765 -97.045 -36.535 -96.045 ;
        RECT -35.185 -97.045 -34.955 -96.045 ;
        RECT -34.695 -97.045 -34.465 -96.045 ;
        RECT -33.375 -97.045 -33.145 -96.045 ;
        RECT -32.885 -97.045 -32.655 -96.045 ;
        RECT -31.905 -97.045 -31.675 -96.045 ;
        RECT -31.415 -97.045 -31.185 -96.045 ;
        RECT -30.355 -97.045 -30.125 -96.045 ;
        RECT -29.865 -97.045 -29.635 -96.045 ;
        RECT -28.810 -97.045 -28.580 -96.045 ;
        RECT -28.320 -97.045 -28.090 -96.045 ;
        RECT -35.070 -98.760 -34.840 -98.260 ;
        RECT -34.580 -98.760 -34.350 -98.260 ;
        RECT -34.090 -98.760 -33.860 -98.260 ;
        RECT -33.600 -98.760 -33.370 -98.260 ;
        RECT -33.110 -98.760 -32.880 -98.260 ;
        RECT -32.620 -98.760 -32.390 -98.260 ;
        RECT -27.415 -98.675 -27.275 -95.480 ;
        RECT -27.505 -99.355 -27.275 -98.675 ;
        RECT -34.580 -100.660 -34.350 -99.660 ;
        RECT -33.600 -100.660 -33.370 -99.660 ;
        RECT -32.620 -100.660 -32.390 -99.660 ;
        RECT -27.055 -100.835 -26.915 -94.795 ;
        RECT -24.730 -94.850 -24.035 -94.785 ;
        RECT -18.940 -94.795 -14.060 -94.655 ;
        RECT -18.940 -94.835 -18.245 -94.795 ;
        RECT -24.730 -94.990 -22.960 -94.850 ;
        RECT -15.865 -94.865 -15.170 -94.795 ;
        RECT -24.730 -95.055 -24.035 -94.990 ;
        RECT -23.100 -95.715 -22.960 -94.990 ;
        RECT -20.985 -94.980 -20.290 -94.935 ;
        RECT -16.800 -94.980 -16.120 -94.935 ;
        RECT -20.985 -95.120 -16.120 -94.980 ;
        RECT -20.985 -95.205 -20.290 -95.120 ;
        RECT -16.800 -95.165 -16.120 -95.120 ;
        RECT -18.330 -95.715 -17.675 -95.655 ;
        RECT -23.100 -95.855 -17.675 -95.715 ;
        RECT -18.330 -95.885 -17.675 -95.855 ;
        RECT -25.595 -96.880 -25.365 -96.200 ;
        RECT -25.590 -99.730 -25.370 -96.880 ;
        RECT -24.755 -97.045 -24.525 -96.045 ;
        RECT -24.265 -97.045 -24.035 -96.045 ;
        RECT -22.685 -97.045 -22.455 -96.045 ;
        RECT -22.195 -97.045 -21.965 -96.045 ;
        RECT -20.875 -97.045 -20.645 -96.045 ;
        RECT -20.385 -97.045 -20.155 -96.045 ;
        RECT -19.405 -97.045 -19.175 -96.045 ;
        RECT -18.915 -97.045 -18.685 -96.045 ;
        RECT -17.855 -97.045 -17.625 -96.045 ;
        RECT -17.365 -97.045 -17.135 -96.045 ;
        RECT -16.310 -97.045 -16.080 -96.045 ;
        RECT -15.820 -97.045 -15.590 -96.045 ;
        RECT -25.595 -100.410 -25.365 -99.730 ;
        RECT -14.200 -100.085 -14.060 -94.795 ;
        RECT -12.230 -94.850 -11.535 -94.785 ;
        RECT -6.440 -94.795 -1.700 -94.655 ;
        RECT -6.440 -94.835 -5.745 -94.795 ;
        RECT -12.230 -94.990 -10.460 -94.850 ;
        RECT -3.365 -94.865 -2.670 -94.795 ;
        RECT -12.230 -95.055 -11.535 -94.990 ;
        RECT -10.600 -95.715 -10.460 -94.990 ;
        RECT -8.485 -94.980 -7.790 -94.935 ;
        RECT -4.300 -94.980 -3.620 -94.935 ;
        RECT -8.485 -95.120 -3.620 -94.980 ;
        RECT -8.485 -95.205 -7.790 -95.120 ;
        RECT -4.300 -95.165 -3.620 -95.120 ;
        RECT -5.830 -95.715 -5.175 -95.655 ;
        RECT -10.600 -95.855 -5.175 -95.715 ;
        RECT -5.830 -95.885 -5.175 -95.855 ;
        RECT -12.855 -96.900 -12.625 -96.220 ;
        RECT -12.850 -98.085 -12.630 -96.900 ;
        RECT -12.255 -97.045 -12.025 -96.045 ;
        RECT -11.765 -97.045 -11.535 -96.045 ;
        RECT -10.185 -97.045 -9.955 -96.045 ;
        RECT -9.695 -97.045 -9.465 -96.045 ;
        RECT -8.375 -97.045 -8.145 -96.045 ;
        RECT -7.885 -97.045 -7.655 -96.045 ;
        RECT -6.905 -97.045 -6.675 -96.045 ;
        RECT -6.415 -97.045 -6.185 -96.045 ;
        RECT -5.355 -97.045 -5.125 -96.045 ;
        RECT -4.865 -97.045 -4.635 -96.045 ;
        RECT -3.810 -97.045 -3.580 -96.045 ;
        RECT -3.320 -97.045 -3.090 -96.045 ;
        RECT -12.030 -98.085 -11.350 -98.080 ;
        RECT -12.855 -98.305 -11.350 -98.085 ;
        RECT -12.030 -98.310 -11.350 -98.305 ;
        RECT -1.840 -99.520 -1.700 -94.795 ;
        RECT 0.270 -94.850 0.965 -94.785 ;
        RECT 6.060 -94.795 10.675 -94.655 ;
        RECT 6.060 -94.835 6.755 -94.795 ;
        RECT 0.270 -94.990 2.040 -94.850 ;
        RECT 9.135 -94.865 9.830 -94.795 ;
        RECT 0.270 -95.055 0.965 -94.990 ;
        RECT 1.900 -95.715 2.040 -94.990 ;
        RECT 4.015 -94.980 4.710 -94.935 ;
        RECT 8.200 -94.980 8.880 -94.935 ;
        RECT 4.015 -95.120 8.880 -94.980 ;
        RECT 4.015 -95.205 4.710 -95.120 ;
        RECT 8.200 -95.165 8.880 -95.120 ;
        RECT 6.670 -95.715 7.325 -95.655 ;
        RECT 1.900 -95.855 7.325 -95.715 ;
        RECT 6.670 -95.885 7.325 -95.855 ;
        RECT -0.455 -96.900 -0.225 -96.220 ;
        RECT -0.450 -98.150 -0.230 -96.900 ;
        RECT 0.245 -97.045 0.475 -96.045 ;
        RECT 0.735 -97.045 0.965 -96.045 ;
        RECT 2.315 -97.045 2.545 -96.045 ;
        RECT 2.805 -97.045 3.035 -96.045 ;
        RECT 4.125 -97.045 4.355 -96.045 ;
        RECT 4.615 -97.045 4.845 -96.045 ;
        RECT 5.595 -97.045 5.825 -96.045 ;
        RECT 6.085 -97.045 6.315 -96.045 ;
        RECT 7.145 -97.045 7.375 -96.045 ;
        RECT 7.635 -97.045 7.865 -96.045 ;
        RECT 8.690 -97.045 8.920 -96.045 ;
        RECT 9.180 -97.045 9.410 -96.045 ;
        RECT 0.455 -98.150 1.135 -98.145 ;
        RECT -0.450 -98.370 1.135 -98.150 ;
        RECT 0.455 -98.375 1.135 -98.370 ;
        RECT 10.535 -98.835 10.675 -94.795 ;
        RECT 12.770 -94.850 13.465 -94.785 ;
        RECT 18.560 -94.795 27.200 -94.655 ;
        RECT 18.560 -94.835 19.255 -94.795 ;
        RECT 12.770 -94.990 14.540 -94.850 ;
        RECT 21.635 -94.865 22.330 -94.795 ;
        RECT 12.770 -95.055 13.465 -94.990 ;
        RECT 14.400 -95.715 14.540 -94.990 ;
        RECT 16.515 -94.980 17.210 -94.935 ;
        RECT 20.700 -94.980 21.380 -94.935 ;
        RECT 16.515 -95.120 21.380 -94.980 ;
        RECT 16.515 -95.205 17.210 -95.120 ;
        RECT 20.700 -95.165 21.380 -95.120 ;
        RECT 19.170 -95.715 19.825 -95.655 ;
        RECT 14.400 -95.855 19.825 -95.715 ;
        RECT 19.170 -95.885 19.825 -95.855 ;
        RECT 11.630 -96.900 11.860 -96.220 ;
        RECT 11.635 -98.460 11.855 -96.900 ;
        RECT 12.745 -97.045 12.975 -96.045 ;
        RECT 13.235 -97.045 13.465 -96.045 ;
        RECT 14.815 -97.045 15.045 -96.045 ;
        RECT 15.305 -97.045 15.535 -96.045 ;
        RECT 16.625 -97.045 16.855 -96.045 ;
        RECT 17.115 -97.045 17.345 -96.045 ;
        RECT 18.095 -97.045 18.325 -96.045 ;
        RECT 18.585 -97.045 18.815 -96.045 ;
        RECT 19.645 -97.045 19.875 -96.045 ;
        RECT 20.135 -97.045 20.365 -96.045 ;
        RECT 21.190 -97.045 21.420 -96.045 ;
        RECT 21.680 -97.045 21.910 -96.045 ;
        RECT 26.155 -96.900 26.385 -96.220 ;
        RECT 26.160 -98.380 26.380 -96.900 ;
        RECT 27.060 -98.170 27.200 -94.795 ;
        RECT 27.770 -94.850 28.465 -94.785 ;
        RECT 33.560 -94.795 47.985 -94.655 ;
        RECT 33.560 -94.835 34.255 -94.795 ;
        RECT 27.770 -94.990 29.540 -94.850 ;
        RECT 36.635 -94.865 37.330 -94.795 ;
        RECT 27.770 -95.055 28.465 -94.990 ;
        RECT 29.400 -95.715 29.540 -94.990 ;
        RECT 31.515 -94.980 32.210 -94.935 ;
        RECT 35.700 -94.980 36.380 -94.935 ;
        RECT 31.515 -95.120 36.380 -94.980 ;
        RECT 31.515 -95.205 32.210 -95.120 ;
        RECT 35.700 -95.165 36.380 -95.120 ;
        RECT 34.170 -95.715 34.825 -95.655 ;
        RECT 29.400 -95.855 34.825 -95.715 ;
        RECT 34.170 -95.885 34.825 -95.855 ;
        RECT 27.745 -97.045 27.975 -96.045 ;
        RECT 28.235 -97.045 28.465 -96.045 ;
        RECT 29.815 -97.045 30.045 -96.045 ;
        RECT 30.305 -97.045 30.535 -96.045 ;
        RECT 31.625 -97.045 31.855 -96.045 ;
        RECT 32.115 -97.045 32.345 -96.045 ;
        RECT 33.095 -97.045 33.325 -96.045 ;
        RECT 33.585 -97.045 33.815 -96.045 ;
        RECT 34.645 -97.045 34.875 -96.045 ;
        RECT 35.135 -97.045 35.365 -96.045 ;
        RECT 36.190 -97.045 36.420 -96.045 ;
        RECT 36.680 -97.045 36.910 -96.045 ;
        RECT 41.200 -98.170 47.160 -97.585 ;
        RECT 27.060 -98.310 47.205 -98.170 ;
        RECT 11.370 -98.690 12.050 -98.460 ;
        RECT 25.895 -98.610 26.575 -98.380 ;
        RECT 10.535 -99.025 46.440 -98.835 ;
        RECT -1.840 -99.660 45.680 -99.520 ;
        RECT -14.200 -100.340 44.885 -100.085 ;
        RECT -27.055 -101.090 44.105 -100.835 ;
        RECT -25.580 -101.685 -24.900 -101.675 ;
        RECT 9.665 -101.685 10.345 -101.665 ;
        RECT -25.580 -101.895 10.345 -101.685 ;
        RECT -25.580 -101.905 -24.900 -101.895 ;
        RECT -37.980 -102.095 -37.300 -102.085 ;
        RECT 9.145 -102.095 9.920 -102.085 ;
        RECT -37.980 -102.305 9.920 -102.095 ;
        RECT -37.980 -102.315 -37.300 -102.305 ;
        RECT 9.145 -102.315 9.920 -102.305 ;
        RECT -6.815 -102.770 43.000 -102.515 ;
        RECT -36.355 -105.175 -36.125 -104.175 ;
        RECT -35.375 -105.175 -35.145 -104.175 ;
        RECT -34.395 -105.175 -34.165 -104.175 ;
        RECT -32.165 -104.750 -31.935 -104.250 ;
        RECT -31.675 -104.750 -31.445 -104.250 ;
        RECT -31.185 -104.750 -30.955 -104.250 ;
        RECT -30.695 -104.750 -30.465 -104.250 ;
        RECT -30.205 -104.750 -29.975 -104.250 ;
        RECT -29.715 -104.750 -29.485 -104.250 ;
        RECT -29.225 -104.750 -28.995 -104.250 ;
        RECT -28.735 -104.750 -28.505 -104.250 ;
        RECT -27.640 -105.175 -27.410 -104.175 ;
        RECT -26.660 -105.175 -26.430 -104.175 ;
        RECT -25.680 -105.175 -25.450 -104.175 ;
        RECT -29.365 -105.440 -28.520 -105.390 ;
        RECT -24.660 -105.440 -24.375 -104.265 ;
        RECT -22.855 -105.175 -22.625 -104.175 ;
        RECT -21.875 -105.175 -21.645 -104.175 ;
        RECT -20.895 -105.175 -20.665 -104.175 ;
        RECT -18.665 -104.750 -18.435 -104.250 ;
        RECT -18.175 -104.750 -17.945 -104.250 ;
        RECT -17.685 -104.750 -17.455 -104.250 ;
        RECT -17.195 -104.750 -16.965 -104.250 ;
        RECT -16.705 -104.750 -16.475 -104.250 ;
        RECT -16.215 -104.750 -15.985 -104.250 ;
        RECT -15.725 -104.750 -15.495 -104.250 ;
        RECT -15.235 -104.750 -15.005 -104.250 ;
        RECT -14.140 -105.175 -13.910 -104.175 ;
        RECT -13.160 -105.175 -12.930 -104.175 ;
        RECT -12.180 -105.175 -11.950 -104.175 ;
        RECT -29.365 -105.725 -24.375 -105.440 ;
        RECT -15.865 -105.440 -15.020 -105.390 ;
        RECT -11.160 -105.440 -10.875 -104.265 ;
        RECT -9.730 -105.175 -9.500 -104.175 ;
        RECT -8.750 -105.175 -8.520 -104.175 ;
        RECT -7.770 -105.175 -7.540 -104.175 ;
        RECT -5.080 -105.260 -4.850 -104.260 ;
        RECT -1.390 -105.260 -1.160 -104.260 ;
        RECT -0.410 -105.260 -0.180 -104.260 ;
        RECT 0.570 -105.260 0.800 -104.260 ;
        RECT 1.700 -105.065 1.930 -105.055 ;
        RECT -29.365 -105.760 -28.520 -105.725 ;
        RECT -36.355 -106.575 -36.125 -106.075 ;
        RECT -35.865 -106.575 -35.635 -106.075 ;
        RECT -35.375 -106.575 -35.145 -106.075 ;
        RECT -34.885 -106.575 -34.655 -106.075 ;
        RECT -34.395 -106.575 -34.165 -106.075 ;
        RECT -33.905 -106.575 -33.675 -106.075 ;
        RECT -32.165 -106.550 -31.935 -106.325 ;
        RECT -35.230 -107.160 -34.570 -106.860 ;
        RECT -36.925 -107.640 -36.625 -107.510 ;
        RECT -38.700 -107.955 -36.625 -107.640 ;
        RECT -38.615 -107.960 -36.625 -107.955 ;
        RECT -36.925 -108.195 -36.625 -107.960 ;
        RECT -35.110 -108.250 -34.635 -107.160 ;
        RECT -32.175 -107.320 -31.935 -106.550 ;
        RECT -31.675 -106.825 -31.445 -106.325 ;
        RECT -31.185 -106.730 -30.955 -106.325 ;
        RECT -31.215 -107.320 -30.910 -106.730 ;
        RECT -30.695 -106.825 -30.465 -106.325 ;
        RECT -30.205 -106.720 -29.975 -106.325 ;
        RECT -30.235 -107.320 -29.930 -106.720 ;
        RECT -29.715 -106.825 -29.485 -106.325 ;
        RECT -29.225 -106.730 -28.995 -106.325 ;
        RECT -29.280 -107.320 -28.975 -106.730 ;
        RECT -28.735 -106.825 -28.505 -106.325 ;
        RECT -27.640 -106.575 -27.410 -106.075 ;
        RECT -27.150 -106.575 -26.920 -106.075 ;
        RECT -26.660 -106.575 -26.430 -106.075 ;
        RECT -26.170 -106.575 -25.940 -106.075 ;
        RECT -25.680 -106.575 -25.450 -106.075 ;
        RECT -25.190 -106.575 -24.960 -106.075 ;
        RECT -33.240 -107.660 -32.580 -107.360 ;
        RECT -32.175 -107.560 -24.520 -107.320 ;
        RECT -35.185 -108.550 -34.500 -108.250 ;
        RECT -36.355 -109.865 -36.125 -109.365 ;
        RECT -35.865 -109.865 -35.635 -109.365 ;
        RECT -35.375 -109.865 -35.145 -109.365 ;
        RECT -34.885 -109.865 -34.655 -109.365 ;
        RECT -34.395 -109.865 -34.165 -109.365 ;
        RECT -33.905 -109.865 -33.675 -109.365 ;
        RECT -33.060 -109.995 -32.760 -107.660 ;
        RECT -32.170 -109.865 -31.940 -109.365 ;
        RECT -31.680 -109.865 -31.450 -109.365 ;
        RECT -31.190 -109.865 -30.960 -109.365 ;
        RECT -30.700 -109.865 -30.470 -109.365 ;
        RECT -30.210 -109.865 -29.980 -109.365 ;
        RECT -29.720 -109.865 -29.490 -109.365 ;
        RECT -28.625 -109.615 -28.395 -109.115 ;
        RECT -28.135 -109.615 -27.905 -109.115 ;
        RECT -27.645 -109.615 -27.415 -109.115 ;
        RECT -27.155 -109.615 -26.925 -109.115 ;
        RECT -26.665 -109.615 -26.435 -109.115 ;
        RECT -26.175 -109.615 -25.945 -109.115 ;
        RECT -25.685 -109.615 -25.455 -109.115 ;
        RECT -25.195 -109.615 -24.965 -109.115 ;
        RECT -24.725 -109.985 -24.520 -107.560 ;
        RECT -24.130 -107.805 -23.830 -105.565 ;
        RECT -23.555 -106.125 -23.255 -105.690 ;
        RECT -15.865 -105.725 -10.875 -105.440 ;
        RECT -15.865 -105.760 -15.020 -105.725 ;
        RECT -23.555 -106.350 -23.250 -106.125 ;
        RECT -24.375 -108.105 -23.690 -107.805 ;
        RECT -28.610 -110.215 -27.765 -110.180 ;
        RECT -32.755 -110.500 -27.765 -110.215 ;
        RECT -25.200 -110.285 -24.515 -109.985 ;
        RECT -23.550 -110.090 -23.250 -106.350 ;
        RECT -22.855 -106.575 -22.625 -106.075 ;
        RECT -22.365 -106.575 -22.135 -106.075 ;
        RECT -21.875 -106.575 -21.645 -106.075 ;
        RECT -21.385 -106.575 -21.155 -106.075 ;
        RECT -20.895 -106.575 -20.665 -106.075 ;
        RECT -20.405 -106.575 -20.175 -106.075 ;
        RECT -18.665 -106.825 -18.420 -106.325 ;
        RECT -18.175 -106.825 -17.945 -106.325 ;
        RECT -17.685 -106.825 -17.455 -106.325 ;
        RECT -17.195 -106.825 -16.965 -106.325 ;
        RECT -16.705 -106.825 -16.475 -106.325 ;
        RECT -16.215 -106.825 -15.985 -106.325 ;
        RECT -15.725 -106.825 -15.495 -106.325 ;
        RECT -15.235 -106.825 -15.005 -106.325 ;
        RECT -14.140 -106.575 -13.910 -106.075 ;
        RECT -13.650 -106.575 -13.420 -106.075 ;
        RECT -13.160 -106.575 -12.930 -106.075 ;
        RECT -12.670 -106.575 -12.440 -106.075 ;
        RECT -12.180 -106.575 -11.950 -106.075 ;
        RECT -11.690 -106.575 -11.460 -106.075 ;
        RECT -22.235 -107.180 -21.550 -106.880 ;
        RECT -22.145 -108.220 -21.670 -107.180 ;
        RECT -18.650 -107.310 -18.420 -106.825 ;
        RECT -17.675 -107.310 -17.465 -106.825 ;
        RECT -16.700 -107.310 -16.490 -106.825 ;
        RECT -15.720 -107.310 -15.510 -106.825 ;
        RECT -18.650 -107.540 -14.850 -107.310 ;
        RECT -19.645 -108.100 -18.985 -107.800 ;
        RECT -22.200 -108.520 -21.515 -108.220 ;
        RECT -22.855 -109.865 -22.625 -109.365 ;
        RECT -22.365 -109.865 -22.135 -109.365 ;
        RECT -21.875 -109.865 -21.645 -109.365 ;
        RECT -21.385 -109.865 -21.155 -109.365 ;
        RECT -20.895 -109.865 -20.665 -109.365 ;
        RECT -20.405 -109.865 -20.175 -109.365 ;
        RECT -19.500 -109.920 -19.200 -108.100 ;
        RECT -15.080 -108.370 -14.850 -107.540 ;
        RECT -11.160 -107.910 -10.875 -105.725 ;
        RECT -10.470 -106.230 -10.170 -105.570 ;
        RECT 1.660 -105.735 1.930 -105.065 ;
        RECT 3.585 -105.105 3.815 -104.325 ;
        RECT 4.565 -105.095 4.795 -104.325 ;
        RECT 4.075 -105.105 5.285 -105.095 ;
        RECT 5.545 -105.105 5.775 -104.325 ;
        RECT 3.460 -105.335 5.775 -105.105 ;
        RECT -10.460 -107.370 -10.170 -106.230 ;
        RECT -9.730 -106.575 -9.500 -106.075 ;
        RECT -9.240 -106.575 -9.010 -106.075 ;
        RECT -8.750 -106.575 -8.520 -106.075 ;
        RECT -8.260 -106.575 -8.030 -106.075 ;
        RECT -7.770 -106.575 -7.540 -106.075 ;
        RECT -7.280 -106.575 -7.050 -106.075 ;
        RECT -5.805 -106.555 -5.100 -106.290 ;
        RECT -8.450 -107.175 -7.765 -106.875 ;
        RECT -10.460 -107.660 -9.265 -107.370 ;
        RECT -9.555 -107.805 -9.265 -107.660 ;
        RECT -11.160 -108.195 -9.830 -107.910 ;
        RECT -9.575 -108.105 -8.915 -107.805 ;
        RECT -15.080 -108.375 -11.025 -108.370 ;
        RECT -15.080 -108.600 -10.985 -108.375 ;
        RECT -18.670 -109.865 -18.440 -109.365 ;
        RECT -18.180 -109.865 -17.950 -109.365 ;
        RECT -17.690 -109.865 -17.460 -109.365 ;
        RECT -17.200 -109.865 -16.970 -109.365 ;
        RECT -16.710 -109.865 -16.480 -109.365 ;
        RECT -16.220 -109.865 -15.990 -109.365 ;
        RECT -15.125 -109.615 -14.895 -109.115 ;
        RECT -14.635 -109.615 -14.405 -109.115 ;
        RECT -14.145 -109.615 -13.915 -109.115 ;
        RECT -13.655 -109.615 -13.425 -109.115 ;
        RECT -13.165 -109.615 -12.935 -109.115 ;
        RECT -12.675 -109.615 -12.445 -109.115 ;
        RECT -12.185 -109.615 -11.955 -109.115 ;
        RECT -11.695 -109.615 -11.465 -109.115 ;
        RECT -11.215 -109.975 -10.985 -108.600 ;
        RECT -10.115 -108.800 -9.830 -108.195 ;
        RECT -8.275 -108.220 -7.800 -107.175 ;
        RECT -8.360 -108.520 -7.700 -108.220 ;
        RECT -5.805 -108.800 -5.520 -106.555 ;
        RECT -5.080 -108.800 -4.850 -107.800 ;
        RECT -4.590 -108.800 -4.360 -107.800 ;
        RECT -3.015 -108.800 -2.785 -107.300 ;
        RECT -2.525 -108.800 -2.295 -107.300 ;
        RECT -2.035 -108.800 -1.805 -107.300 ;
        RECT -1.470 -108.800 -1.240 -107.300 ;
        RECT -0.980 -108.800 -0.750 -107.300 ;
        RECT -0.490 -108.800 -0.260 -107.300 ;
        RECT 0.080 -108.795 0.310 -107.295 ;
        RECT 0.570 -108.795 0.800 -107.295 ;
        RECT 1.060 -108.795 1.290 -107.295 ;
        RECT -10.115 -109.085 -5.520 -108.800 ;
        RECT -24.725 -110.290 -24.520 -110.285 ;
        RECT -23.550 -110.390 -22.835 -110.090 ;
        RECT -15.110 -110.215 -14.265 -110.180 ;
        RECT -23.550 -110.420 -23.250 -110.390 ;
        RECT -35.865 -111.765 -35.635 -110.765 ;
        RECT -34.885 -111.765 -34.655 -110.765 ;
        RECT -33.905 -111.765 -33.675 -110.765 ;
        RECT -32.755 -111.675 -32.470 -110.500 ;
        RECT -28.610 -110.550 -27.765 -110.500 ;
        RECT -19.255 -110.500 -14.265 -110.215 ;
        RECT -11.755 -110.275 -10.985 -109.975 ;
        RECT 1.660 -109.760 1.890 -105.735 ;
        RECT 2.105 -106.155 2.785 -105.925 ;
        RECT 4.075 -105.980 4.305 -105.335 ;
        RECT 4.565 -105.980 4.795 -105.480 ;
        RECT 5.055 -105.980 5.285 -105.335 ;
        RECT 5.545 -105.980 5.775 -105.480 ;
        RECT 2.425 -109.200 2.655 -106.155 ;
        RECT 7.120 -108.695 7.350 -107.015 ;
        RECT 7.610 -108.515 7.840 -104.330 ;
        RECT 8.590 -105.830 8.820 -104.330 ;
        RECT 11.610 -105.115 11.840 -104.335 ;
        RECT 12.590 -105.105 12.820 -104.335 ;
        RECT 12.100 -105.115 13.310 -105.105 ;
        RECT 13.570 -105.115 13.800 -104.335 ;
        RECT 11.485 -105.345 13.800 -105.115 ;
        RECT 12.100 -105.990 12.330 -105.345 ;
        RECT 12.590 -105.990 12.820 -105.490 ;
        RECT 13.080 -105.990 13.310 -105.345 ;
        RECT 13.570 -105.990 13.800 -105.490 ;
        RECT 8.100 -108.695 8.330 -107.015 ;
        RECT 8.590 -108.515 8.820 -107.015 ;
        RECT 9.080 -108.510 9.310 -107.015 ;
        RECT 9.080 -108.695 9.315 -108.510 ;
        RECT 7.120 -108.930 9.315 -108.695 ;
        RECT 15.145 -108.705 15.375 -107.025 ;
        RECT 15.635 -108.525 15.865 -104.340 ;
        RECT 16.615 -105.840 16.845 -104.340 ;
        RECT 19.730 -105.215 19.960 -104.215 ;
        RECT 23.420 -105.215 23.650 -104.215 ;
        RECT 24.400 -105.215 24.630 -104.215 ;
        RECT 25.380 -105.215 25.610 -104.215 ;
        RECT 27.795 -105.270 28.025 -104.270 ;
        RECT 28.285 -105.425 28.515 -104.270 ;
        RECT 28.775 -105.270 29.005 -104.270 ;
        RECT 29.375 -105.270 29.605 -104.270 ;
        RECT 29.865 -105.270 30.095 -104.270 ;
        RECT 30.355 -105.270 30.585 -104.270 ;
        RECT 32.165 -105.270 32.395 -104.270 ;
        RECT 33.145 -105.270 33.375 -104.270 ;
        RECT 34.695 -105.270 34.925 -104.270 ;
        RECT 36.240 -105.270 36.470 -104.270 ;
        RECT 25.755 -105.655 28.515 -105.425 ;
        RECT 25.775 -105.700 26.455 -105.655 ;
        RECT 33.610 -105.910 34.305 -105.820 ;
        RECT 36.685 -105.875 37.380 -105.850 ;
        RECT 41.340 -105.875 42.430 -105.580 ;
        RECT 36.685 -105.910 42.430 -105.875 ;
        RECT 33.610 -106.015 42.430 -105.910 ;
        RECT 27.820 -106.105 28.515 -106.040 ;
        RECT 33.610 -106.050 37.885 -106.015 ;
        RECT 41.340 -106.025 42.430 -106.015 ;
        RECT 33.610 -106.090 34.305 -106.050 ;
        RECT 27.820 -106.245 29.590 -106.105 ;
        RECT 36.685 -106.120 37.380 -106.050 ;
        RECT 27.820 -106.310 28.515 -106.245 ;
        RECT 29.450 -106.970 29.590 -106.245 ;
        RECT 31.565 -106.235 32.260 -106.190 ;
        RECT 35.750 -106.235 36.430 -106.190 ;
        RECT 31.565 -106.375 36.430 -106.235 ;
        RECT 31.565 -106.460 32.260 -106.375 ;
        RECT 35.750 -106.420 36.430 -106.375 ;
        RECT 34.220 -106.970 34.875 -106.910 ;
        RECT 16.125 -108.705 16.355 -107.025 ;
        RECT 16.615 -108.525 16.845 -107.025 ;
        RECT 17.105 -108.520 17.335 -107.025 ;
        RECT 29.450 -107.110 34.875 -106.970 ;
        RECT 34.220 -107.140 34.875 -107.110 ;
        RECT 17.105 -108.705 17.340 -108.520 ;
        RECT 15.145 -108.940 17.340 -108.705 ;
        RECT 19.730 -108.755 19.960 -107.755 ;
        RECT 20.220 -108.755 20.450 -107.755 ;
        RECT 21.795 -108.755 22.025 -107.255 ;
        RECT 22.285 -108.755 22.515 -107.255 ;
        RECT 22.775 -108.755 23.005 -107.255 ;
        RECT 23.340 -108.755 23.570 -107.255 ;
        RECT 23.830 -108.755 24.060 -107.255 ;
        RECT 24.320 -108.755 24.550 -107.255 ;
        RECT 24.890 -108.750 25.120 -107.250 ;
        RECT 25.380 -108.750 25.610 -107.250 ;
        RECT 25.870 -108.750 26.100 -107.250 ;
        RECT 27.795 -108.300 28.025 -107.300 ;
        RECT 28.285 -108.300 28.515 -107.300 ;
        RECT 29.865 -108.300 30.095 -107.300 ;
        RECT 30.355 -108.300 30.585 -107.300 ;
        RECT 31.675 -108.300 31.905 -107.300 ;
        RECT 32.165 -108.300 32.395 -107.300 ;
        RECT 33.145 -108.300 33.375 -107.300 ;
        RECT 33.635 -108.300 33.865 -107.300 ;
        RECT 34.695 -108.300 34.925 -107.300 ;
        RECT 35.185 -108.300 35.415 -107.300 ;
        RECT 36.240 -108.300 36.470 -107.300 ;
        RECT 36.730 -108.300 36.960 -107.300 ;
        RECT 2.425 -109.430 11.170 -109.200 ;
        RECT 1.660 -109.990 19.010 -109.760 ;
        RECT -31.680 -111.765 -31.450 -110.765 ;
        RECT -30.700 -111.765 -30.470 -110.765 ;
        RECT -29.720 -111.765 -29.490 -110.765 ;
        RECT -28.625 -111.690 -28.395 -111.190 ;
        RECT -28.135 -111.690 -27.905 -111.190 ;
        RECT -27.645 -111.690 -27.415 -111.190 ;
        RECT -27.155 -111.690 -26.925 -111.190 ;
        RECT -26.665 -111.690 -26.435 -111.190 ;
        RECT -26.175 -111.690 -25.945 -111.190 ;
        RECT -25.685 -111.690 -25.455 -111.190 ;
        RECT -25.195 -111.690 -24.965 -111.190 ;
        RECT -22.365 -111.765 -22.135 -110.765 ;
        RECT -21.385 -111.765 -21.155 -110.765 ;
        RECT -20.405 -111.765 -20.175 -110.765 ;
        RECT -19.255 -111.675 -18.970 -110.500 ;
        RECT -15.110 -110.550 -14.265 -110.500 ;
        RECT -18.180 -111.765 -17.950 -110.765 ;
        RECT -17.200 -111.765 -16.970 -110.765 ;
        RECT -16.220 -111.765 -15.990 -110.765 ;
        RECT -15.125 -111.690 -14.895 -111.190 ;
        RECT -14.635 -111.690 -14.405 -111.190 ;
        RECT -14.145 -111.690 -13.915 -111.190 ;
        RECT -13.655 -111.690 -13.425 -111.190 ;
        RECT -13.165 -111.690 -12.935 -111.190 ;
        RECT -12.675 -111.690 -12.445 -111.190 ;
        RECT -12.185 -111.690 -11.955 -111.190 ;
        RECT -11.695 -111.690 -11.465 -111.190 ;
        RECT -35.865 -118.955 -35.635 -117.955 ;
        RECT -34.885 -118.955 -34.655 -117.955 ;
        RECT -33.905 -118.955 -33.675 -117.955 ;
        RECT -32.755 -119.220 -32.470 -118.045 ;
        RECT -31.680 -118.955 -31.450 -117.955 ;
        RECT -30.700 -118.955 -30.470 -117.955 ;
        RECT -29.720 -118.955 -29.490 -117.955 ;
        RECT -28.625 -118.530 -28.395 -118.030 ;
        RECT -28.135 -118.530 -27.905 -118.030 ;
        RECT -27.645 -118.530 -27.415 -118.030 ;
        RECT -27.155 -118.530 -26.925 -118.030 ;
        RECT -26.665 -118.530 -26.435 -118.030 ;
        RECT -26.175 -118.530 -25.945 -118.030 ;
        RECT -25.685 -118.530 -25.455 -118.030 ;
        RECT -25.195 -118.530 -24.965 -118.030 ;
        RECT -22.365 -118.955 -22.135 -117.955 ;
        RECT -21.385 -118.955 -21.155 -117.955 ;
        RECT -20.405 -118.955 -20.175 -117.955 ;
        RECT -28.610 -119.220 -27.765 -119.170 ;
        RECT -32.755 -119.505 -27.765 -119.220 ;
        RECT -19.255 -119.220 -18.970 -118.045 ;
        RECT -18.180 -118.955 -17.950 -117.955 ;
        RECT -17.200 -118.955 -16.970 -117.955 ;
        RECT -16.220 -118.955 -15.990 -117.955 ;
        RECT -15.125 -118.530 -14.895 -118.030 ;
        RECT -14.635 -118.530 -14.405 -118.030 ;
        RECT -14.145 -118.530 -13.915 -118.030 ;
        RECT -13.655 -118.530 -13.425 -118.030 ;
        RECT -13.165 -118.530 -12.935 -118.030 ;
        RECT -12.675 -118.530 -12.445 -118.030 ;
        RECT -12.185 -118.530 -11.955 -118.030 ;
        RECT -11.695 -118.530 -11.465 -118.030 ;
        RECT -15.110 -119.220 -14.265 -119.170 ;
        RECT -23.550 -119.330 -23.250 -119.300 ;
        RECT -24.725 -119.435 -24.520 -119.430 ;
        RECT -28.610 -119.540 -27.765 -119.505 ;
        RECT -36.355 -120.355 -36.125 -119.855 ;
        RECT -35.865 -120.355 -35.635 -119.855 ;
        RECT -35.375 -120.355 -35.145 -119.855 ;
        RECT -34.885 -120.355 -34.655 -119.855 ;
        RECT -34.395 -120.355 -34.165 -119.855 ;
        RECT -33.905 -120.355 -33.675 -119.855 ;
        RECT -38.655 -121.760 -37.780 -120.665 ;
        RECT -35.185 -121.470 -34.500 -121.170 ;
        RECT -36.925 -121.760 -36.625 -121.525 ;
        RECT -38.655 -122.080 -36.625 -121.760 ;
        RECT -38.655 -122.235 -37.780 -122.080 ;
        RECT -36.925 -122.210 -36.625 -122.080 ;
        RECT -35.110 -122.410 -34.635 -121.470 ;
        RECT -33.060 -122.060 -32.760 -119.725 ;
        RECT -25.200 -119.735 -24.515 -119.435 ;
        RECT -23.550 -119.630 -22.835 -119.330 ;
        RECT -19.255 -119.505 -14.265 -119.220 ;
        RECT -15.110 -119.540 -14.265 -119.505 ;
        RECT -32.170 -120.355 -31.940 -119.855 ;
        RECT -31.680 -120.355 -31.450 -119.855 ;
        RECT -31.190 -120.355 -30.960 -119.855 ;
        RECT -30.700 -120.355 -30.470 -119.855 ;
        RECT -30.210 -120.355 -29.980 -119.855 ;
        RECT -29.720 -120.355 -29.490 -119.855 ;
        RECT -28.625 -120.605 -28.395 -120.105 ;
        RECT -28.135 -120.605 -27.905 -120.105 ;
        RECT -27.645 -120.605 -27.415 -120.105 ;
        RECT -27.155 -120.605 -26.925 -120.105 ;
        RECT -26.665 -120.605 -26.435 -120.105 ;
        RECT -26.175 -120.605 -25.945 -120.105 ;
        RECT -25.685 -120.605 -25.455 -120.105 ;
        RECT -25.195 -120.605 -24.965 -120.105 ;
        RECT -33.240 -122.360 -32.580 -122.060 ;
        RECT -24.725 -122.160 -24.520 -119.735 ;
        RECT -24.375 -121.915 -23.690 -121.615 ;
        RECT -37.545 -122.560 -34.635 -122.410 ;
        RECT -32.175 -122.400 -24.520 -122.160 ;
        RECT -37.545 -122.860 -34.570 -122.560 ;
        RECT -37.545 -122.885 -34.635 -122.860 ;
        RECT -37.545 -123.280 -37.070 -122.885 ;
        RECT -38.620 -123.755 -37.070 -123.280 ;
        RECT -36.355 -123.645 -36.125 -123.145 ;
        RECT -35.865 -123.645 -35.635 -123.145 ;
        RECT -35.375 -123.645 -35.145 -123.145 ;
        RECT -34.885 -123.645 -34.655 -123.145 ;
        RECT -34.395 -123.645 -34.165 -123.145 ;
        RECT -33.905 -123.645 -33.675 -123.145 ;
        RECT -32.175 -123.170 -31.935 -122.400 ;
        RECT -32.165 -123.395 -31.935 -123.170 ;
        RECT -31.675 -123.395 -31.445 -122.895 ;
        RECT -31.215 -122.990 -30.910 -122.400 ;
        RECT -31.185 -123.395 -30.955 -122.990 ;
        RECT -30.695 -123.395 -30.465 -122.895 ;
        RECT -30.235 -123.000 -29.930 -122.400 ;
        RECT -30.205 -123.395 -29.975 -123.000 ;
        RECT -29.715 -123.395 -29.485 -122.895 ;
        RECT -29.280 -122.990 -28.975 -122.400 ;
        RECT -29.225 -123.395 -28.995 -122.990 ;
        RECT -28.735 -123.395 -28.505 -122.895 ;
        RECT -27.640 -123.645 -27.410 -123.145 ;
        RECT -27.150 -123.645 -26.920 -123.145 ;
        RECT -26.660 -123.645 -26.430 -123.145 ;
        RECT -26.170 -123.645 -25.940 -123.145 ;
        RECT -25.680 -123.645 -25.450 -123.145 ;
        RECT -25.190 -123.645 -24.960 -123.145 ;
        RECT -29.365 -123.995 -28.520 -123.960 ;
        RECT -29.365 -124.280 -24.375 -123.995 ;
        RECT -24.130 -124.155 -23.830 -121.915 ;
        RECT -23.550 -123.370 -23.250 -119.630 ;
        RECT -11.755 -119.745 -10.985 -119.445 ;
        RECT -22.855 -120.355 -22.625 -119.855 ;
        RECT -22.365 -120.355 -22.135 -119.855 ;
        RECT -21.875 -120.355 -21.645 -119.855 ;
        RECT -21.385 -120.355 -21.155 -119.855 ;
        RECT -20.895 -120.355 -20.665 -119.855 ;
        RECT -20.405 -120.355 -20.175 -119.855 ;
        RECT -22.200 -121.500 -21.515 -121.200 ;
        RECT -22.145 -122.540 -21.670 -121.500 ;
        RECT -19.500 -121.620 -19.200 -119.800 ;
        RECT -18.670 -120.355 -18.440 -119.855 ;
        RECT -18.180 -120.355 -17.950 -119.855 ;
        RECT -17.690 -120.355 -17.460 -119.855 ;
        RECT -17.200 -120.355 -16.970 -119.855 ;
        RECT -16.710 -120.355 -16.480 -119.855 ;
        RECT -16.220 -120.355 -15.990 -119.855 ;
        RECT -15.125 -120.605 -14.895 -120.105 ;
        RECT -14.635 -120.605 -14.405 -120.105 ;
        RECT -14.145 -120.605 -13.915 -120.105 ;
        RECT -13.655 -120.605 -13.425 -120.105 ;
        RECT -13.165 -120.605 -12.935 -120.105 ;
        RECT -12.675 -120.605 -12.445 -120.105 ;
        RECT -12.185 -120.605 -11.955 -120.105 ;
        RECT -11.695 -120.605 -11.465 -120.105 ;
        RECT -11.215 -121.120 -10.985 -119.745 ;
        RECT 1.660 -119.960 19.010 -119.730 ;
        RECT -15.080 -121.345 -10.985 -121.120 ;
        RECT -10.115 -120.920 -5.520 -120.635 ;
        RECT -15.080 -121.350 -11.025 -121.345 ;
        RECT -19.645 -121.920 -18.985 -121.620 ;
        RECT -15.080 -122.180 -14.850 -121.350 ;
        RECT -10.115 -121.525 -9.830 -120.920 ;
        RECT -9.010 -121.500 -8.350 -121.200 ;
        RECT -18.650 -122.410 -14.850 -122.180 ;
        RECT -11.160 -121.810 -9.830 -121.525 ;
        RECT -22.235 -122.840 -21.550 -122.540 ;
        RECT -18.650 -122.895 -18.420 -122.410 ;
        RECT -17.675 -122.895 -17.465 -122.410 ;
        RECT -16.700 -122.895 -16.490 -122.410 ;
        RECT -15.720 -122.895 -15.510 -122.410 ;
        RECT -23.555 -123.595 -23.250 -123.370 ;
        RECT -23.555 -124.030 -23.255 -123.595 ;
        RECT -22.855 -123.645 -22.625 -123.145 ;
        RECT -22.365 -123.645 -22.135 -123.145 ;
        RECT -21.875 -123.645 -21.645 -123.145 ;
        RECT -21.385 -123.645 -21.155 -123.145 ;
        RECT -20.895 -123.645 -20.665 -123.145 ;
        RECT -20.405 -123.645 -20.175 -123.145 ;
        RECT -18.665 -123.395 -18.420 -122.895 ;
        RECT -18.175 -123.395 -17.945 -122.895 ;
        RECT -17.685 -123.395 -17.455 -122.895 ;
        RECT -17.195 -123.395 -16.965 -122.895 ;
        RECT -16.705 -123.395 -16.475 -122.895 ;
        RECT -16.215 -123.395 -15.985 -122.895 ;
        RECT -15.725 -123.395 -15.495 -122.895 ;
        RECT -15.235 -123.395 -15.005 -122.895 ;
        RECT -14.140 -123.645 -13.910 -123.145 ;
        RECT -13.650 -123.645 -13.420 -123.145 ;
        RECT -13.160 -123.645 -12.930 -123.145 ;
        RECT -12.670 -123.645 -12.440 -123.145 ;
        RECT -12.180 -123.645 -11.950 -123.145 ;
        RECT -11.690 -123.645 -11.460 -123.145 ;
        RECT -15.865 -123.995 -15.020 -123.960 ;
        RECT -11.160 -123.995 -10.875 -121.810 ;
        RECT -10.625 -122.350 -9.965 -122.050 ;
        RECT -10.460 -123.490 -10.170 -122.350 ;
        RECT -8.925 -122.545 -8.450 -121.500 ;
        RECT -9.100 -122.845 -8.415 -122.545 ;
        RECT -29.365 -124.330 -28.520 -124.280 ;
        RECT -36.355 -125.545 -36.125 -124.545 ;
        RECT -35.375 -125.545 -35.145 -124.545 ;
        RECT -34.395 -125.545 -34.165 -124.545 ;
        RECT -32.165 -125.470 -31.935 -124.970 ;
        RECT -31.675 -125.470 -31.445 -124.970 ;
        RECT -31.185 -125.470 -30.955 -124.970 ;
        RECT -30.695 -125.470 -30.465 -124.970 ;
        RECT -30.205 -125.470 -29.975 -124.970 ;
        RECT -29.715 -125.470 -29.485 -124.970 ;
        RECT -29.225 -125.470 -28.995 -124.970 ;
        RECT -28.735 -125.470 -28.505 -124.970 ;
        RECT -27.640 -125.545 -27.410 -124.545 ;
        RECT -26.660 -125.545 -26.430 -124.545 ;
        RECT -25.680 -125.545 -25.450 -124.545 ;
        RECT -24.660 -125.455 -24.375 -124.280 ;
        RECT -15.865 -124.280 -10.875 -123.995 ;
        RECT -10.470 -124.150 -10.170 -123.490 ;
        RECT -9.730 -123.645 -9.500 -123.145 ;
        RECT -9.240 -123.645 -9.010 -123.145 ;
        RECT -8.750 -123.645 -8.520 -123.145 ;
        RECT -8.260 -123.645 -8.030 -123.145 ;
        RECT -7.770 -123.645 -7.540 -123.145 ;
        RECT -7.280 -123.645 -7.050 -123.145 ;
        RECT -5.805 -123.165 -5.520 -120.920 ;
        RECT -5.080 -121.920 -4.850 -120.920 ;
        RECT -4.590 -121.920 -4.360 -120.920 ;
        RECT -3.015 -122.420 -2.785 -120.920 ;
        RECT -2.525 -122.420 -2.295 -120.920 ;
        RECT -2.035 -122.420 -1.805 -120.920 ;
        RECT -1.470 -122.420 -1.240 -120.920 ;
        RECT -0.980 -122.420 -0.750 -120.920 ;
        RECT -0.490 -122.420 -0.260 -120.920 ;
        RECT 0.080 -122.425 0.310 -120.925 ;
        RECT 0.570 -122.425 0.800 -120.925 ;
        RECT 1.060 -122.425 1.290 -120.925 ;
        RECT -5.805 -123.430 -5.100 -123.165 ;
        RECT 1.660 -123.985 1.890 -119.960 ;
        RECT 2.425 -120.520 11.170 -120.290 ;
        RECT 2.425 -123.565 2.655 -120.520 ;
        RECT 7.120 -121.025 9.315 -120.790 ;
        RECT 7.120 -122.705 7.350 -121.025 ;
        RECT 2.105 -123.795 2.785 -123.565 ;
        RECT -15.865 -124.330 -15.020 -124.280 ;
        RECT -22.855 -125.545 -22.625 -124.545 ;
        RECT -21.875 -125.545 -21.645 -124.545 ;
        RECT -20.895 -125.545 -20.665 -124.545 ;
        RECT -18.665 -125.470 -18.435 -124.970 ;
        RECT -18.175 -125.470 -17.945 -124.970 ;
        RECT -17.685 -125.470 -17.455 -124.970 ;
        RECT -17.195 -125.470 -16.965 -124.970 ;
        RECT -16.705 -125.470 -16.475 -124.970 ;
        RECT -16.215 -125.470 -15.985 -124.970 ;
        RECT -15.725 -125.470 -15.495 -124.970 ;
        RECT -15.235 -125.470 -15.005 -124.970 ;
        RECT -14.140 -125.545 -13.910 -124.545 ;
        RECT -13.160 -125.545 -12.930 -124.545 ;
        RECT -12.180 -125.545 -11.950 -124.545 ;
        RECT -11.160 -125.455 -10.875 -124.280 ;
        RECT -9.730 -125.545 -9.500 -124.545 ;
        RECT -8.750 -125.545 -8.520 -124.545 ;
        RECT -7.770 -125.545 -7.540 -124.545 ;
        RECT -5.080 -125.460 -4.850 -124.460 ;
        RECT -1.390 -125.460 -1.160 -124.460 ;
        RECT -0.410 -125.460 -0.180 -124.460 ;
        RECT 0.570 -125.460 0.800 -124.460 ;
        RECT 1.660 -124.655 1.930 -123.985 ;
        RECT 4.075 -124.385 4.305 -123.740 ;
        RECT 4.565 -124.240 4.795 -123.740 ;
        RECT 5.055 -124.385 5.285 -123.740 ;
        RECT 5.545 -124.240 5.775 -123.740 ;
        RECT 3.460 -124.615 5.775 -124.385 ;
        RECT 1.700 -124.665 1.930 -124.655 ;
        RECT 3.585 -125.395 3.815 -124.615 ;
        RECT 4.075 -124.625 5.285 -124.615 ;
        RECT 4.565 -125.395 4.795 -124.625 ;
        RECT 5.545 -125.395 5.775 -124.615 ;
        RECT 7.610 -125.390 7.840 -121.205 ;
        RECT 8.100 -122.705 8.330 -121.025 ;
        RECT 8.590 -122.705 8.820 -121.205 ;
        RECT 9.080 -121.210 9.315 -121.025 ;
        RECT 15.145 -121.015 17.340 -120.780 ;
        RECT 9.080 -122.705 9.310 -121.210 ;
        RECT 15.145 -122.695 15.375 -121.015 ;
        RECT 8.590 -125.390 8.820 -123.890 ;
        RECT 12.100 -124.375 12.330 -123.730 ;
        RECT 12.590 -124.230 12.820 -123.730 ;
        RECT 13.080 -124.375 13.310 -123.730 ;
        RECT 13.570 -124.230 13.800 -123.730 ;
        RECT 11.485 -124.605 13.800 -124.375 ;
        RECT 11.610 -125.385 11.840 -124.605 ;
        RECT 12.100 -124.615 13.310 -124.605 ;
        RECT 12.590 -125.385 12.820 -124.615 ;
        RECT 13.570 -125.385 13.800 -124.605 ;
        RECT 15.635 -125.380 15.865 -121.195 ;
        RECT 16.125 -122.695 16.355 -121.015 ;
        RECT 16.615 -122.695 16.845 -121.195 ;
        RECT 17.105 -121.200 17.340 -121.015 ;
        RECT 17.105 -122.695 17.335 -121.200 ;
        RECT 19.730 -121.965 19.960 -120.965 ;
        RECT 20.220 -121.965 20.450 -120.965 ;
        RECT 21.795 -122.465 22.025 -120.965 ;
        RECT 22.285 -122.465 22.515 -120.965 ;
        RECT 22.775 -122.465 23.005 -120.965 ;
        RECT 23.340 -122.465 23.570 -120.965 ;
        RECT 23.830 -122.465 24.060 -120.965 ;
        RECT 24.320 -122.465 24.550 -120.965 ;
        RECT 24.890 -122.470 25.120 -120.970 ;
        RECT 25.380 -122.470 25.610 -120.970 ;
        RECT 25.870 -122.470 26.100 -120.970 ;
        RECT 27.795 -122.420 28.025 -121.420 ;
        RECT 28.285 -122.420 28.515 -121.420 ;
        RECT 29.865 -122.420 30.095 -121.420 ;
        RECT 30.355 -122.420 30.585 -121.420 ;
        RECT 31.675 -122.420 31.905 -121.420 ;
        RECT 32.165 -122.420 32.395 -121.420 ;
        RECT 33.145 -122.420 33.375 -121.420 ;
        RECT 33.635 -122.420 33.865 -121.420 ;
        RECT 34.695 -122.420 34.925 -121.420 ;
        RECT 35.185 -122.420 35.415 -121.420 ;
        RECT 36.240 -122.420 36.470 -121.420 ;
        RECT 36.730 -122.420 36.960 -121.420 ;
        RECT 34.220 -122.610 34.875 -122.580 ;
        RECT 29.450 -122.750 34.875 -122.610 ;
        RECT 27.820 -123.475 28.515 -123.410 ;
        RECT 29.450 -123.475 29.590 -122.750 ;
        RECT 34.220 -122.810 34.875 -122.750 ;
        RECT 27.820 -123.615 29.590 -123.475 ;
        RECT 31.565 -123.345 32.260 -123.260 ;
        RECT 35.750 -123.345 36.430 -123.300 ;
        RECT 31.565 -123.485 36.430 -123.345 ;
        RECT 31.565 -123.530 32.260 -123.485 ;
        RECT 35.750 -123.530 36.430 -123.485 ;
        RECT 27.820 -123.680 28.515 -123.615 ;
        RECT 33.610 -123.670 34.305 -123.630 ;
        RECT 36.685 -123.670 37.380 -123.600 ;
        RECT 33.610 -123.705 37.885 -123.670 ;
        RECT 42.175 -123.705 42.315 -106.025 ;
        RECT 33.610 -123.810 42.315 -123.705 ;
        RECT 16.615 -125.380 16.845 -123.880 ;
        RECT 33.610 -123.900 34.305 -123.810 ;
        RECT 36.685 -123.845 42.315 -123.810 ;
        RECT 36.685 -123.870 37.380 -123.845 ;
        RECT 25.775 -124.065 26.455 -124.020 ;
        RECT 25.755 -124.295 28.515 -124.065 ;
        RECT 19.730 -125.505 19.960 -124.505 ;
        RECT 23.420 -125.505 23.650 -124.505 ;
        RECT 24.400 -125.505 24.630 -124.505 ;
        RECT 25.380 -125.505 25.610 -124.505 ;
        RECT 27.795 -125.450 28.025 -124.450 ;
        RECT 28.285 -125.450 28.515 -124.295 ;
        RECT 28.775 -125.450 29.005 -124.450 ;
        RECT 29.375 -125.450 29.605 -124.450 ;
        RECT 29.865 -125.450 30.095 -124.450 ;
        RECT 30.355 -125.450 30.585 -124.450 ;
        RECT 32.165 -125.450 32.395 -124.450 ;
        RECT 33.145 -125.450 33.375 -124.450 ;
        RECT 34.695 -125.450 34.925 -124.450 ;
        RECT 36.240 -125.450 36.470 -124.450 ;
        RECT 42.745 -126.950 43.000 -102.770 ;
        RECT 43.850 -119.480 44.105 -101.090 ;
        RECT 43.835 -119.955 44.130 -119.480 ;
        RECT -6.815 -127.205 43.000 -126.950 ;
        RECT 9.145 -127.415 9.920 -127.405 ;
        RECT -37.360 -127.450 9.920 -127.415 ;
        RECT -37.980 -127.625 9.920 -127.450 ;
        RECT 42.745 -127.560 43.000 -127.205 ;
        RECT -37.980 -127.680 -37.300 -127.625 ;
        RECT 9.145 -127.635 9.920 -127.625 ;
        RECT -25.580 -127.825 -24.900 -127.815 ;
        RECT -25.580 -128.035 10.345 -127.825 ;
        RECT -25.580 -128.045 -24.900 -128.035 ;
        RECT 9.665 -128.055 10.345 -128.035 ;
        RECT 42.145 -128.095 43.100 -127.560 ;
        RECT 43.850 -128.630 44.105 -119.955 ;
        RECT 44.630 -123.440 44.885 -100.340 ;
        RECT 45.540 -117.880 45.680 -99.660 ;
        RECT 46.250 -106.695 46.440 -99.025 ;
        RECT 46.250 -107.360 46.500 -106.695 ;
        RECT 45.440 -118.470 45.760 -117.880 ;
        RECT 44.600 -124.135 44.945 -123.440 ;
        RECT -27.055 -128.860 44.105 -128.630 ;
        RECT -27.055 -128.885 41.985 -128.860 ;
        RECT -37.255 -133.675 -37.025 -132.675 ;
        RECT -36.765 -133.675 -36.535 -132.675 ;
        RECT -35.185 -133.675 -34.955 -132.675 ;
        RECT -34.695 -133.675 -34.465 -132.675 ;
        RECT -33.375 -133.675 -33.145 -132.675 ;
        RECT -32.885 -133.675 -32.655 -132.675 ;
        RECT -31.905 -133.675 -31.675 -132.675 ;
        RECT -31.415 -133.675 -31.185 -132.675 ;
        RECT -30.355 -133.675 -30.125 -132.675 ;
        RECT -29.865 -133.675 -29.635 -132.675 ;
        RECT -28.810 -133.675 -28.580 -132.675 ;
        RECT -28.320 -133.675 -28.090 -132.675 ;
        RECT -30.830 -133.865 -30.175 -133.835 ;
        RECT -35.600 -134.005 -30.175 -133.865 ;
        RECT -37.230 -134.730 -36.535 -134.665 ;
        RECT -35.600 -134.730 -35.460 -134.005 ;
        RECT -30.830 -134.065 -30.175 -134.005 ;
        RECT -37.230 -134.870 -35.460 -134.730 ;
        RECT -33.485 -134.600 -32.790 -134.515 ;
        RECT -29.300 -134.600 -28.620 -134.555 ;
        RECT -33.485 -134.740 -28.620 -134.600 ;
        RECT -33.485 -134.785 -32.790 -134.740 ;
        RECT -29.300 -134.785 -28.620 -134.740 ;
        RECT -37.230 -134.935 -36.535 -134.870 ;
        RECT -31.440 -134.925 -30.745 -134.885 ;
        RECT -28.365 -134.925 -27.670 -134.855 ;
        RECT -27.055 -134.925 -26.915 -128.885 ;
        RECT -25.595 -129.990 -25.365 -129.310 ;
        RECT 44.630 -129.380 44.885 -124.135 ;
        RECT -14.200 -129.535 44.885 -129.380 ;
        RECT -14.200 -129.635 41.985 -129.535 ;
        RECT 42.950 -129.570 44.885 -129.535 ;
        RECT -25.590 -132.840 -25.370 -129.990 ;
        RECT -25.595 -133.520 -25.365 -132.840 ;
        RECT -24.755 -133.675 -24.525 -132.675 ;
        RECT -24.265 -133.675 -24.035 -132.675 ;
        RECT -22.685 -133.675 -22.455 -132.675 ;
        RECT -22.195 -133.675 -21.965 -132.675 ;
        RECT -20.875 -133.675 -20.645 -132.675 ;
        RECT -20.385 -133.675 -20.155 -132.675 ;
        RECT -19.405 -133.675 -19.175 -132.675 ;
        RECT -18.915 -133.675 -18.685 -132.675 ;
        RECT -17.855 -133.675 -17.625 -132.675 ;
        RECT -17.365 -133.675 -17.135 -132.675 ;
        RECT -16.310 -133.675 -16.080 -132.675 ;
        RECT -15.820 -133.675 -15.590 -132.675 ;
        RECT -18.330 -133.865 -17.675 -133.835 ;
        RECT -23.100 -134.005 -17.675 -133.865 ;
        RECT -31.440 -135.065 -26.915 -134.925 ;
        RECT -24.730 -134.730 -24.035 -134.665 ;
        RECT -23.100 -134.730 -22.960 -134.005 ;
        RECT -18.330 -134.065 -17.675 -134.005 ;
        RECT -24.730 -134.870 -22.960 -134.730 ;
        RECT -20.985 -134.600 -20.290 -134.515 ;
        RECT -16.800 -134.600 -16.120 -134.555 ;
        RECT -20.985 -134.740 -16.120 -134.600 ;
        RECT -20.985 -134.785 -20.290 -134.740 ;
        RECT -16.800 -134.785 -16.120 -134.740 ;
        RECT -24.730 -134.935 -24.035 -134.870 ;
        RECT -18.940 -134.925 -18.245 -134.885 ;
        RECT -15.865 -134.925 -15.170 -134.855 ;
        RECT -14.200 -134.925 -14.060 -129.635 ;
        RECT 45.540 -130.060 45.680 -118.470 ;
        RECT -1.840 -130.200 45.680 -130.060 ;
        RECT -12.030 -131.415 -11.350 -131.410 ;
        RECT -12.855 -131.635 -11.350 -131.415 ;
        RECT -12.850 -132.820 -12.630 -131.635 ;
        RECT -12.030 -131.640 -11.350 -131.635 ;
        RECT -12.855 -133.500 -12.625 -132.820 ;
        RECT -12.255 -133.675 -12.025 -132.675 ;
        RECT -11.765 -133.675 -11.535 -132.675 ;
        RECT -10.185 -133.675 -9.955 -132.675 ;
        RECT -9.695 -133.675 -9.465 -132.675 ;
        RECT -8.375 -133.675 -8.145 -132.675 ;
        RECT -7.885 -133.675 -7.655 -132.675 ;
        RECT -6.905 -133.675 -6.675 -132.675 ;
        RECT -6.415 -133.675 -6.185 -132.675 ;
        RECT -5.355 -133.675 -5.125 -132.675 ;
        RECT -4.865 -133.675 -4.635 -132.675 ;
        RECT -3.810 -133.675 -3.580 -132.675 ;
        RECT -3.320 -133.675 -3.090 -132.675 ;
        RECT -5.830 -133.865 -5.175 -133.835 ;
        RECT -10.600 -134.005 -5.175 -133.865 ;
        RECT -18.940 -135.065 -14.060 -134.925 ;
        RECT -12.230 -134.730 -11.535 -134.665 ;
        RECT -10.600 -134.730 -10.460 -134.005 ;
        RECT -5.830 -134.065 -5.175 -134.005 ;
        RECT -12.230 -134.870 -10.460 -134.730 ;
        RECT -8.485 -134.600 -7.790 -134.515 ;
        RECT -4.300 -134.600 -3.620 -134.555 ;
        RECT -8.485 -134.740 -3.620 -134.600 ;
        RECT -8.485 -134.785 -7.790 -134.740 ;
        RECT -4.300 -134.785 -3.620 -134.740 ;
        RECT -12.230 -134.935 -11.535 -134.870 ;
        RECT -6.440 -134.925 -5.745 -134.885 ;
        RECT -3.365 -134.925 -2.670 -134.855 ;
        RECT -1.840 -134.925 -1.700 -130.200 ;
        RECT 46.250 -130.695 46.440 -107.360 ;
        RECT 10.535 -130.745 39.025 -130.695 ;
        RECT 42.425 -130.745 46.440 -130.695 ;
        RECT 10.535 -130.885 46.440 -130.745 ;
        RECT 0.455 -131.350 1.135 -131.345 ;
        RECT -0.450 -131.570 1.135 -131.350 ;
        RECT -0.450 -132.820 -0.230 -131.570 ;
        RECT 0.455 -131.575 1.135 -131.570 ;
        RECT -0.455 -133.500 -0.225 -132.820 ;
        RECT 0.245 -133.675 0.475 -132.675 ;
        RECT 0.735 -133.675 0.965 -132.675 ;
        RECT 2.315 -133.675 2.545 -132.675 ;
        RECT 2.805 -133.675 3.035 -132.675 ;
        RECT 4.125 -133.675 4.355 -132.675 ;
        RECT 4.615 -133.675 4.845 -132.675 ;
        RECT 5.595 -133.675 5.825 -132.675 ;
        RECT 6.085 -133.675 6.315 -132.675 ;
        RECT 7.145 -133.675 7.375 -132.675 ;
        RECT 7.635 -133.675 7.865 -132.675 ;
        RECT 8.690 -133.675 8.920 -132.675 ;
        RECT 9.180 -133.675 9.410 -132.675 ;
        RECT 6.670 -133.865 7.325 -133.835 ;
        RECT 1.900 -134.005 7.325 -133.865 ;
        RECT -6.440 -135.065 -1.700 -134.925 ;
        RECT 0.270 -134.730 0.965 -134.665 ;
        RECT 1.900 -134.730 2.040 -134.005 ;
        RECT 6.670 -134.065 7.325 -134.005 ;
        RECT 0.270 -134.870 2.040 -134.730 ;
        RECT 4.015 -134.600 4.710 -134.515 ;
        RECT 8.200 -134.600 8.880 -134.555 ;
        RECT 4.015 -134.740 8.880 -134.600 ;
        RECT 4.015 -134.785 4.710 -134.740 ;
        RECT 8.200 -134.785 8.880 -134.740 ;
        RECT 0.270 -134.935 0.965 -134.870 ;
        RECT 6.060 -134.925 6.755 -134.885 ;
        RECT 9.135 -134.925 9.830 -134.855 ;
        RECT 10.535 -134.925 10.675 -130.885 ;
        RECT 11.370 -131.260 12.050 -131.030 ;
        RECT 11.635 -132.820 11.855 -131.260 ;
        RECT 25.895 -131.340 26.575 -131.110 ;
        RECT 11.630 -133.500 11.860 -132.820 ;
        RECT 12.745 -133.675 12.975 -132.675 ;
        RECT 13.235 -133.675 13.465 -132.675 ;
        RECT 14.815 -133.675 15.045 -132.675 ;
        RECT 15.305 -133.675 15.535 -132.675 ;
        RECT 16.625 -133.675 16.855 -132.675 ;
        RECT 17.115 -133.675 17.345 -132.675 ;
        RECT 18.095 -133.675 18.325 -132.675 ;
        RECT 18.585 -133.675 18.815 -132.675 ;
        RECT 19.645 -133.675 19.875 -132.675 ;
        RECT 20.135 -133.675 20.365 -132.675 ;
        RECT 21.190 -133.675 21.420 -132.675 ;
        RECT 21.680 -133.675 21.910 -132.675 ;
        RECT 26.160 -132.820 26.380 -131.340 ;
        RECT 47.065 -131.410 47.205 -98.310 ;
        RECT 27.060 -131.550 47.205 -131.410 ;
        RECT 26.155 -133.500 26.385 -132.820 ;
        RECT 19.170 -133.865 19.825 -133.835 ;
        RECT 14.400 -134.005 19.825 -133.865 ;
        RECT 6.060 -135.065 10.675 -134.925 ;
        RECT 12.770 -134.730 13.465 -134.665 ;
        RECT 14.400 -134.730 14.540 -134.005 ;
        RECT 19.170 -134.065 19.825 -134.005 ;
        RECT 12.770 -134.870 14.540 -134.730 ;
        RECT 16.515 -134.600 17.210 -134.515 ;
        RECT 20.700 -134.600 21.380 -134.555 ;
        RECT 16.515 -134.740 21.380 -134.600 ;
        RECT 16.515 -134.785 17.210 -134.740 ;
        RECT 20.700 -134.785 21.380 -134.740 ;
        RECT 12.770 -134.935 13.465 -134.870 ;
        RECT 18.560 -134.925 19.255 -134.885 ;
        RECT 21.635 -134.925 22.330 -134.855 ;
        RECT 27.060 -134.925 27.200 -131.550 ;
        RECT 27.745 -133.675 27.975 -132.675 ;
        RECT 28.235 -133.675 28.465 -132.675 ;
        RECT 29.815 -133.675 30.045 -132.675 ;
        RECT 30.305 -133.675 30.535 -132.675 ;
        RECT 31.625 -133.675 31.855 -132.675 ;
        RECT 32.115 -133.675 32.345 -132.675 ;
        RECT 33.095 -133.675 33.325 -132.675 ;
        RECT 33.585 -133.675 33.815 -132.675 ;
        RECT 34.645 -133.675 34.875 -132.675 ;
        RECT 35.135 -133.675 35.365 -132.675 ;
        RECT 36.190 -133.675 36.420 -132.675 ;
        RECT 36.680 -133.675 36.910 -132.675 ;
        RECT 34.170 -133.865 34.825 -133.835 ;
        RECT 29.400 -134.005 34.825 -133.865 ;
        RECT 18.560 -135.065 27.200 -134.925 ;
        RECT 27.770 -134.730 28.465 -134.665 ;
        RECT 29.400 -134.730 29.540 -134.005 ;
        RECT 34.170 -134.065 34.825 -134.005 ;
        RECT 27.770 -134.870 29.540 -134.730 ;
        RECT 31.515 -134.600 32.210 -134.515 ;
        RECT 35.700 -134.600 36.380 -134.555 ;
        RECT 31.515 -134.740 36.380 -134.600 ;
        RECT 31.515 -134.785 32.210 -134.740 ;
        RECT 35.700 -134.785 36.380 -134.740 ;
        RECT 27.770 -134.935 28.465 -134.870 ;
        RECT 33.560 -134.925 34.255 -134.885 ;
        RECT 36.635 -134.925 37.330 -134.855 ;
        RECT 47.845 -134.925 47.985 -94.795 ;
        RECT 33.560 -135.065 47.985 -134.925 ;
        RECT -31.440 -135.155 -30.745 -135.065 ;
        RECT -28.365 -135.125 -27.670 -135.065 ;
        RECT -18.940 -135.155 -18.245 -135.065 ;
        RECT -15.865 -135.125 -15.170 -135.065 ;
        RECT -6.440 -135.155 -5.745 -135.065 ;
        RECT -3.365 -135.125 -2.670 -135.065 ;
        RECT 6.060 -135.155 6.755 -135.065 ;
        RECT 9.135 -135.125 9.830 -135.065 ;
        RECT 18.560 -135.155 19.255 -135.065 ;
        RECT 21.635 -135.125 22.330 -135.065 ;
        RECT 33.560 -135.155 34.255 -135.065 ;
        RECT 36.635 -135.125 37.330 -135.065 ;
        RECT -37.255 -136.705 -37.025 -135.705 ;
        RECT -36.765 -136.705 -36.535 -135.705 ;
        RECT -36.275 -136.705 -36.045 -135.705 ;
        RECT -35.675 -136.705 -35.445 -135.705 ;
        RECT -35.185 -136.705 -34.955 -135.705 ;
        RECT -34.695 -136.705 -34.465 -135.705 ;
        RECT -32.885 -136.705 -32.655 -135.705 ;
        RECT -31.905 -136.705 -31.675 -135.705 ;
        RECT -30.355 -136.705 -30.125 -135.705 ;
        RECT -28.810 -136.705 -28.580 -135.705 ;
        RECT -24.755 -136.705 -24.525 -135.705 ;
        RECT -24.265 -136.705 -24.035 -135.705 ;
        RECT -23.775 -136.705 -23.545 -135.705 ;
        RECT -23.175 -136.705 -22.945 -135.705 ;
        RECT -22.685 -136.705 -22.455 -135.705 ;
        RECT -22.195 -136.705 -21.965 -135.705 ;
        RECT -20.385 -136.705 -20.155 -135.705 ;
        RECT -19.405 -136.705 -19.175 -135.705 ;
        RECT -17.855 -136.705 -17.625 -135.705 ;
        RECT -16.310 -136.705 -16.080 -135.705 ;
        RECT -12.255 -136.705 -12.025 -135.705 ;
        RECT -11.765 -136.705 -11.535 -135.705 ;
        RECT -11.275 -136.705 -11.045 -135.705 ;
        RECT -10.675 -136.705 -10.445 -135.705 ;
        RECT -10.185 -136.705 -9.955 -135.705 ;
        RECT -9.695 -136.705 -9.465 -135.705 ;
        RECT -7.885 -136.705 -7.655 -135.705 ;
        RECT -6.905 -136.705 -6.675 -135.705 ;
        RECT -5.355 -136.705 -5.125 -135.705 ;
        RECT -3.810 -136.705 -3.580 -135.705 ;
        RECT 0.245 -136.705 0.475 -135.705 ;
        RECT 0.735 -136.705 0.965 -135.705 ;
        RECT 1.225 -136.705 1.455 -135.705 ;
        RECT 1.825 -136.705 2.055 -135.705 ;
        RECT 2.315 -136.705 2.545 -135.705 ;
        RECT 2.805 -136.705 3.035 -135.705 ;
        RECT 4.615 -136.705 4.845 -135.705 ;
        RECT 5.595 -136.705 5.825 -135.705 ;
        RECT 7.145 -136.705 7.375 -135.705 ;
        RECT 8.690 -136.705 8.920 -135.705 ;
        RECT 12.745 -136.705 12.975 -135.705 ;
        RECT 13.235 -136.705 13.465 -135.705 ;
        RECT 13.725 -136.705 13.955 -135.705 ;
        RECT 14.325 -136.705 14.555 -135.705 ;
        RECT 14.815 -136.705 15.045 -135.705 ;
        RECT 15.305 -136.705 15.535 -135.705 ;
        RECT 17.115 -136.705 17.345 -135.705 ;
        RECT 18.095 -136.705 18.325 -135.705 ;
        RECT 19.645 -136.705 19.875 -135.705 ;
        RECT 21.190 -136.705 21.420 -135.705 ;
        RECT 27.745 -136.705 27.975 -135.705 ;
        RECT 28.235 -136.705 28.465 -135.705 ;
        RECT 28.725 -136.705 28.955 -135.705 ;
        RECT 29.325 -136.705 29.555 -135.705 ;
        RECT 29.815 -136.705 30.045 -135.705 ;
        RECT 30.305 -136.705 30.535 -135.705 ;
        RECT 32.115 -136.705 32.345 -135.705 ;
        RECT 33.095 -136.705 33.325 -135.705 ;
        RECT 34.645 -136.705 34.875 -135.705 ;
        RECT 36.190 -136.705 36.420 -135.705 ;
        RECT 49.295 -137.020 50.770 -100.570 ;
        RECT -98.520 -138.430 -97.830 -137.745 ;
        RECT -40.045 -138.520 -39.230 -137.645 ;
        RECT 44.035 -138.365 50.770 -137.020 ;
        RECT -99.210 -138.920 -98.525 -138.630 ;
        RECT -121.005 -149.725 -119.940 -148.835 ;
        RECT -39.990 -150.295 -39.330 -138.520 ;
        RECT 49.295 -149.675 50.770 -138.365 ;
        RECT 51.055 -132.925 52.055 -102.645 ;
        RECT 60.375 -120.355 61.720 -77.225 ;
        RECT 65.335 -81.890 390.960 -80.335 ;
        RECT 60.070 -122.060 62.000 -120.355 ;
        RECT 65.335 -121.805 66.590 -81.890 ;
        RECT 68.270 -84.140 344.620 -83.255 ;
        RECT 68.270 -115.555 69.925 -84.140 ;
        RECT 73.830 -86.935 301.075 -85.830 ;
        RECT 73.830 -106.655 74.280 -86.935 ;
        RECT 80.735 -89.720 255.130 -88.590 ;
        RECT 78.775 -92.120 211.005 -90.795 ;
        RECT 77.365 -94.150 168.600 -92.905 ;
        RECT 77.495 -97.550 80.320 -97.545 ;
        RECT 76.070 -98.250 80.320 -97.550 ;
        RECT 129.495 -99.710 161.820 -98.865 ;
        RECT 75.980 -100.355 127.145 -100.155 ;
        RECT 75.980 -101.825 128.045 -100.355 ;
        RECT 75.980 -101.915 127.870 -101.825 ;
        RECT 75.905 -102.860 77.240 -102.470 ;
        RECT 75.905 -103.635 125.475 -102.860 ;
        RECT 75.905 -103.960 77.240 -103.635 ;
        RECT 77.220 -106.180 81.355 -105.425 ;
        RECT 85.200 -106.135 86.095 -105.755 ;
        RECT 97.885 -106.095 98.115 -105.595 ;
        RECT 98.375 -106.095 98.605 -105.595 ;
        RECT 98.865 -106.095 99.095 -105.595 ;
        RECT 99.355 -106.095 99.585 -105.595 ;
        RECT 99.845 -106.095 100.075 -105.595 ;
        RECT 100.335 -106.095 100.565 -105.595 ;
        RECT 100.825 -106.095 101.055 -105.595 ;
        RECT 101.315 -106.095 101.545 -105.595 ;
        RECT 85.200 -106.510 93.550 -106.135 ;
        RECT 73.810 -107.475 74.300 -106.655 ;
        RECT 85.200 -106.700 86.095 -106.510 ;
        RECT 67.750 -117.680 70.320 -115.555 ;
        RECT 73.830 -118.300 74.280 -107.475 ;
        RECT 87.355 -107.690 87.585 -106.690 ;
        RECT 87.845 -107.690 88.075 -106.690 ;
        RECT 88.335 -107.690 88.565 -106.690 ;
        RECT 88.825 -107.690 89.055 -106.690 ;
        RECT 93.175 -106.885 93.550 -106.510 ;
        RECT 102.410 -106.520 102.640 -105.520 ;
        RECT 103.390 -106.520 103.620 -105.520 ;
        RECT 104.370 -106.520 104.600 -105.520 ;
        RECT 100.685 -106.785 101.530 -106.735 ;
        RECT 105.390 -106.785 105.675 -105.610 ;
        RECT 106.595 -106.520 106.825 -105.520 ;
        RECT 107.575 -106.520 107.805 -105.520 ;
        RECT 108.555 -106.520 108.785 -105.520 ;
        RECT 111.385 -106.095 111.615 -105.595 ;
        RECT 111.875 -106.095 112.105 -105.595 ;
        RECT 112.365 -106.095 112.595 -105.595 ;
        RECT 112.855 -106.095 113.085 -105.595 ;
        RECT 113.345 -106.095 113.575 -105.595 ;
        RECT 113.835 -106.095 114.065 -105.595 ;
        RECT 114.325 -106.095 114.555 -105.595 ;
        RECT 114.815 -106.095 115.045 -105.595 ;
        RECT 115.910 -106.520 116.140 -105.520 ;
        RECT 116.890 -106.520 117.120 -105.520 ;
        RECT 117.870 -106.520 118.100 -105.520 ;
        RECT 93.040 -107.560 93.700 -106.885 ;
        RECT 97.405 -107.310 98.175 -107.010 ;
        RECT 100.685 -107.070 105.675 -106.785 ;
        RECT 114.185 -106.785 115.030 -106.735 ;
        RECT 118.890 -106.785 119.175 -105.610 ;
        RECT 120.095 -106.520 120.325 -105.520 ;
        RECT 121.075 -106.520 121.305 -105.520 ;
        RECT 122.055 -106.520 122.285 -105.520 ;
        RECT 109.670 -106.895 109.970 -106.865 ;
        RECT 100.685 -107.105 101.530 -107.070 ;
        RECT 109.255 -107.195 109.970 -106.895 ;
        RECT 110.940 -107.000 111.145 -106.995 ;
        RECT 91.535 -107.880 91.745 -107.860 ;
        RECT 91.125 -108.180 91.785 -107.880 ;
        RECT 87.355 -112.510 87.585 -109.510 ;
        RECT 88.415 -112.510 88.645 -109.510 ;
        RECT 88.905 -112.510 89.135 -109.510 ;
        RECT 89.395 -112.510 89.625 -109.510 ;
        RECT 89.960 -112.510 90.190 -109.510 ;
        RECT 90.450 -112.510 90.680 -109.510 ;
        RECT 90.940 -112.510 91.170 -109.510 ;
        RECT 76.530 -117.195 87.080 -116.215 ;
        RECT 86.100 -117.225 87.080 -117.195 ;
        RECT 86.100 -117.995 87.090 -117.225 ;
        RECT 86.065 -118.205 91.250 -117.995 ;
        RECT 73.830 -118.365 83.745 -118.300 ;
        RECT 73.830 -118.575 90.800 -118.365 ;
        RECT 73.830 -118.750 83.745 -118.575 ;
        RECT 87.330 -120.780 87.560 -119.780 ;
        RECT 87.820 -120.780 88.050 -119.780 ;
        RECT 88.310 -120.780 88.540 -119.780 ;
        RECT 89.380 -121.305 90.040 -121.005 ;
        RECT 65.255 -122.955 66.695 -121.805 ;
        RECT 89.815 -121.870 90.025 -121.305 ;
        RECT 90.590 -121.430 90.800 -118.575 ;
        RECT 91.040 -121.010 91.250 -118.205 ;
        RECT 91.535 -118.350 91.745 -108.180 ;
        RECT 91.985 -108.485 96.535 -108.200 ;
        RECT 91.985 -115.240 92.270 -108.485 ;
        RECT 94.770 -109.065 95.430 -108.765 ;
        RECT 94.870 -110.110 95.345 -109.065 ;
        RECT 96.250 -109.090 96.535 -108.485 ;
        RECT 97.405 -108.685 97.635 -107.310 ;
        RECT 97.885 -108.170 98.115 -107.670 ;
        RECT 98.375 -108.170 98.605 -107.670 ;
        RECT 98.865 -108.170 99.095 -107.670 ;
        RECT 99.355 -108.170 99.585 -107.670 ;
        RECT 99.845 -108.170 100.075 -107.670 ;
        RECT 100.335 -108.170 100.565 -107.670 ;
        RECT 100.825 -108.170 101.055 -107.670 ;
        RECT 101.315 -108.170 101.545 -107.670 ;
        RECT 102.410 -107.920 102.640 -107.420 ;
        RECT 102.900 -107.920 103.130 -107.420 ;
        RECT 103.390 -107.920 103.620 -107.420 ;
        RECT 103.880 -107.920 104.110 -107.420 ;
        RECT 104.370 -107.920 104.600 -107.420 ;
        RECT 104.860 -107.920 105.090 -107.420 ;
        RECT 97.405 -108.910 101.500 -108.685 ;
        RECT 97.445 -108.915 101.500 -108.910 ;
        RECT 96.250 -109.375 97.580 -109.090 ;
        RECT 96.385 -109.915 97.045 -109.615 ;
        RECT 94.835 -110.410 95.520 -110.110 ;
        RECT 93.470 -111.210 93.700 -110.710 ;
        RECT 93.960 -111.210 94.190 -110.710 ;
        RECT 94.450 -111.210 94.680 -110.710 ;
        RECT 94.940 -111.210 95.170 -110.710 ;
        RECT 95.430 -111.210 95.660 -110.710 ;
        RECT 95.920 -111.210 96.150 -110.710 ;
        RECT 96.590 -111.055 96.880 -109.915 ;
        RECT 96.590 -111.715 96.890 -111.055 ;
        RECT 97.295 -111.560 97.580 -109.375 ;
        RECT 101.270 -109.745 101.500 -108.915 ;
        RECT 105.620 -109.185 105.920 -107.365 ;
        RECT 106.595 -107.920 106.825 -107.420 ;
        RECT 107.085 -107.920 107.315 -107.420 ;
        RECT 107.575 -107.920 107.805 -107.420 ;
        RECT 108.065 -107.920 108.295 -107.420 ;
        RECT 108.555 -107.920 108.785 -107.420 ;
        RECT 109.045 -107.920 109.275 -107.420 ;
        RECT 107.935 -109.065 108.620 -108.765 ;
        RECT 105.405 -109.485 106.065 -109.185 ;
        RECT 101.270 -109.975 105.070 -109.745 ;
        RECT 101.930 -110.460 102.140 -109.975 ;
        RECT 102.910 -110.460 103.120 -109.975 ;
        RECT 103.885 -110.460 104.095 -109.975 ;
        RECT 104.840 -110.460 105.070 -109.975 ;
        RECT 108.090 -110.105 108.565 -109.065 ;
        RECT 107.970 -110.405 108.655 -110.105 ;
        RECT 97.880 -111.210 98.110 -110.710 ;
        RECT 98.370 -111.210 98.600 -110.710 ;
        RECT 98.860 -111.210 99.090 -110.710 ;
        RECT 99.350 -111.210 99.580 -110.710 ;
        RECT 99.840 -111.210 100.070 -110.710 ;
        RECT 100.330 -111.210 100.560 -110.710 ;
        RECT 101.425 -110.960 101.655 -110.460 ;
        RECT 101.915 -110.960 102.145 -110.460 ;
        RECT 102.405 -110.960 102.635 -110.460 ;
        RECT 102.895 -110.960 103.125 -110.460 ;
        RECT 103.385 -110.960 103.615 -110.460 ;
        RECT 103.875 -110.960 104.105 -110.460 ;
        RECT 104.365 -110.960 104.595 -110.460 ;
        RECT 104.840 -110.960 105.085 -110.460 ;
        RECT 106.595 -111.210 106.825 -110.710 ;
        RECT 107.085 -111.210 107.315 -110.710 ;
        RECT 107.575 -111.210 107.805 -110.710 ;
        RECT 108.065 -111.210 108.295 -110.710 ;
        RECT 108.555 -111.210 108.785 -110.710 ;
        RECT 109.045 -111.210 109.275 -110.710 ;
        RECT 109.670 -110.935 109.970 -107.195 ;
        RECT 110.935 -107.300 111.620 -107.000 ;
        RECT 114.185 -107.070 119.175 -106.785 ;
        RECT 114.185 -107.105 115.030 -107.070 ;
        RECT 110.110 -109.480 110.795 -109.180 ;
        RECT 109.670 -111.160 109.975 -110.935 ;
        RECT 101.440 -111.560 102.285 -111.525 ;
        RECT 97.295 -111.845 102.285 -111.560 ;
        RECT 109.675 -111.595 109.975 -111.160 ;
        RECT 110.250 -111.720 110.550 -109.480 ;
        RECT 110.940 -109.725 111.145 -107.300 ;
        RECT 111.385 -108.170 111.615 -107.670 ;
        RECT 111.875 -108.170 112.105 -107.670 ;
        RECT 112.365 -108.170 112.595 -107.670 ;
        RECT 112.855 -108.170 113.085 -107.670 ;
        RECT 113.345 -108.170 113.575 -107.670 ;
        RECT 113.835 -108.170 114.065 -107.670 ;
        RECT 114.325 -108.170 114.555 -107.670 ;
        RECT 114.815 -108.170 115.045 -107.670 ;
        RECT 115.910 -107.920 116.140 -107.420 ;
        RECT 116.400 -107.920 116.630 -107.420 ;
        RECT 116.890 -107.920 117.120 -107.420 ;
        RECT 117.380 -107.920 117.610 -107.420 ;
        RECT 117.870 -107.920 118.100 -107.420 ;
        RECT 118.360 -107.920 118.590 -107.420 ;
        RECT 119.180 -109.625 119.480 -107.290 ;
        RECT 120.095 -107.920 120.325 -107.420 ;
        RECT 120.585 -107.920 120.815 -107.420 ;
        RECT 121.075 -107.920 121.305 -107.420 ;
        RECT 121.565 -107.920 121.795 -107.420 ;
        RECT 122.055 -107.920 122.285 -107.420 ;
        RECT 122.545 -107.920 122.775 -107.420 ;
        RECT 120.920 -109.035 121.605 -108.735 ;
        RECT 110.940 -109.965 118.595 -109.725 ;
        RECT 119.000 -109.925 119.660 -109.625 ;
        RECT 111.380 -111.210 111.610 -110.710 ;
        RECT 111.870 -111.210 112.100 -110.710 ;
        RECT 112.360 -111.210 112.590 -110.710 ;
        RECT 112.850 -111.210 113.080 -110.710 ;
        RECT 113.340 -111.210 113.570 -110.710 ;
        RECT 113.830 -111.210 114.060 -110.710 ;
        RECT 114.925 -110.960 115.155 -110.460 ;
        RECT 115.395 -110.555 115.700 -109.965 ;
        RECT 115.415 -110.960 115.645 -110.555 ;
        RECT 115.905 -110.960 116.135 -110.460 ;
        RECT 116.350 -110.565 116.655 -109.965 ;
        RECT 116.395 -110.960 116.625 -110.565 ;
        RECT 116.885 -110.960 117.115 -110.460 ;
        RECT 117.330 -110.555 117.635 -109.965 ;
        RECT 117.375 -110.960 117.605 -110.555 ;
        RECT 117.865 -110.960 118.095 -110.460 ;
        RECT 118.355 -110.735 118.595 -109.965 ;
        RECT 121.055 -110.125 121.530 -109.035 ;
        RECT 123.045 -109.325 123.345 -109.090 ;
        RECT 123.045 -109.645 124.390 -109.325 ;
        RECT 123.045 -109.775 123.775 -109.645 ;
        RECT 120.990 -110.425 121.650 -110.125 ;
        RECT 118.355 -110.960 118.585 -110.735 ;
        RECT 120.095 -111.210 120.325 -110.710 ;
        RECT 120.585 -111.210 120.815 -110.710 ;
        RECT 121.075 -111.210 121.305 -110.710 ;
        RECT 121.565 -111.210 121.795 -110.710 ;
        RECT 122.055 -111.210 122.285 -110.710 ;
        RECT 122.545 -111.210 122.775 -110.710 ;
        RECT 114.940 -111.560 115.785 -111.525 ;
        RECT 93.960 -113.110 94.190 -112.110 ;
        RECT 94.940 -113.110 95.170 -112.110 ;
        RECT 95.920 -113.110 96.150 -112.110 ;
        RECT 97.295 -113.020 97.580 -111.845 ;
        RECT 101.440 -111.895 102.285 -111.845 ;
        RECT 110.795 -111.845 115.785 -111.560 ;
        RECT 98.370 -113.110 98.600 -112.110 ;
        RECT 99.350 -113.110 99.580 -112.110 ;
        RECT 100.330 -113.110 100.560 -112.110 ;
        RECT 101.425 -113.035 101.655 -112.535 ;
        RECT 101.915 -113.035 102.145 -112.535 ;
        RECT 102.405 -113.035 102.635 -112.535 ;
        RECT 102.895 -113.035 103.125 -112.535 ;
        RECT 103.385 -113.035 103.615 -112.535 ;
        RECT 103.875 -113.035 104.105 -112.535 ;
        RECT 104.365 -113.035 104.595 -112.535 ;
        RECT 104.855 -113.035 105.085 -112.535 ;
        RECT 107.085 -113.110 107.315 -112.110 ;
        RECT 108.065 -113.110 108.295 -112.110 ;
        RECT 109.045 -113.110 109.275 -112.110 ;
        RECT 110.795 -113.020 111.080 -111.845 ;
        RECT 114.940 -111.895 115.785 -111.845 ;
        RECT 111.870 -113.110 112.100 -112.110 ;
        RECT 112.850 -113.110 113.080 -112.110 ;
        RECT 113.830 -113.110 114.060 -112.110 ;
        RECT 114.925 -113.035 115.155 -112.535 ;
        RECT 115.415 -113.035 115.645 -112.535 ;
        RECT 115.905 -113.035 116.135 -112.535 ;
        RECT 116.395 -113.035 116.625 -112.535 ;
        RECT 116.885 -113.035 117.115 -112.535 ;
        RECT 117.375 -113.035 117.605 -112.535 ;
        RECT 117.865 -113.035 118.095 -112.535 ;
        RECT 118.355 -113.035 118.585 -112.535 ;
        RECT 120.585 -113.110 120.815 -112.110 ;
        RECT 121.565 -113.110 121.795 -112.110 ;
        RECT 122.545 -113.110 122.775 -112.110 ;
        RECT 123.325 -113.995 123.775 -109.775 ;
        RECT 103.615 -114.445 123.775 -113.995 ;
        RECT 103.615 -114.900 104.415 -114.445 ;
        RECT 91.985 -115.525 108.345 -115.240 ;
        RECT 103.600 -116.475 104.400 -115.815 ;
        RECT 91.535 -118.560 95.385 -118.350 ;
        RECT 103.085 -118.390 103.745 -118.090 ;
        RECT 92.060 -120.780 92.290 -119.780 ;
        RECT 92.550 -120.780 92.780 -119.780 ;
        RECT 93.040 -120.780 93.270 -119.780 ;
        RECT 91.620 -121.010 92.280 -120.975 ;
        RECT 91.040 -121.220 92.280 -121.010 ;
        RECT 91.620 -121.275 92.280 -121.220 ;
        RECT 92.735 -121.430 93.395 -121.375 ;
        RECT 90.590 -121.640 93.395 -121.430 ;
        RECT 92.735 -121.675 93.395 -121.640 ;
        RECT 94.560 -121.870 94.860 -121.720 ;
        RECT 89.815 -122.080 94.860 -121.870 ;
        RECT 87.330 -124.240 87.560 -122.240 ;
        RECT 88.385 -124.240 88.615 -122.240 ;
        RECT 88.875 -124.240 89.105 -122.240 ;
        RECT 89.365 -124.240 89.595 -122.240 ;
        RECT 92.060 -124.240 92.290 -122.240 ;
        RECT 93.115 -124.240 93.345 -122.240 ;
        RECT 93.605 -124.240 93.835 -122.240 ;
        RECT 94.095 -124.240 94.325 -122.240 ;
        RECT 94.560 -122.380 94.860 -122.080 ;
        RECT 95.175 -122.970 95.385 -118.560 ;
        RECT 96.150 -121.375 96.380 -119.875 ;
        RECT 96.640 -121.375 96.870 -119.875 ;
        RECT 97.130 -121.375 97.360 -119.875 ;
        RECT 97.700 -121.370 97.930 -119.870 ;
        RECT 98.190 -121.370 98.420 -119.870 ;
        RECT 98.680 -121.370 98.910 -119.870 ;
        RECT 99.245 -121.370 99.475 -119.870 ;
        RECT 99.735 -121.370 99.965 -119.870 ;
        RECT 100.225 -121.370 100.455 -119.870 ;
        RECT 101.800 -120.870 102.030 -119.870 ;
        RECT 102.290 -120.870 102.520 -119.870 ;
        RECT 103.245 -121.815 103.545 -118.390 ;
        RECT 103.940 -118.595 104.240 -116.475 ;
        RECT 106.185 -117.870 106.415 -115.870 ;
        RECT 107.165 -117.870 107.395 -115.870 ;
        RECT 108.060 -118.135 108.345 -115.525 ;
        RECT 124.700 -115.580 125.475 -103.635 ;
        RECT 109.040 -115.930 125.475 -115.580 ;
        RECT 109.040 -116.825 109.390 -115.930 ;
        RECT 103.940 -118.600 105.645 -118.595 ;
        RECT 103.940 -118.890 105.650 -118.600 ;
        RECT 107.915 -118.805 108.345 -118.135 ;
        RECT 103.940 -118.895 105.645 -118.890 ;
        RECT 103.050 -122.115 103.705 -121.815 ;
        RECT 103.940 -122.665 104.240 -118.895 ;
        RECT 105.695 -120.140 105.925 -119.140 ;
        RECT 106.185 -120.140 106.415 -119.140 ;
        RECT 106.745 -120.140 106.975 -119.140 ;
        RECT 107.235 -120.140 107.465 -119.140 ;
        RECT 109.845 -119.595 110.075 -116.095 ;
        RECT 110.335 -119.595 110.565 -116.095 ;
        RECT 111.845 -119.595 112.075 -116.095 ;
        RECT 112.335 -119.595 112.565 -116.095 ;
        RECT 114.260 -119.580 114.610 -115.930 ;
        RECT 114.845 -119.595 115.075 -116.095 ;
        RECT 115.335 -119.595 115.565 -116.095 ;
        RECT 116.845 -119.595 117.075 -116.095 ;
        RECT 117.335 -119.595 117.565 -116.095 ;
        RECT 119.215 -119.585 119.565 -115.930 ;
        RECT 119.845 -119.595 120.075 -116.095 ;
        RECT 120.335 -119.595 120.565 -116.095 ;
        RECT 121.845 -119.595 122.075 -116.095 ;
        RECT 122.335 -119.595 122.565 -116.095 ;
        RECT 112.905 -119.845 113.495 -119.785 ;
        RECT 112.905 -120.015 113.940 -119.845 ;
        RECT 122.770 -119.880 123.360 -119.860 ;
        RECT 125.525 -119.880 126.130 -119.765 ;
        RECT 112.905 -120.075 113.495 -120.015 ;
        RECT 105.445 -122.475 105.675 -121.975 ;
        RECT 105.935 -122.475 106.165 -121.975 ;
        RECT 106.425 -122.475 106.655 -121.975 ;
        RECT 106.915 -122.475 107.145 -121.975 ;
        RECT 107.405 -122.475 107.635 -121.975 ;
        RECT 107.895 -122.475 108.125 -121.975 ;
        RECT 103.940 -122.965 105.575 -122.665 ;
        RECT 95.135 -123.630 95.435 -122.970 ;
        RECT 96.640 -124.410 96.870 -123.410 ;
        RECT 97.620 -124.410 97.850 -123.410 ;
        RECT 98.600 -124.410 98.830 -123.410 ;
        RECT 102.290 -124.410 102.520 -123.410 ;
        RECT 105.935 -124.375 106.165 -123.375 ;
        RECT 106.915 -124.375 107.145 -123.375 ;
        RECT 107.895 -124.375 108.125 -123.375 ;
        RECT 110.335 -124.020 110.565 -120.520 ;
        RECT 112.335 -124.020 112.565 -120.520 ;
        RECT 113.770 -124.520 113.940 -120.015 ;
        RECT 118.290 -120.210 118.880 -119.920 ;
        RECT 122.770 -120.105 126.130 -119.880 ;
        RECT 122.770 -120.150 123.360 -120.105 ;
        RECT 115.335 -124.020 115.565 -120.520 ;
        RECT 117.335 -124.020 117.565 -120.520 ;
        RECT 118.320 -124.195 118.490 -120.210 ;
        RECT 120.335 -124.020 120.565 -120.520 ;
        RECT 122.335 -124.020 122.565 -120.520 ;
        RECT 118.320 -124.365 124.860 -124.195 ;
        RECT 113.770 -124.690 124.420 -124.520 ;
        RECT 53.320 -129.300 53.550 -128.300 ;
        RECT 54.300 -129.300 54.530 -128.300 ;
        RECT 55.280 -129.300 55.510 -128.300 ;
        RECT 56.655 -129.565 56.940 -128.390 ;
        RECT 57.730 -129.300 57.960 -128.300 ;
        RECT 58.710 -129.300 58.940 -128.300 ;
        RECT 59.690 -129.300 59.920 -128.300 ;
        RECT 60.785 -128.875 61.015 -128.375 ;
        RECT 61.275 -128.875 61.505 -128.375 ;
        RECT 61.765 -128.875 61.995 -128.375 ;
        RECT 62.255 -128.875 62.485 -128.375 ;
        RECT 62.745 -128.875 62.975 -128.375 ;
        RECT 63.235 -128.875 63.465 -128.375 ;
        RECT 63.725 -128.875 63.955 -128.375 ;
        RECT 64.215 -128.875 64.445 -128.375 ;
        RECT 66.445 -129.300 66.675 -128.300 ;
        RECT 67.425 -129.300 67.655 -128.300 ;
        RECT 68.405 -129.300 68.635 -128.300 ;
        RECT 60.800 -129.565 61.645 -129.515 ;
        RECT 52.830 -130.700 53.060 -130.200 ;
        RECT 53.320 -130.700 53.550 -130.200 ;
        RECT 53.810 -130.700 54.040 -130.200 ;
        RECT 54.300 -130.700 54.530 -130.200 ;
        RECT 54.790 -130.700 55.020 -130.200 ;
        RECT 55.280 -130.700 55.510 -130.200 ;
        RECT 55.950 -130.355 56.250 -129.695 ;
        RECT 56.655 -129.850 61.645 -129.565 ;
        RECT 70.155 -129.565 70.440 -128.390 ;
        RECT 71.230 -129.300 71.460 -128.300 ;
        RECT 72.210 -129.300 72.440 -128.300 ;
        RECT 73.190 -129.300 73.420 -128.300 ;
        RECT 74.285 -128.875 74.515 -128.375 ;
        RECT 74.775 -128.875 75.005 -128.375 ;
        RECT 75.265 -128.875 75.495 -128.375 ;
        RECT 75.755 -128.875 75.985 -128.375 ;
        RECT 76.245 -128.875 76.475 -128.375 ;
        RECT 76.735 -128.875 76.965 -128.375 ;
        RECT 77.225 -128.875 77.455 -128.375 ;
        RECT 77.715 -128.875 77.945 -128.375 ;
        RECT 79.945 -129.300 80.175 -128.300 ;
        RECT 80.925 -129.300 81.155 -128.300 ;
        RECT 81.905 -129.300 82.135 -128.300 ;
        RECT 74.300 -129.565 75.145 -129.515 ;
        RECT 54.195 -131.300 54.880 -131.000 ;
        RECT 54.230 -132.345 54.705 -131.300 ;
        RECT 55.950 -131.495 56.240 -130.355 ;
        RECT 55.745 -131.795 56.405 -131.495 ;
        RECT 56.655 -132.035 56.940 -129.850 ;
        RECT 60.800 -129.885 61.645 -129.850 ;
        RECT 57.240 -130.700 57.470 -130.200 ;
        RECT 57.730 -130.700 57.960 -130.200 ;
        RECT 58.220 -130.700 58.450 -130.200 ;
        RECT 58.710 -130.700 58.940 -130.200 ;
        RECT 59.200 -130.700 59.430 -130.200 ;
        RECT 59.690 -130.700 59.920 -130.200 ;
        RECT 60.785 -130.950 61.015 -130.450 ;
        RECT 61.275 -130.950 61.505 -130.450 ;
        RECT 61.765 -130.950 61.995 -130.450 ;
        RECT 62.255 -130.950 62.485 -130.450 ;
        RECT 62.745 -130.950 62.975 -130.450 ;
        RECT 63.235 -130.950 63.465 -130.450 ;
        RECT 63.725 -130.950 63.955 -130.450 ;
        RECT 64.200 -130.950 64.445 -130.450 ;
        RECT 65.955 -130.700 66.185 -130.200 ;
        RECT 66.445 -130.700 66.675 -130.200 ;
        RECT 66.935 -130.700 67.165 -130.200 ;
        RECT 67.425 -130.700 67.655 -130.200 ;
        RECT 67.915 -130.700 68.145 -130.200 ;
        RECT 68.405 -130.700 68.635 -130.200 ;
        RECT 69.035 -130.250 69.335 -129.815 ;
        RECT 69.030 -130.475 69.335 -130.250 ;
        RECT 61.290 -131.435 61.500 -130.950 ;
        RECT 62.270 -131.435 62.480 -130.950 ;
        RECT 63.245 -131.435 63.455 -130.950 ;
        RECT 64.200 -131.435 64.430 -130.950 ;
        RECT 67.330 -131.305 68.015 -131.005 ;
        RECT 55.610 -132.320 56.940 -132.035 ;
        RECT 60.630 -131.665 64.430 -131.435 ;
        RECT 54.130 -132.645 54.790 -132.345 ;
        RECT 55.610 -132.925 55.895 -132.320 ;
        RECT 60.630 -132.495 60.860 -131.665 ;
        RECT 64.765 -132.225 65.425 -131.925 ;
        RECT 56.805 -132.500 60.860 -132.495 ;
        RECT 51.055 -133.210 55.895 -132.925 ;
        RECT 56.765 -132.725 60.860 -132.500 ;
        RECT -39.990 -150.975 -39.310 -150.295 ;
        RECT 51.055 -152.160 52.055 -133.210 ;
        RECT 56.765 -134.100 56.995 -132.725 ;
        RECT 57.245 -133.740 57.475 -133.240 ;
        RECT 57.735 -133.740 57.965 -133.240 ;
        RECT 58.225 -133.740 58.455 -133.240 ;
        RECT 58.715 -133.740 58.945 -133.240 ;
        RECT 59.205 -133.740 59.435 -133.240 ;
        RECT 59.695 -133.740 59.925 -133.240 ;
        RECT 60.185 -133.740 60.415 -133.240 ;
        RECT 60.675 -133.740 60.905 -133.240 ;
        RECT 61.770 -133.990 62.000 -133.490 ;
        RECT 62.260 -133.990 62.490 -133.490 ;
        RECT 62.750 -133.990 62.980 -133.490 ;
        RECT 63.240 -133.990 63.470 -133.490 ;
        RECT 63.730 -133.990 63.960 -133.490 ;
        RECT 64.220 -133.990 64.450 -133.490 ;
        RECT 64.980 -134.045 65.280 -132.225 ;
        RECT 67.450 -132.345 67.925 -131.305 ;
        RECT 67.295 -132.645 67.980 -132.345 ;
        RECT 65.955 -133.990 66.185 -133.490 ;
        RECT 66.445 -133.990 66.675 -133.490 ;
        RECT 66.935 -133.990 67.165 -133.490 ;
        RECT 67.425 -133.990 67.655 -133.490 ;
        RECT 67.915 -133.990 68.145 -133.490 ;
        RECT 68.405 -133.990 68.635 -133.490 ;
        RECT 56.765 -134.400 57.535 -134.100 ;
        RECT 69.030 -134.215 69.330 -130.475 ;
        RECT 69.610 -131.930 69.910 -129.690 ;
        RECT 70.155 -129.850 75.145 -129.565 ;
        RECT 74.300 -129.885 75.145 -129.850 ;
        RECT 70.740 -130.700 70.970 -130.200 ;
        RECT 71.230 -130.700 71.460 -130.200 ;
        RECT 71.720 -130.700 71.950 -130.200 ;
        RECT 72.210 -130.700 72.440 -130.200 ;
        RECT 72.700 -130.700 72.930 -130.200 ;
        RECT 73.190 -130.700 73.420 -130.200 ;
        RECT 74.285 -130.950 74.515 -130.450 ;
        RECT 74.775 -130.855 75.005 -130.450 ;
        RECT 74.755 -131.445 75.060 -130.855 ;
        RECT 75.265 -130.950 75.495 -130.450 ;
        RECT 75.755 -130.845 75.985 -130.450 ;
        RECT 75.710 -131.445 76.015 -130.845 ;
        RECT 76.245 -130.950 76.475 -130.450 ;
        RECT 76.735 -130.855 76.965 -130.450 ;
        RECT 76.690 -131.445 76.995 -130.855 ;
        RECT 77.225 -130.950 77.455 -130.450 ;
        RECT 77.715 -130.675 77.945 -130.450 ;
        RECT 77.715 -131.445 77.955 -130.675 ;
        RECT 79.455 -130.700 79.685 -130.200 ;
        RECT 79.945 -130.700 80.175 -130.200 ;
        RECT 80.435 -130.700 80.665 -130.200 ;
        RECT 80.925 -130.700 81.155 -130.200 ;
        RECT 81.415 -130.700 81.645 -130.200 ;
        RECT 81.905 -130.700 82.135 -130.200 ;
        RECT 80.350 -131.285 81.010 -130.985 ;
        RECT 70.300 -131.685 77.955 -131.445 ;
        RECT 69.470 -132.230 70.155 -131.930 ;
        RECT 70.300 -134.110 70.505 -131.685 ;
        RECT 78.360 -131.785 79.020 -131.485 ;
        RECT 70.745 -133.740 70.975 -133.240 ;
        RECT 71.235 -133.740 71.465 -133.240 ;
        RECT 71.725 -133.740 71.955 -133.240 ;
        RECT 72.215 -133.740 72.445 -133.240 ;
        RECT 72.705 -133.740 72.935 -133.240 ;
        RECT 73.195 -133.740 73.425 -133.240 ;
        RECT 73.685 -133.740 73.915 -133.240 ;
        RECT 74.175 -133.740 74.405 -133.240 ;
        RECT 75.270 -133.990 75.500 -133.490 ;
        RECT 75.760 -133.990 75.990 -133.490 ;
        RECT 76.250 -133.990 76.480 -133.490 ;
        RECT 76.740 -133.990 76.970 -133.490 ;
        RECT 77.230 -133.990 77.460 -133.490 ;
        RECT 77.720 -133.990 77.950 -133.490 ;
        RECT 60.045 -134.340 60.890 -134.305 ;
        RECT 60.045 -134.625 65.035 -134.340 ;
        RECT 68.615 -134.515 69.330 -134.215 ;
        RECT 70.295 -134.410 70.980 -134.110 ;
        RECT 78.540 -134.120 78.840 -131.785 ;
        RECT 80.415 -132.375 80.890 -131.285 ;
        RECT 82.405 -131.765 82.705 -131.635 ;
        RECT 82.405 -132.085 84.685 -131.765 ;
        RECT 82.405 -132.320 82.705 -132.085 ;
        RECT 80.280 -132.675 80.965 -132.375 ;
        RECT 79.455 -133.990 79.685 -133.490 ;
        RECT 79.945 -133.990 80.175 -133.490 ;
        RECT 80.435 -133.990 80.665 -133.490 ;
        RECT 80.925 -133.990 81.155 -133.490 ;
        RECT 81.415 -133.990 81.645 -133.490 ;
        RECT 81.905 -133.990 82.135 -133.490 ;
        RECT 73.545 -134.340 74.390 -134.305 ;
        RECT 70.300 -134.415 70.505 -134.410 ;
        RECT 69.030 -134.545 69.330 -134.515 ;
        RECT 60.045 -134.675 60.890 -134.625 ;
        RECT 57.245 -135.815 57.475 -135.315 ;
        RECT 57.735 -135.815 57.965 -135.315 ;
        RECT 58.225 -135.815 58.455 -135.315 ;
        RECT 58.715 -135.815 58.945 -135.315 ;
        RECT 59.205 -135.815 59.435 -135.315 ;
        RECT 59.695 -135.815 59.925 -135.315 ;
        RECT 60.185 -135.815 60.415 -135.315 ;
        RECT 60.675 -135.815 60.905 -135.315 ;
        RECT 61.770 -135.890 62.000 -134.890 ;
        RECT 62.750 -135.890 62.980 -134.890 ;
        RECT 63.730 -135.890 63.960 -134.890 ;
        RECT 64.750 -135.800 65.035 -134.625 ;
        RECT 73.545 -134.625 78.535 -134.340 ;
        RECT 73.545 -134.675 74.390 -134.625 ;
        RECT 65.955 -135.890 66.185 -134.890 ;
        RECT 66.935 -135.890 67.165 -134.890 ;
        RECT 67.915 -135.890 68.145 -134.890 ;
        RECT 70.745 -135.815 70.975 -135.315 ;
        RECT 71.235 -135.815 71.465 -135.315 ;
        RECT 71.725 -135.815 71.955 -135.315 ;
        RECT 72.215 -135.815 72.445 -135.315 ;
        RECT 72.705 -135.815 72.935 -135.315 ;
        RECT 73.195 -135.815 73.425 -135.315 ;
        RECT 73.685 -135.815 73.915 -135.315 ;
        RECT 74.175 -135.815 74.405 -135.315 ;
        RECT 75.270 -135.890 75.500 -134.890 ;
        RECT 76.250 -135.890 76.480 -134.890 ;
        RECT 77.230 -135.890 77.460 -134.890 ;
        RECT 78.250 -135.800 78.535 -134.625 ;
        RECT 79.455 -135.890 79.685 -134.890 ;
        RECT 80.435 -135.890 80.665 -134.890 ;
        RECT 81.415 -135.890 81.645 -134.890 ;
        RECT 84.045 -150.295 84.685 -132.085 ;
        RECT 121.555 -135.545 121.905 -124.690 ;
        RECT 124.690 -125.005 124.860 -124.365 ;
        RECT 120.960 -136.645 122.815 -135.545 ;
        RECT 124.385 -138.290 124.990 -125.005 ;
        RECT 84.020 -150.975 84.685 -150.295 ;
        RECT 117.985 -138.895 124.990 -138.290 ;
        RECT 117.985 -153.110 118.590 -138.895 ;
        RECT 125.525 -150.100 126.130 -120.105 ;
        RECT 126.645 -137.410 127.870 -101.915 ;
        RECT 129.495 -117.950 130.340 -99.710 ;
        RECT 130.985 -101.115 132.050 -100.920 ;
        RECT 139.620 -101.035 141.815 -100.800 ;
        RECT 130.985 -101.385 138.175 -101.115 ;
        RECT 139.620 -101.220 139.855 -101.035 ;
        RECT 130.985 -101.585 132.050 -101.385 ;
        RECT 133.820 -103.585 134.470 -102.835 ;
        RECT 135.250 -103.105 135.480 -102.105 ;
        RECT 135.740 -103.245 135.970 -102.105 ;
        RECT 136.230 -103.105 136.460 -102.105 ;
        RECT 136.720 -103.245 136.950 -102.105 ;
        RECT 137.905 -102.835 138.175 -101.385 ;
        RECT 139.625 -102.715 139.855 -101.220 ;
        RECT 140.115 -102.715 140.345 -101.215 ;
        RECT 140.605 -102.715 140.835 -101.035 ;
        RECT 137.905 -103.105 139.545 -102.835 ;
        RECT 135.250 -103.475 138.435 -103.245 ;
        RECT 139.275 -103.380 139.545 -103.105 ;
        RECT 130.990 -110.720 132.285 -109.405 ;
        RECT 134.070 -110.605 134.340 -103.585 ;
        RECT 135.250 -104.755 135.480 -103.475 ;
        RECT 135.740 -103.485 136.950 -103.475 ;
        RECT 136.230 -104.755 136.460 -103.485 ;
        RECT 137.210 -104.755 137.440 -103.475 ;
        RECT 139.145 -103.670 139.940 -103.380 ;
        RECT 140.115 -105.400 140.345 -103.900 ;
        RECT 141.095 -105.400 141.325 -101.215 ;
        RECT 141.585 -102.715 141.815 -101.035 ;
        RECT 145.095 -103.575 148.635 -103.010 ;
        RECT 143.160 -104.250 143.390 -103.750 ;
        RECT 143.650 -104.395 143.880 -103.750 ;
        RECT 144.140 -104.250 144.370 -103.750 ;
        RECT 144.630 -104.395 144.860 -103.750 ;
        RECT 143.160 -104.625 146.345 -104.395 ;
        RECT 143.160 -105.405 143.390 -104.625 ;
        RECT 143.650 -104.635 144.860 -104.625 ;
        RECT 144.140 -105.405 144.370 -104.635 ;
        RECT 145.120 -105.405 145.350 -104.625 ;
        RECT 135.120 -109.900 135.350 -108.400 ;
        RECT 133.355 -110.875 134.340 -110.605 ;
        RECT 134.630 -112.580 134.860 -111.085 ;
        RECT 134.625 -112.765 134.860 -112.580 ;
        RECT 135.120 -112.585 135.350 -111.085 ;
        RECT 135.610 -112.765 135.840 -111.085 ;
        RECT 136.100 -112.585 136.330 -108.400 ;
        RECT 138.165 -109.175 138.395 -108.395 ;
        RECT 139.145 -109.165 139.375 -108.395 ;
        RECT 138.655 -109.175 139.865 -109.165 ;
        RECT 140.125 -109.175 140.355 -108.395 ;
        RECT 138.165 -109.405 141.350 -109.175 ;
        RECT 138.165 -110.050 138.395 -109.550 ;
        RECT 138.655 -110.050 138.885 -109.405 ;
        RECT 139.145 -110.050 139.375 -109.550 ;
        RECT 139.635 -110.050 139.865 -109.405 ;
        RECT 142.355 -110.955 142.585 -107.955 ;
        RECT 143.410 -110.955 143.640 -107.955 ;
        RECT 143.900 -110.955 144.130 -107.955 ;
        RECT 144.390 -110.955 144.620 -107.955 ;
        RECT 145.450 -110.955 145.680 -107.955 ;
        RECT 136.590 -112.765 136.820 -111.085 ;
        RECT 146.605 -111.610 147.130 -111.250 ;
        RECT 146.635 -112.025 146.960 -111.610 ;
        RECT 141.860 -112.350 146.960 -112.025 ;
        RECT 134.625 -113.000 136.820 -112.765 ;
        RECT 142.355 -114.015 142.585 -112.515 ;
        RECT 142.845 -114.015 143.075 -112.515 ;
        RECT 143.335 -114.015 143.565 -112.515 ;
        RECT 144.545 -114.015 144.775 -112.515 ;
        RECT 145.035 -114.015 145.265 -112.515 ;
        RECT 146.200 -114.555 146.765 -114.550 ;
        RECT 148.070 -114.555 148.635 -103.575 ;
        RECT 152.315 -109.745 152.545 -107.245 ;
        RECT 153.660 -109.745 153.890 -107.245 ;
        RECT 154.150 -109.745 154.380 -107.245 ;
        RECT 154.640 -109.745 154.870 -107.245 ;
        RECT 155.290 -109.745 155.520 -107.245 ;
        RECT 156.920 -109.745 157.150 -107.245 ;
        RECT 158.060 -108.745 158.290 -107.245 ;
        RECT 151.160 -110.545 151.850 -110.525 ;
        RECT 155.190 -110.545 155.880 -110.525 ;
        RECT 157.115 -110.545 157.385 -110.180 ;
        RECT 151.160 -110.765 157.385 -110.545 ;
        RECT 151.160 -110.795 151.850 -110.765 ;
        RECT 155.190 -110.795 155.880 -110.765 ;
        RECT 157.115 -110.870 157.385 -110.765 ;
        RECT 157.975 -110.945 158.305 -110.885 ;
        RECT 160.975 -110.945 161.820 -99.710 ;
        RECT 167.355 -100.320 168.600 -94.150 ;
        RECT 169.410 -99.450 204.820 -98.495 ;
        RECT 166.900 -101.000 168.685 -100.320 ;
        RECT 166.900 -101.270 168.715 -101.000 ;
        RECT 166.900 -101.655 168.685 -101.270 ;
        RECT 150.355 -112.480 150.870 -112.025 ;
        RECT 145.250 -115.120 148.635 -114.555 ;
        RECT 129.495 -118.380 131.245 -117.950 ;
        RECT 139.580 -118.300 141.775 -118.065 ;
        RECT 129.495 -118.650 138.135 -118.380 ;
        RECT 139.580 -118.485 139.815 -118.300 ;
        RECT 129.495 -118.795 131.245 -118.650 ;
        RECT 133.780 -120.850 134.430 -120.100 ;
        RECT 135.210 -120.370 135.440 -119.370 ;
        RECT 135.700 -120.510 135.930 -119.370 ;
        RECT 136.190 -120.370 136.420 -119.370 ;
        RECT 136.680 -120.510 136.910 -119.370 ;
        RECT 137.865 -120.100 138.135 -118.650 ;
        RECT 139.585 -119.980 139.815 -118.485 ;
        RECT 140.075 -119.980 140.305 -118.480 ;
        RECT 140.565 -119.980 140.795 -118.300 ;
        RECT 137.865 -120.370 139.505 -120.100 ;
        RECT 135.210 -120.740 138.395 -120.510 ;
        RECT 139.235 -120.645 139.505 -120.370 ;
        RECT 134.030 -127.870 134.300 -120.850 ;
        RECT 135.210 -122.020 135.440 -120.740 ;
        RECT 135.700 -120.750 136.910 -120.740 ;
        RECT 136.190 -122.020 136.420 -120.750 ;
        RECT 137.170 -122.020 137.400 -120.740 ;
        RECT 139.105 -120.935 139.900 -120.645 ;
        RECT 140.075 -122.665 140.305 -121.165 ;
        RECT 141.055 -122.665 141.285 -118.480 ;
        RECT 141.545 -119.980 141.775 -118.300 ;
        RECT 146.200 -120.275 146.765 -115.120 ;
        RECT 150.415 -115.645 150.810 -112.480 ;
        RECT 151.825 -113.725 152.055 -112.225 ;
        RECT 152.315 -113.725 152.545 -112.225 ;
        RECT 154.175 -113.725 154.405 -111.225 ;
        RECT 154.665 -113.725 154.895 -111.225 ;
        RECT 155.290 -113.725 155.520 -111.225 ;
        RECT 155.780 -113.725 156.010 -111.225 ;
        RECT 156.430 -113.725 156.660 -111.225 ;
        RECT 156.920 -113.725 157.150 -111.225 ;
        RECT 157.410 -113.725 157.640 -111.225 ;
        RECT 157.975 -111.255 166.085 -110.945 ;
        RECT 157.975 -111.300 158.305 -111.255 ;
        RECT 158.060 -113.725 158.290 -112.225 ;
        RECT 158.550 -113.725 158.780 -112.225 ;
        RECT 147.915 -116.040 150.810 -115.645 ;
        RECT 147.915 -117.815 148.310 -116.040 ;
        RECT 147.785 -118.300 148.365 -117.815 ;
        RECT 157.920 -118.455 160.115 -118.220 ;
        RECT 150.930 -118.535 151.415 -118.505 ;
        RECT 150.930 -118.805 156.475 -118.535 ;
        RECT 157.920 -118.640 158.155 -118.455 ;
        RECT 150.930 -118.835 151.415 -118.805 ;
        RECT 145.055 -120.840 148.595 -120.275 ;
        RECT 143.120 -121.515 143.350 -121.015 ;
        RECT 143.610 -121.660 143.840 -121.015 ;
        RECT 144.100 -121.515 144.330 -121.015 ;
        RECT 144.590 -121.660 144.820 -121.015 ;
        RECT 143.120 -121.890 146.305 -121.660 ;
        RECT 143.120 -122.670 143.350 -121.890 ;
        RECT 143.610 -121.900 144.820 -121.890 ;
        RECT 144.100 -122.670 144.330 -121.900 ;
        RECT 145.080 -122.670 145.310 -121.890 ;
        RECT 135.080 -127.165 135.310 -125.665 ;
        RECT 133.315 -128.140 134.300 -127.870 ;
        RECT 134.590 -129.845 134.820 -128.350 ;
        RECT 134.585 -130.030 134.820 -129.845 ;
        RECT 135.080 -129.850 135.310 -128.350 ;
        RECT 135.570 -130.030 135.800 -128.350 ;
        RECT 136.060 -129.850 136.290 -125.665 ;
        RECT 138.125 -126.440 138.355 -125.660 ;
        RECT 139.105 -126.430 139.335 -125.660 ;
        RECT 138.615 -126.440 139.825 -126.430 ;
        RECT 140.085 -126.440 140.315 -125.660 ;
        RECT 138.125 -126.670 141.310 -126.440 ;
        RECT 138.125 -127.315 138.355 -126.815 ;
        RECT 138.615 -127.315 138.845 -126.670 ;
        RECT 139.105 -127.315 139.335 -126.815 ;
        RECT 139.595 -127.315 139.825 -126.670 ;
        RECT 142.315 -128.220 142.545 -125.220 ;
        RECT 143.370 -128.220 143.600 -125.220 ;
        RECT 143.860 -128.220 144.090 -125.220 ;
        RECT 144.350 -128.220 144.580 -125.220 ;
        RECT 145.410 -128.220 145.640 -125.220 ;
        RECT 136.550 -130.030 136.780 -128.350 ;
        RECT 146.565 -128.875 147.090 -128.515 ;
        RECT 146.595 -129.290 146.920 -128.875 ;
        RECT 141.820 -129.615 146.920 -129.290 ;
        RECT 134.585 -130.265 136.780 -130.030 ;
        RECT 142.315 -131.280 142.545 -129.780 ;
        RECT 142.805 -131.280 143.035 -129.780 ;
        RECT 143.295 -131.280 143.525 -129.780 ;
        RECT 144.505 -131.280 144.735 -129.780 ;
        RECT 144.995 -131.280 145.225 -129.780 ;
        RECT 148.030 -131.820 148.595 -120.840 ;
        RECT 152.120 -121.005 152.770 -120.255 ;
        RECT 153.550 -120.525 153.780 -119.525 ;
        RECT 154.040 -120.665 154.270 -119.525 ;
        RECT 154.530 -120.525 154.760 -119.525 ;
        RECT 155.020 -120.665 155.250 -119.525 ;
        RECT 156.205 -120.255 156.475 -118.805 ;
        RECT 157.925 -120.135 158.155 -118.640 ;
        RECT 158.415 -120.135 158.645 -118.635 ;
        RECT 158.905 -120.135 159.135 -118.455 ;
        RECT 156.205 -120.525 157.845 -120.255 ;
        RECT 153.550 -120.895 156.735 -120.665 ;
        RECT 157.575 -120.800 157.845 -120.525 ;
        RECT 152.370 -128.025 152.640 -121.005 ;
        RECT 153.550 -122.175 153.780 -120.895 ;
        RECT 154.040 -120.905 155.250 -120.895 ;
        RECT 154.530 -122.175 154.760 -120.905 ;
        RECT 155.510 -122.175 155.740 -120.895 ;
        RECT 157.445 -121.090 158.240 -120.800 ;
        RECT 158.415 -122.820 158.645 -121.320 ;
        RECT 159.395 -122.820 159.625 -118.635 ;
        RECT 159.885 -120.135 160.115 -118.455 ;
        RECT 163.395 -120.995 166.935 -120.430 ;
        RECT 161.460 -121.670 161.690 -121.170 ;
        RECT 161.950 -121.815 162.180 -121.170 ;
        RECT 162.440 -121.670 162.670 -121.170 ;
        RECT 162.930 -121.815 163.160 -121.170 ;
        RECT 161.460 -122.045 164.645 -121.815 ;
        RECT 161.460 -122.825 161.690 -122.045 ;
        RECT 161.950 -122.055 163.160 -122.045 ;
        RECT 162.440 -122.825 162.670 -122.055 ;
        RECT 163.420 -122.825 163.650 -122.045 ;
        RECT 153.420 -127.320 153.650 -125.820 ;
        RECT 151.655 -128.295 152.640 -128.025 ;
        RECT 152.930 -130.000 153.160 -128.505 ;
        RECT 152.925 -130.185 153.160 -130.000 ;
        RECT 153.420 -130.005 153.650 -128.505 ;
        RECT 153.910 -130.185 154.140 -128.505 ;
        RECT 154.400 -130.005 154.630 -125.820 ;
        RECT 156.465 -126.595 156.695 -125.815 ;
        RECT 157.445 -126.585 157.675 -125.815 ;
        RECT 156.955 -126.595 158.165 -126.585 ;
        RECT 158.425 -126.595 158.655 -125.815 ;
        RECT 156.465 -126.825 159.650 -126.595 ;
        RECT 156.465 -127.470 156.695 -126.970 ;
        RECT 156.955 -127.470 157.185 -126.825 ;
        RECT 157.445 -127.470 157.675 -126.970 ;
        RECT 157.935 -127.470 158.165 -126.825 ;
        RECT 160.655 -128.375 160.885 -125.375 ;
        RECT 161.710 -128.375 161.940 -125.375 ;
        RECT 162.200 -128.375 162.430 -125.375 ;
        RECT 162.690 -128.375 162.920 -125.375 ;
        RECT 163.750 -128.375 163.980 -125.375 ;
        RECT 154.890 -130.185 155.120 -128.505 ;
        RECT 164.905 -129.030 165.430 -128.670 ;
        RECT 164.935 -129.445 165.260 -129.030 ;
        RECT 160.160 -129.770 165.260 -129.445 ;
        RECT 152.925 -130.420 155.120 -130.185 ;
        RECT 160.655 -131.435 160.885 -129.935 ;
        RECT 161.145 -131.435 161.375 -129.935 ;
        RECT 161.635 -131.435 161.865 -129.935 ;
        RECT 162.845 -131.435 163.075 -129.935 ;
        RECT 163.335 -131.435 163.565 -129.935 ;
        RECT 145.210 -131.975 148.595 -131.820 ;
        RECT 166.370 -131.975 166.935 -120.995 ;
        RECT 167.355 -129.100 168.600 -101.655 ;
        RECT 169.410 -118.020 170.365 -99.450 ;
        RECT 172.790 -101.170 174.575 -100.490 ;
        RECT 181.820 -101.090 184.015 -100.855 ;
        RECT 172.790 -101.440 180.375 -101.170 ;
        RECT 181.820 -101.275 182.055 -101.090 ;
        RECT 172.790 -101.825 174.575 -101.440 ;
        RECT 176.020 -103.640 176.670 -102.890 ;
        RECT 177.450 -103.160 177.680 -102.160 ;
        RECT 177.940 -103.300 178.170 -102.160 ;
        RECT 178.430 -103.160 178.660 -102.160 ;
        RECT 178.920 -103.300 179.150 -102.160 ;
        RECT 180.105 -102.890 180.375 -101.440 ;
        RECT 181.825 -102.770 182.055 -101.275 ;
        RECT 182.315 -102.770 182.545 -101.270 ;
        RECT 182.805 -102.770 183.035 -101.090 ;
        RECT 180.105 -103.160 181.745 -102.890 ;
        RECT 177.450 -103.530 180.635 -103.300 ;
        RECT 181.475 -103.435 181.745 -103.160 ;
        RECT 176.270 -110.660 176.540 -103.640 ;
        RECT 177.450 -104.810 177.680 -103.530 ;
        RECT 177.940 -103.540 179.150 -103.530 ;
        RECT 178.430 -104.810 178.660 -103.540 ;
        RECT 179.410 -104.810 179.640 -103.530 ;
        RECT 181.345 -103.725 182.140 -103.435 ;
        RECT 182.315 -105.455 182.545 -103.955 ;
        RECT 183.295 -105.455 183.525 -101.270 ;
        RECT 183.785 -102.770 184.015 -101.090 ;
        RECT 187.295 -103.630 190.835 -103.065 ;
        RECT 185.360 -104.305 185.590 -103.805 ;
        RECT 185.850 -104.450 186.080 -103.805 ;
        RECT 186.340 -104.305 186.570 -103.805 ;
        RECT 186.830 -104.450 187.060 -103.805 ;
        RECT 185.360 -104.680 188.545 -104.450 ;
        RECT 185.360 -105.460 185.590 -104.680 ;
        RECT 185.850 -104.690 187.060 -104.680 ;
        RECT 186.340 -105.460 186.570 -104.690 ;
        RECT 187.320 -105.460 187.550 -104.680 ;
        RECT 177.320 -109.955 177.550 -108.455 ;
        RECT 175.555 -110.930 176.540 -110.660 ;
        RECT 176.830 -112.635 177.060 -111.140 ;
        RECT 176.825 -112.820 177.060 -112.635 ;
        RECT 177.320 -112.640 177.550 -111.140 ;
        RECT 177.810 -112.820 178.040 -111.140 ;
        RECT 178.300 -112.640 178.530 -108.455 ;
        RECT 180.365 -109.230 180.595 -108.450 ;
        RECT 181.345 -109.220 181.575 -108.450 ;
        RECT 180.855 -109.230 182.065 -109.220 ;
        RECT 182.325 -109.230 182.555 -108.450 ;
        RECT 180.365 -109.460 183.550 -109.230 ;
        RECT 180.365 -110.105 180.595 -109.605 ;
        RECT 180.855 -110.105 181.085 -109.460 ;
        RECT 181.345 -110.105 181.575 -109.605 ;
        RECT 181.835 -110.105 182.065 -109.460 ;
        RECT 184.555 -111.010 184.785 -108.010 ;
        RECT 185.610 -111.010 185.840 -108.010 ;
        RECT 186.100 -111.010 186.330 -108.010 ;
        RECT 186.590 -111.010 186.820 -108.010 ;
        RECT 187.650 -111.010 187.880 -108.010 ;
        RECT 178.790 -112.820 179.020 -111.140 ;
        RECT 188.805 -111.665 189.330 -111.305 ;
        RECT 188.835 -112.080 189.160 -111.665 ;
        RECT 184.060 -112.405 189.160 -112.080 ;
        RECT 176.825 -113.055 179.020 -112.820 ;
        RECT 184.555 -114.070 184.785 -112.570 ;
        RECT 185.045 -114.070 185.275 -112.570 ;
        RECT 185.535 -114.070 185.765 -112.570 ;
        RECT 186.745 -114.070 186.975 -112.570 ;
        RECT 187.235 -114.070 187.465 -112.570 ;
        RECT 188.400 -114.610 188.965 -114.605 ;
        RECT 190.270 -114.610 190.835 -103.630 ;
        RECT 194.515 -109.800 194.745 -107.300 ;
        RECT 195.860 -109.800 196.090 -107.300 ;
        RECT 196.350 -109.800 196.580 -107.300 ;
        RECT 196.840 -109.800 197.070 -107.300 ;
        RECT 197.490 -109.800 197.720 -107.300 ;
        RECT 199.120 -109.800 199.350 -107.300 ;
        RECT 200.260 -108.800 200.490 -107.300 ;
        RECT 193.360 -110.600 194.050 -110.580 ;
        RECT 197.390 -110.600 198.080 -110.580 ;
        RECT 199.315 -110.600 199.585 -110.235 ;
        RECT 193.360 -110.820 199.585 -110.600 ;
        RECT 193.360 -110.850 194.050 -110.820 ;
        RECT 197.390 -110.850 198.080 -110.820 ;
        RECT 199.315 -110.925 199.585 -110.820 ;
        RECT 200.175 -111.000 200.505 -110.940 ;
        RECT 203.740 -111.000 204.820 -99.450 ;
        RECT 192.555 -112.535 193.070 -112.080 ;
        RECT 187.450 -115.175 190.835 -114.610 ;
        RECT 169.410 -118.435 173.660 -118.020 ;
        RECT 181.780 -118.355 183.975 -118.120 ;
        RECT 169.410 -118.705 180.335 -118.435 ;
        RECT 181.780 -118.540 182.015 -118.355 ;
        RECT 169.410 -118.975 173.660 -118.705 ;
        RECT 175.980 -120.905 176.630 -120.155 ;
        RECT 177.410 -120.425 177.640 -119.425 ;
        RECT 177.900 -120.565 178.130 -119.425 ;
        RECT 178.390 -120.425 178.620 -119.425 ;
        RECT 178.880 -120.565 179.110 -119.425 ;
        RECT 180.065 -120.155 180.335 -118.705 ;
        RECT 181.785 -120.035 182.015 -118.540 ;
        RECT 182.275 -120.035 182.505 -118.535 ;
        RECT 182.765 -120.035 182.995 -118.355 ;
        RECT 180.065 -120.425 181.705 -120.155 ;
        RECT 177.410 -120.795 180.595 -120.565 ;
        RECT 181.435 -120.700 181.705 -120.425 ;
        RECT 176.230 -127.925 176.500 -120.905 ;
        RECT 177.410 -122.075 177.640 -120.795 ;
        RECT 177.900 -120.805 179.110 -120.795 ;
        RECT 178.390 -122.075 178.620 -120.805 ;
        RECT 179.370 -122.075 179.600 -120.795 ;
        RECT 181.305 -120.990 182.100 -120.700 ;
        RECT 182.275 -122.720 182.505 -121.220 ;
        RECT 183.255 -122.720 183.485 -118.535 ;
        RECT 183.745 -120.035 183.975 -118.355 ;
        RECT 188.400 -120.330 188.965 -115.175 ;
        RECT 192.615 -115.700 193.010 -112.535 ;
        RECT 194.025 -113.780 194.255 -112.280 ;
        RECT 194.515 -113.780 194.745 -112.280 ;
        RECT 196.375 -113.780 196.605 -111.280 ;
        RECT 196.865 -113.780 197.095 -111.280 ;
        RECT 197.490 -113.780 197.720 -111.280 ;
        RECT 197.980 -113.780 198.210 -111.280 ;
        RECT 198.630 -113.780 198.860 -111.280 ;
        RECT 199.120 -113.780 199.350 -111.280 ;
        RECT 199.610 -113.780 199.840 -111.280 ;
        RECT 200.175 -111.310 208.285 -111.000 ;
        RECT 200.175 -111.355 200.505 -111.310 ;
        RECT 200.260 -113.780 200.490 -112.280 ;
        RECT 200.750 -113.780 200.980 -112.280 ;
        RECT 190.115 -116.095 193.010 -115.700 ;
        RECT 190.115 -117.870 190.510 -116.095 ;
        RECT 189.985 -118.355 190.565 -117.870 ;
        RECT 200.120 -118.510 202.315 -118.275 ;
        RECT 193.130 -118.590 193.615 -118.560 ;
        RECT 193.130 -118.860 198.675 -118.590 ;
        RECT 200.120 -118.695 200.355 -118.510 ;
        RECT 193.130 -118.890 193.615 -118.860 ;
        RECT 187.255 -120.895 190.795 -120.330 ;
        RECT 185.320 -121.570 185.550 -121.070 ;
        RECT 185.810 -121.715 186.040 -121.070 ;
        RECT 186.300 -121.570 186.530 -121.070 ;
        RECT 186.790 -121.715 187.020 -121.070 ;
        RECT 185.320 -121.945 188.505 -121.715 ;
        RECT 185.320 -122.725 185.550 -121.945 ;
        RECT 185.810 -121.955 187.020 -121.945 ;
        RECT 186.300 -122.725 186.530 -121.955 ;
        RECT 187.280 -122.725 187.510 -121.945 ;
        RECT 177.280 -127.220 177.510 -125.720 ;
        RECT 175.515 -128.195 176.500 -127.925 ;
        RECT 167.435 -129.945 168.550 -129.100 ;
        RECT 176.790 -129.900 177.020 -128.405 ;
        RECT 176.785 -130.085 177.020 -129.900 ;
        RECT 177.280 -129.905 177.510 -128.405 ;
        RECT 177.770 -130.085 178.000 -128.405 ;
        RECT 178.260 -129.905 178.490 -125.720 ;
        RECT 180.325 -126.495 180.555 -125.715 ;
        RECT 181.305 -126.485 181.535 -125.715 ;
        RECT 180.815 -126.495 182.025 -126.485 ;
        RECT 182.285 -126.495 182.515 -125.715 ;
        RECT 180.325 -126.725 183.510 -126.495 ;
        RECT 180.325 -127.370 180.555 -126.870 ;
        RECT 180.815 -127.370 181.045 -126.725 ;
        RECT 181.305 -127.370 181.535 -126.870 ;
        RECT 181.795 -127.370 182.025 -126.725 ;
        RECT 184.515 -128.275 184.745 -125.275 ;
        RECT 185.570 -128.275 185.800 -125.275 ;
        RECT 186.060 -128.275 186.290 -125.275 ;
        RECT 186.550 -128.275 186.780 -125.275 ;
        RECT 187.610 -128.275 187.840 -125.275 ;
        RECT 178.750 -130.085 178.980 -128.405 ;
        RECT 188.765 -128.930 189.290 -128.570 ;
        RECT 188.795 -129.345 189.120 -128.930 ;
        RECT 184.020 -129.670 189.120 -129.345 ;
        RECT 176.785 -130.320 178.980 -130.085 ;
        RECT 184.515 -131.335 184.745 -129.835 ;
        RECT 185.005 -131.335 185.235 -129.835 ;
        RECT 185.495 -131.335 185.725 -129.835 ;
        RECT 186.705 -131.335 186.935 -129.835 ;
        RECT 187.195 -131.335 187.425 -129.835 ;
        RECT 190.230 -131.875 190.795 -120.895 ;
        RECT 194.320 -121.060 194.970 -120.310 ;
        RECT 195.750 -120.580 195.980 -119.580 ;
        RECT 196.240 -120.720 196.470 -119.580 ;
        RECT 196.730 -120.580 196.960 -119.580 ;
        RECT 197.220 -120.720 197.450 -119.580 ;
        RECT 198.405 -120.310 198.675 -118.860 ;
        RECT 200.125 -120.190 200.355 -118.695 ;
        RECT 200.615 -120.190 200.845 -118.690 ;
        RECT 201.105 -120.190 201.335 -118.510 ;
        RECT 198.405 -120.580 200.045 -120.310 ;
        RECT 195.750 -120.950 198.935 -120.720 ;
        RECT 199.775 -120.855 200.045 -120.580 ;
        RECT 194.570 -128.080 194.840 -121.060 ;
        RECT 195.750 -122.230 195.980 -120.950 ;
        RECT 196.240 -120.960 197.450 -120.950 ;
        RECT 196.730 -122.230 196.960 -120.960 ;
        RECT 197.710 -122.230 197.940 -120.950 ;
        RECT 199.645 -121.145 200.440 -120.855 ;
        RECT 200.615 -122.875 200.845 -121.375 ;
        RECT 201.595 -122.875 201.825 -118.690 ;
        RECT 202.085 -120.190 202.315 -118.510 ;
        RECT 205.595 -121.050 209.135 -120.485 ;
        RECT 203.660 -121.725 203.890 -121.225 ;
        RECT 204.150 -121.870 204.380 -121.225 ;
        RECT 204.640 -121.725 204.870 -121.225 ;
        RECT 205.130 -121.870 205.360 -121.225 ;
        RECT 203.660 -122.100 206.845 -121.870 ;
        RECT 203.660 -122.880 203.890 -122.100 ;
        RECT 204.150 -122.110 205.360 -122.100 ;
        RECT 204.640 -122.880 204.870 -122.110 ;
        RECT 205.620 -122.880 205.850 -122.100 ;
        RECT 195.620 -127.375 195.850 -125.875 ;
        RECT 193.855 -128.350 194.840 -128.080 ;
        RECT 195.130 -130.055 195.360 -128.560 ;
        RECT 195.125 -130.240 195.360 -130.055 ;
        RECT 195.620 -130.060 195.850 -128.560 ;
        RECT 196.110 -130.240 196.340 -128.560 ;
        RECT 196.600 -130.060 196.830 -125.875 ;
        RECT 198.665 -126.650 198.895 -125.870 ;
        RECT 199.645 -126.640 199.875 -125.870 ;
        RECT 199.155 -126.650 200.365 -126.640 ;
        RECT 200.625 -126.650 200.855 -125.870 ;
        RECT 198.665 -126.880 201.850 -126.650 ;
        RECT 198.665 -127.525 198.895 -127.025 ;
        RECT 199.155 -127.525 199.385 -126.880 ;
        RECT 199.645 -127.525 199.875 -127.025 ;
        RECT 200.135 -127.525 200.365 -126.880 ;
        RECT 202.855 -128.430 203.085 -125.430 ;
        RECT 203.910 -128.430 204.140 -125.430 ;
        RECT 204.400 -128.430 204.630 -125.430 ;
        RECT 204.890 -128.430 205.120 -125.430 ;
        RECT 205.950 -128.430 206.180 -125.430 ;
        RECT 197.090 -130.240 197.320 -128.560 ;
        RECT 207.105 -129.085 207.630 -128.725 ;
        RECT 207.135 -129.500 207.460 -129.085 ;
        RECT 202.360 -129.825 207.460 -129.500 ;
        RECT 195.125 -130.475 197.320 -130.240 ;
        RECT 202.855 -131.490 203.085 -129.990 ;
        RECT 203.345 -131.490 203.575 -129.990 ;
        RECT 203.835 -131.490 204.065 -129.990 ;
        RECT 205.045 -131.490 205.275 -129.990 ;
        RECT 205.535 -131.490 205.765 -129.990 ;
        RECT 145.210 -132.385 166.935 -131.975 ;
        RECT 145.230 -132.540 166.935 -132.385 ;
        RECT 187.410 -132.030 190.795 -131.875 ;
        RECT 208.570 -132.030 209.135 -121.050 ;
        RECT 209.680 -128.785 211.005 -92.120 ;
        RECT 211.890 -99.415 251.695 -98.405 ;
        RECT 211.890 -118.365 212.900 -99.415 ;
        RECT 217.310 -101.365 218.795 -100.935 ;
        RECT 226.135 -101.285 228.330 -101.050 ;
        RECT 217.310 -101.635 224.690 -101.365 ;
        RECT 226.135 -101.470 226.370 -101.285 ;
        RECT 217.310 -102.045 218.795 -101.635 ;
        RECT 220.335 -103.835 220.985 -103.085 ;
        RECT 221.765 -103.355 221.995 -102.355 ;
        RECT 222.255 -103.495 222.485 -102.355 ;
        RECT 222.745 -103.355 222.975 -102.355 ;
        RECT 223.235 -103.495 223.465 -102.355 ;
        RECT 224.420 -103.085 224.690 -101.635 ;
        RECT 226.140 -102.965 226.370 -101.470 ;
        RECT 226.630 -102.965 226.860 -101.465 ;
        RECT 227.120 -102.965 227.350 -101.285 ;
        RECT 224.420 -103.355 226.060 -103.085 ;
        RECT 221.765 -103.725 224.950 -103.495 ;
        RECT 225.790 -103.630 226.060 -103.355 ;
        RECT 220.585 -110.855 220.855 -103.835 ;
        RECT 221.765 -105.005 221.995 -103.725 ;
        RECT 222.255 -103.735 223.465 -103.725 ;
        RECT 222.745 -105.005 222.975 -103.735 ;
        RECT 223.725 -105.005 223.955 -103.725 ;
        RECT 225.660 -103.920 226.455 -103.630 ;
        RECT 226.630 -105.650 226.860 -104.150 ;
        RECT 227.610 -105.650 227.840 -101.465 ;
        RECT 228.100 -102.965 228.330 -101.285 ;
        RECT 231.610 -103.825 235.150 -103.260 ;
        RECT 229.675 -104.500 229.905 -104.000 ;
        RECT 230.165 -104.645 230.395 -104.000 ;
        RECT 230.655 -104.500 230.885 -104.000 ;
        RECT 231.145 -104.645 231.375 -104.000 ;
        RECT 229.675 -104.875 232.860 -104.645 ;
        RECT 229.675 -105.655 229.905 -104.875 ;
        RECT 230.165 -104.885 231.375 -104.875 ;
        RECT 230.655 -105.655 230.885 -104.885 ;
        RECT 231.635 -105.655 231.865 -104.875 ;
        RECT 221.635 -110.150 221.865 -108.650 ;
        RECT 219.870 -111.125 220.855 -110.855 ;
        RECT 221.145 -112.830 221.375 -111.335 ;
        RECT 221.140 -113.015 221.375 -112.830 ;
        RECT 221.635 -112.835 221.865 -111.335 ;
        RECT 222.125 -113.015 222.355 -111.335 ;
        RECT 222.615 -112.835 222.845 -108.650 ;
        RECT 224.680 -109.425 224.910 -108.645 ;
        RECT 225.660 -109.415 225.890 -108.645 ;
        RECT 225.170 -109.425 226.380 -109.415 ;
        RECT 226.640 -109.425 226.870 -108.645 ;
        RECT 224.680 -109.655 227.865 -109.425 ;
        RECT 224.680 -110.300 224.910 -109.800 ;
        RECT 225.170 -110.300 225.400 -109.655 ;
        RECT 225.660 -110.300 225.890 -109.800 ;
        RECT 226.150 -110.300 226.380 -109.655 ;
        RECT 228.870 -111.205 229.100 -108.205 ;
        RECT 229.925 -111.205 230.155 -108.205 ;
        RECT 230.415 -111.205 230.645 -108.205 ;
        RECT 230.905 -111.205 231.135 -108.205 ;
        RECT 231.965 -111.205 232.195 -108.205 ;
        RECT 223.105 -113.015 223.335 -111.335 ;
        RECT 233.120 -111.860 233.645 -111.500 ;
        RECT 233.150 -112.275 233.475 -111.860 ;
        RECT 228.375 -112.600 233.475 -112.275 ;
        RECT 221.140 -113.250 223.335 -113.015 ;
        RECT 228.870 -114.265 229.100 -112.765 ;
        RECT 229.360 -114.265 229.590 -112.765 ;
        RECT 229.850 -114.265 230.080 -112.765 ;
        RECT 231.060 -114.265 231.290 -112.765 ;
        RECT 231.550 -114.265 231.780 -112.765 ;
        RECT 232.715 -114.805 233.280 -114.800 ;
        RECT 234.585 -114.805 235.150 -103.825 ;
        RECT 238.830 -109.995 239.060 -107.495 ;
        RECT 240.175 -109.995 240.405 -107.495 ;
        RECT 240.665 -109.995 240.895 -107.495 ;
        RECT 241.155 -109.995 241.385 -107.495 ;
        RECT 241.805 -109.995 242.035 -107.495 ;
        RECT 243.435 -109.995 243.665 -107.495 ;
        RECT 244.575 -108.995 244.805 -107.495 ;
        RECT 237.675 -110.795 238.365 -110.775 ;
        RECT 241.705 -110.795 242.395 -110.775 ;
        RECT 243.630 -110.795 243.900 -110.430 ;
        RECT 237.675 -111.015 243.900 -110.795 ;
        RECT 237.675 -111.045 238.365 -111.015 ;
        RECT 241.705 -111.045 242.395 -111.015 ;
        RECT 243.630 -111.120 243.900 -111.015 ;
        RECT 244.490 -111.195 244.820 -111.135 ;
        RECT 250.685 -111.195 251.695 -99.415 ;
        RECT 236.870 -112.730 237.385 -112.275 ;
        RECT 231.765 -115.370 235.150 -114.805 ;
        RECT 211.890 -118.630 218.540 -118.365 ;
        RECT 226.095 -118.550 228.290 -118.315 ;
        RECT 211.890 -118.900 224.650 -118.630 ;
        RECT 226.095 -118.735 226.330 -118.550 ;
        RECT 211.890 -119.375 218.540 -118.900 ;
        RECT 220.295 -121.100 220.945 -120.350 ;
        RECT 221.725 -120.620 221.955 -119.620 ;
        RECT 222.215 -120.760 222.445 -119.620 ;
        RECT 222.705 -120.620 222.935 -119.620 ;
        RECT 223.195 -120.760 223.425 -119.620 ;
        RECT 224.380 -120.350 224.650 -118.900 ;
        RECT 226.100 -120.230 226.330 -118.735 ;
        RECT 226.590 -120.230 226.820 -118.730 ;
        RECT 227.080 -120.230 227.310 -118.550 ;
        RECT 224.380 -120.620 226.020 -120.350 ;
        RECT 221.725 -120.990 224.910 -120.760 ;
        RECT 225.750 -120.895 226.020 -120.620 ;
        RECT 220.545 -128.120 220.815 -121.100 ;
        RECT 221.725 -122.270 221.955 -120.990 ;
        RECT 222.215 -121.000 223.425 -120.990 ;
        RECT 222.705 -122.270 222.935 -121.000 ;
        RECT 223.685 -122.270 223.915 -120.990 ;
        RECT 225.620 -121.185 226.415 -120.895 ;
        RECT 226.590 -122.915 226.820 -121.415 ;
        RECT 227.570 -122.915 227.800 -118.730 ;
        RECT 228.060 -120.230 228.290 -118.550 ;
        RECT 232.715 -120.525 233.280 -115.370 ;
        RECT 236.930 -115.895 237.325 -112.730 ;
        RECT 238.340 -113.975 238.570 -112.475 ;
        RECT 238.830 -113.975 239.060 -112.475 ;
        RECT 240.690 -113.975 240.920 -111.475 ;
        RECT 241.180 -113.975 241.410 -111.475 ;
        RECT 241.805 -113.975 242.035 -111.475 ;
        RECT 242.295 -113.975 242.525 -111.475 ;
        RECT 242.945 -113.975 243.175 -111.475 ;
        RECT 243.435 -113.975 243.665 -111.475 ;
        RECT 243.925 -113.975 244.155 -111.475 ;
        RECT 244.490 -111.505 252.600 -111.195 ;
        RECT 244.490 -111.550 244.820 -111.505 ;
        RECT 244.575 -113.975 244.805 -112.475 ;
        RECT 245.065 -113.975 245.295 -112.475 ;
        RECT 234.430 -116.290 237.325 -115.895 ;
        RECT 234.430 -118.065 234.825 -116.290 ;
        RECT 234.300 -118.550 234.880 -118.065 ;
        RECT 244.435 -118.705 246.630 -118.470 ;
        RECT 237.445 -118.785 237.930 -118.755 ;
        RECT 237.445 -119.055 242.990 -118.785 ;
        RECT 244.435 -118.890 244.670 -118.705 ;
        RECT 237.445 -119.085 237.930 -119.055 ;
        RECT 231.570 -121.090 235.110 -120.525 ;
        RECT 229.635 -121.765 229.865 -121.265 ;
        RECT 230.125 -121.910 230.355 -121.265 ;
        RECT 230.615 -121.765 230.845 -121.265 ;
        RECT 231.105 -121.910 231.335 -121.265 ;
        RECT 229.635 -122.140 232.820 -121.910 ;
        RECT 229.635 -122.920 229.865 -122.140 ;
        RECT 230.125 -122.150 231.335 -122.140 ;
        RECT 230.615 -122.920 230.845 -122.150 ;
        RECT 231.595 -122.920 231.825 -122.140 ;
        RECT 221.595 -127.415 221.825 -125.915 ;
        RECT 219.830 -128.390 220.815 -128.120 ;
        RECT 209.680 -130.440 211.365 -128.785 ;
        RECT 221.105 -130.095 221.335 -128.600 ;
        RECT 221.100 -130.280 221.335 -130.095 ;
        RECT 221.595 -130.100 221.825 -128.600 ;
        RECT 222.085 -130.280 222.315 -128.600 ;
        RECT 222.575 -130.100 222.805 -125.915 ;
        RECT 224.640 -126.690 224.870 -125.910 ;
        RECT 225.620 -126.680 225.850 -125.910 ;
        RECT 225.130 -126.690 226.340 -126.680 ;
        RECT 226.600 -126.690 226.830 -125.910 ;
        RECT 224.640 -126.920 227.825 -126.690 ;
        RECT 224.640 -127.565 224.870 -127.065 ;
        RECT 225.130 -127.565 225.360 -126.920 ;
        RECT 225.620 -127.565 225.850 -127.065 ;
        RECT 226.110 -127.565 226.340 -126.920 ;
        RECT 228.830 -128.470 229.060 -125.470 ;
        RECT 229.885 -128.470 230.115 -125.470 ;
        RECT 230.375 -128.470 230.605 -125.470 ;
        RECT 230.865 -128.470 231.095 -125.470 ;
        RECT 231.925 -128.470 232.155 -125.470 ;
        RECT 223.065 -130.280 223.295 -128.600 ;
        RECT 233.080 -129.125 233.605 -128.765 ;
        RECT 233.110 -129.540 233.435 -129.125 ;
        RECT 228.335 -129.865 233.435 -129.540 ;
        RECT 221.100 -130.515 223.295 -130.280 ;
        RECT 228.830 -131.530 229.060 -130.030 ;
        RECT 229.320 -131.530 229.550 -130.030 ;
        RECT 229.810 -131.530 230.040 -130.030 ;
        RECT 231.020 -131.530 231.250 -130.030 ;
        RECT 231.510 -131.530 231.740 -130.030 ;
        RECT 187.410 -132.440 209.135 -132.030 ;
        RECT 234.545 -132.070 235.110 -121.090 ;
        RECT 238.635 -121.255 239.285 -120.505 ;
        RECT 240.065 -120.775 240.295 -119.775 ;
        RECT 240.555 -120.915 240.785 -119.775 ;
        RECT 241.045 -120.775 241.275 -119.775 ;
        RECT 241.535 -120.915 241.765 -119.775 ;
        RECT 242.720 -120.505 242.990 -119.055 ;
        RECT 244.440 -120.385 244.670 -118.890 ;
        RECT 244.930 -120.385 245.160 -118.885 ;
        RECT 245.420 -120.385 245.650 -118.705 ;
        RECT 242.720 -120.775 244.360 -120.505 ;
        RECT 240.065 -121.145 243.250 -120.915 ;
        RECT 244.090 -121.050 244.360 -120.775 ;
        RECT 238.885 -128.275 239.155 -121.255 ;
        RECT 240.065 -122.425 240.295 -121.145 ;
        RECT 240.555 -121.155 241.765 -121.145 ;
        RECT 241.045 -122.425 241.275 -121.155 ;
        RECT 242.025 -122.425 242.255 -121.145 ;
        RECT 243.960 -121.340 244.755 -121.050 ;
        RECT 244.930 -123.070 245.160 -121.570 ;
        RECT 245.910 -123.070 246.140 -118.885 ;
        RECT 246.400 -120.385 246.630 -118.705 ;
        RECT 249.910 -121.245 253.450 -120.680 ;
        RECT 247.975 -121.920 248.205 -121.420 ;
        RECT 248.465 -122.065 248.695 -121.420 ;
        RECT 248.955 -121.920 249.185 -121.420 ;
        RECT 249.445 -122.065 249.675 -121.420 ;
        RECT 247.975 -122.295 251.160 -122.065 ;
        RECT 247.975 -123.075 248.205 -122.295 ;
        RECT 248.465 -122.305 249.675 -122.295 ;
        RECT 248.955 -123.075 249.185 -122.305 ;
        RECT 249.935 -123.075 250.165 -122.295 ;
        RECT 239.935 -127.570 240.165 -126.070 ;
        RECT 238.170 -128.545 239.155 -128.275 ;
        RECT 239.445 -130.250 239.675 -128.755 ;
        RECT 239.440 -130.435 239.675 -130.250 ;
        RECT 239.935 -130.255 240.165 -128.755 ;
        RECT 240.425 -130.435 240.655 -128.755 ;
        RECT 240.915 -130.255 241.145 -126.070 ;
        RECT 242.980 -126.845 243.210 -126.065 ;
        RECT 243.960 -126.835 244.190 -126.065 ;
        RECT 243.470 -126.845 244.680 -126.835 ;
        RECT 244.940 -126.845 245.170 -126.065 ;
        RECT 242.980 -127.075 246.165 -126.845 ;
        RECT 242.980 -127.720 243.210 -127.220 ;
        RECT 243.470 -127.720 243.700 -127.075 ;
        RECT 243.960 -127.720 244.190 -127.220 ;
        RECT 244.450 -127.720 244.680 -127.075 ;
        RECT 247.170 -128.625 247.400 -125.625 ;
        RECT 248.225 -128.625 248.455 -125.625 ;
        RECT 248.715 -128.625 248.945 -125.625 ;
        RECT 249.205 -128.625 249.435 -125.625 ;
        RECT 250.265 -128.625 250.495 -125.625 ;
        RECT 241.405 -130.435 241.635 -128.755 ;
        RECT 251.420 -129.280 251.945 -128.920 ;
        RECT 251.450 -129.695 251.775 -129.280 ;
        RECT 246.675 -130.020 251.775 -129.695 ;
        RECT 239.440 -130.670 241.635 -130.435 ;
        RECT 247.170 -131.685 247.400 -130.185 ;
        RECT 247.660 -131.685 247.890 -130.185 ;
        RECT 248.150 -131.685 248.380 -130.185 ;
        RECT 249.360 -131.685 249.590 -130.185 ;
        RECT 249.850 -131.685 250.080 -130.185 ;
        RECT 187.430 -132.595 209.135 -132.440 ;
        RECT 231.725 -132.225 235.110 -132.070 ;
        RECT 252.885 -132.225 253.450 -121.245 ;
        RECT 254.000 -128.090 255.130 -89.720 ;
        RECT 258.285 -99.740 298.215 -98.445 ;
        RECT 258.285 -117.760 259.580 -99.740 ;
        RECT 262.265 -101.195 263.495 -100.715 ;
        RECT 272.125 -101.115 274.320 -100.880 ;
        RECT 262.265 -101.465 270.680 -101.195 ;
        RECT 272.125 -101.300 272.360 -101.115 ;
        RECT 262.265 -101.815 263.495 -101.465 ;
        RECT 266.325 -103.665 266.975 -102.915 ;
        RECT 267.755 -103.185 267.985 -102.185 ;
        RECT 268.245 -103.325 268.475 -102.185 ;
        RECT 268.735 -103.185 268.965 -102.185 ;
        RECT 269.225 -103.325 269.455 -102.185 ;
        RECT 270.410 -102.915 270.680 -101.465 ;
        RECT 272.130 -102.795 272.360 -101.300 ;
        RECT 272.620 -102.795 272.850 -101.295 ;
        RECT 273.110 -102.795 273.340 -101.115 ;
        RECT 270.410 -103.185 272.050 -102.915 ;
        RECT 267.755 -103.555 270.940 -103.325 ;
        RECT 271.780 -103.460 272.050 -103.185 ;
        RECT 266.575 -110.685 266.845 -103.665 ;
        RECT 267.755 -104.835 267.985 -103.555 ;
        RECT 268.245 -103.565 269.455 -103.555 ;
        RECT 268.735 -104.835 268.965 -103.565 ;
        RECT 269.715 -104.835 269.945 -103.555 ;
        RECT 271.650 -103.750 272.445 -103.460 ;
        RECT 272.620 -105.480 272.850 -103.980 ;
        RECT 273.600 -105.480 273.830 -101.295 ;
        RECT 274.090 -102.795 274.320 -101.115 ;
        RECT 277.600 -103.655 281.140 -103.090 ;
        RECT 275.665 -104.330 275.895 -103.830 ;
        RECT 276.155 -104.475 276.385 -103.830 ;
        RECT 276.645 -104.330 276.875 -103.830 ;
        RECT 277.135 -104.475 277.365 -103.830 ;
        RECT 275.665 -104.705 278.850 -104.475 ;
        RECT 275.665 -105.485 275.895 -104.705 ;
        RECT 276.155 -104.715 277.365 -104.705 ;
        RECT 276.645 -105.485 276.875 -104.715 ;
        RECT 277.625 -105.485 277.855 -104.705 ;
        RECT 267.625 -109.980 267.855 -108.480 ;
        RECT 265.860 -110.955 266.845 -110.685 ;
        RECT 267.135 -112.660 267.365 -111.165 ;
        RECT 267.130 -112.845 267.365 -112.660 ;
        RECT 267.625 -112.665 267.855 -111.165 ;
        RECT 268.115 -112.845 268.345 -111.165 ;
        RECT 268.605 -112.665 268.835 -108.480 ;
        RECT 270.670 -109.255 270.900 -108.475 ;
        RECT 271.650 -109.245 271.880 -108.475 ;
        RECT 271.160 -109.255 272.370 -109.245 ;
        RECT 272.630 -109.255 272.860 -108.475 ;
        RECT 270.670 -109.485 273.855 -109.255 ;
        RECT 270.670 -110.130 270.900 -109.630 ;
        RECT 271.160 -110.130 271.390 -109.485 ;
        RECT 271.650 -110.130 271.880 -109.630 ;
        RECT 272.140 -110.130 272.370 -109.485 ;
        RECT 274.860 -111.035 275.090 -108.035 ;
        RECT 275.915 -111.035 276.145 -108.035 ;
        RECT 276.405 -111.035 276.635 -108.035 ;
        RECT 276.895 -111.035 277.125 -108.035 ;
        RECT 277.955 -111.035 278.185 -108.035 ;
        RECT 269.095 -112.845 269.325 -111.165 ;
        RECT 279.110 -111.690 279.635 -111.330 ;
        RECT 279.140 -112.105 279.465 -111.690 ;
        RECT 274.365 -112.430 279.465 -112.105 ;
        RECT 267.130 -113.080 269.325 -112.845 ;
        RECT 274.860 -114.095 275.090 -112.595 ;
        RECT 275.350 -114.095 275.580 -112.595 ;
        RECT 275.840 -114.095 276.070 -112.595 ;
        RECT 277.050 -114.095 277.280 -112.595 ;
        RECT 277.540 -114.095 277.770 -112.595 ;
        RECT 278.705 -114.635 279.270 -114.630 ;
        RECT 280.575 -114.635 281.140 -103.655 ;
        RECT 284.820 -109.825 285.050 -107.325 ;
        RECT 286.165 -109.825 286.395 -107.325 ;
        RECT 286.655 -109.825 286.885 -107.325 ;
        RECT 287.145 -109.825 287.375 -107.325 ;
        RECT 287.795 -109.825 288.025 -107.325 ;
        RECT 289.425 -109.825 289.655 -107.325 ;
        RECT 290.565 -108.825 290.795 -107.325 ;
        RECT 283.665 -110.625 284.355 -110.605 ;
        RECT 287.695 -110.625 288.385 -110.605 ;
        RECT 289.620 -110.625 289.890 -110.260 ;
        RECT 283.665 -110.845 289.890 -110.625 ;
        RECT 283.665 -110.875 284.355 -110.845 ;
        RECT 287.695 -110.875 288.385 -110.845 ;
        RECT 289.620 -110.950 289.890 -110.845 ;
        RECT 290.480 -111.025 290.810 -110.965 ;
        RECT 296.920 -111.025 298.215 -99.740 ;
        RECT 299.970 -100.025 301.075 -86.935 ;
        RECT 302.230 -99.840 342.150 -98.650 ;
        RECT 299.455 -101.595 301.335 -100.025 ;
        RECT 282.860 -112.560 283.375 -112.105 ;
        RECT 277.755 -115.200 281.140 -114.635 ;
        RECT 258.285 -118.460 264.325 -117.760 ;
        RECT 272.085 -118.380 274.280 -118.145 ;
        RECT 258.285 -118.730 270.640 -118.460 ;
        RECT 272.085 -118.565 272.320 -118.380 ;
        RECT 258.285 -119.055 264.325 -118.730 ;
        RECT 266.285 -120.930 266.935 -120.180 ;
        RECT 267.715 -120.450 267.945 -119.450 ;
        RECT 268.205 -120.590 268.435 -119.450 ;
        RECT 268.695 -120.450 268.925 -119.450 ;
        RECT 269.185 -120.590 269.415 -119.450 ;
        RECT 270.370 -120.180 270.640 -118.730 ;
        RECT 272.090 -120.060 272.320 -118.565 ;
        RECT 272.580 -120.060 272.810 -118.560 ;
        RECT 273.070 -120.060 273.300 -118.380 ;
        RECT 270.370 -120.450 272.010 -120.180 ;
        RECT 267.715 -120.820 270.900 -120.590 ;
        RECT 271.740 -120.725 272.010 -120.450 ;
        RECT 266.535 -127.950 266.805 -120.930 ;
        RECT 267.715 -122.100 267.945 -120.820 ;
        RECT 268.205 -120.830 269.415 -120.820 ;
        RECT 268.695 -122.100 268.925 -120.830 ;
        RECT 269.675 -122.100 269.905 -120.820 ;
        RECT 271.610 -121.015 272.405 -120.725 ;
        RECT 272.580 -122.745 272.810 -121.245 ;
        RECT 273.560 -122.745 273.790 -118.560 ;
        RECT 274.050 -120.060 274.280 -118.380 ;
        RECT 278.705 -120.355 279.270 -115.200 ;
        RECT 282.920 -115.725 283.315 -112.560 ;
        RECT 284.330 -113.805 284.560 -112.305 ;
        RECT 284.820 -113.805 285.050 -112.305 ;
        RECT 286.680 -113.805 286.910 -111.305 ;
        RECT 287.170 -113.805 287.400 -111.305 ;
        RECT 287.795 -113.805 288.025 -111.305 ;
        RECT 288.285 -113.805 288.515 -111.305 ;
        RECT 288.935 -113.805 289.165 -111.305 ;
        RECT 289.425 -113.805 289.655 -111.305 ;
        RECT 289.915 -113.805 290.145 -111.305 ;
        RECT 290.480 -111.335 298.590 -111.025 ;
        RECT 290.480 -111.380 290.810 -111.335 ;
        RECT 290.565 -113.805 290.795 -112.305 ;
        RECT 291.055 -113.805 291.285 -112.305 ;
        RECT 280.420 -116.120 283.315 -115.725 ;
        RECT 280.420 -117.895 280.815 -116.120 ;
        RECT 280.290 -118.380 280.870 -117.895 ;
        RECT 290.425 -118.535 292.620 -118.300 ;
        RECT 283.435 -118.615 283.920 -118.585 ;
        RECT 283.435 -118.885 288.980 -118.615 ;
        RECT 290.425 -118.720 290.660 -118.535 ;
        RECT 283.435 -118.915 283.920 -118.885 ;
        RECT 277.560 -120.920 281.100 -120.355 ;
        RECT 275.625 -121.595 275.855 -121.095 ;
        RECT 276.115 -121.740 276.345 -121.095 ;
        RECT 276.605 -121.595 276.835 -121.095 ;
        RECT 277.095 -121.740 277.325 -121.095 ;
        RECT 275.625 -121.970 278.810 -121.740 ;
        RECT 275.625 -122.750 275.855 -121.970 ;
        RECT 276.115 -121.980 277.325 -121.970 ;
        RECT 276.605 -122.750 276.835 -121.980 ;
        RECT 277.585 -122.750 277.815 -121.970 ;
        RECT 267.585 -127.245 267.815 -125.745 ;
        RECT 253.890 -130.590 255.380 -128.090 ;
        RECT 265.820 -128.220 266.805 -127.950 ;
        RECT 267.095 -129.925 267.325 -128.430 ;
        RECT 267.090 -130.110 267.325 -129.925 ;
        RECT 267.585 -129.930 267.815 -128.430 ;
        RECT 268.075 -130.110 268.305 -128.430 ;
        RECT 268.565 -129.930 268.795 -125.745 ;
        RECT 270.630 -126.520 270.860 -125.740 ;
        RECT 271.610 -126.510 271.840 -125.740 ;
        RECT 271.120 -126.520 272.330 -126.510 ;
        RECT 272.590 -126.520 272.820 -125.740 ;
        RECT 270.630 -126.750 273.815 -126.520 ;
        RECT 270.630 -127.395 270.860 -126.895 ;
        RECT 271.120 -127.395 271.350 -126.750 ;
        RECT 271.610 -127.395 271.840 -126.895 ;
        RECT 272.100 -127.395 272.330 -126.750 ;
        RECT 274.820 -128.300 275.050 -125.300 ;
        RECT 275.875 -128.300 276.105 -125.300 ;
        RECT 276.365 -128.300 276.595 -125.300 ;
        RECT 276.855 -128.300 277.085 -125.300 ;
        RECT 277.915 -128.300 278.145 -125.300 ;
        RECT 269.055 -130.110 269.285 -128.430 ;
        RECT 279.070 -128.955 279.595 -128.595 ;
        RECT 279.100 -129.370 279.425 -128.955 ;
        RECT 274.325 -129.695 279.425 -129.370 ;
        RECT 267.090 -130.345 269.285 -130.110 ;
        RECT 274.820 -131.360 275.050 -129.860 ;
        RECT 275.310 -131.360 275.540 -129.860 ;
        RECT 275.800 -131.360 276.030 -129.860 ;
        RECT 277.010 -131.360 277.240 -129.860 ;
        RECT 277.500 -131.360 277.730 -129.860 ;
        RECT 280.535 -131.900 281.100 -120.920 ;
        RECT 284.625 -121.085 285.275 -120.335 ;
        RECT 286.055 -120.605 286.285 -119.605 ;
        RECT 286.545 -120.745 286.775 -119.605 ;
        RECT 287.035 -120.605 287.265 -119.605 ;
        RECT 287.525 -120.745 287.755 -119.605 ;
        RECT 288.710 -120.335 288.980 -118.885 ;
        RECT 290.430 -120.215 290.660 -118.720 ;
        RECT 290.920 -120.215 291.150 -118.715 ;
        RECT 291.410 -120.215 291.640 -118.535 ;
        RECT 288.710 -120.605 290.350 -120.335 ;
        RECT 286.055 -120.975 289.240 -120.745 ;
        RECT 290.080 -120.880 290.350 -120.605 ;
        RECT 284.875 -128.105 285.145 -121.085 ;
        RECT 286.055 -122.255 286.285 -120.975 ;
        RECT 286.545 -120.985 287.755 -120.975 ;
        RECT 287.035 -122.255 287.265 -120.985 ;
        RECT 288.015 -122.255 288.245 -120.975 ;
        RECT 289.950 -121.170 290.745 -120.880 ;
        RECT 290.920 -122.900 291.150 -121.400 ;
        RECT 291.900 -122.900 292.130 -118.715 ;
        RECT 292.390 -120.215 292.620 -118.535 ;
        RECT 295.900 -121.075 299.440 -120.510 ;
        RECT 293.965 -121.750 294.195 -121.250 ;
        RECT 294.455 -121.895 294.685 -121.250 ;
        RECT 294.945 -121.750 295.175 -121.250 ;
        RECT 295.435 -121.895 295.665 -121.250 ;
        RECT 293.965 -122.125 297.150 -121.895 ;
        RECT 293.965 -122.905 294.195 -122.125 ;
        RECT 294.455 -122.135 295.665 -122.125 ;
        RECT 294.945 -122.905 295.175 -122.135 ;
        RECT 295.925 -122.905 296.155 -122.125 ;
        RECT 285.925 -127.400 286.155 -125.900 ;
        RECT 284.160 -128.375 285.145 -128.105 ;
        RECT 285.435 -130.080 285.665 -128.585 ;
        RECT 285.430 -130.265 285.665 -130.080 ;
        RECT 285.925 -130.085 286.155 -128.585 ;
        RECT 286.415 -130.265 286.645 -128.585 ;
        RECT 286.905 -130.085 287.135 -125.900 ;
        RECT 288.970 -126.675 289.200 -125.895 ;
        RECT 289.950 -126.665 290.180 -125.895 ;
        RECT 289.460 -126.675 290.670 -126.665 ;
        RECT 290.930 -126.675 291.160 -125.895 ;
        RECT 288.970 -126.905 292.155 -126.675 ;
        RECT 288.970 -127.550 289.200 -127.050 ;
        RECT 289.460 -127.550 289.690 -126.905 ;
        RECT 289.950 -127.550 290.180 -127.050 ;
        RECT 290.440 -127.550 290.670 -126.905 ;
        RECT 293.160 -128.455 293.390 -125.455 ;
        RECT 294.215 -128.455 294.445 -125.455 ;
        RECT 294.705 -128.455 294.935 -125.455 ;
        RECT 295.195 -128.455 295.425 -125.455 ;
        RECT 296.255 -128.455 296.485 -125.455 ;
        RECT 287.395 -130.265 287.625 -128.585 ;
        RECT 297.410 -129.110 297.935 -128.750 ;
        RECT 297.440 -129.525 297.765 -129.110 ;
        RECT 292.665 -129.850 297.765 -129.525 ;
        RECT 285.430 -130.500 287.625 -130.265 ;
        RECT 293.160 -131.515 293.390 -130.015 ;
        RECT 293.650 -131.515 293.880 -130.015 ;
        RECT 294.140 -131.515 294.370 -130.015 ;
        RECT 295.350 -131.515 295.580 -130.015 ;
        RECT 295.840 -131.515 296.070 -130.015 ;
        RECT 231.725 -132.635 253.450 -132.225 ;
        RECT 277.715 -132.055 281.100 -131.900 ;
        RECT 298.875 -132.055 299.440 -121.075 ;
        RECT 299.970 -128.780 301.075 -101.595 ;
        RECT 302.230 -117.460 303.420 -99.840 ;
        RECT 307.460 -100.865 308.710 -100.365 ;
        RECT 315.895 -100.785 318.090 -100.550 ;
        RECT 307.460 -101.135 314.450 -100.865 ;
        RECT 315.895 -100.970 316.130 -100.785 ;
        RECT 307.460 -101.510 308.710 -101.135 ;
        RECT 310.095 -103.335 310.745 -102.585 ;
        RECT 311.525 -102.855 311.755 -101.855 ;
        RECT 312.015 -102.995 312.245 -101.855 ;
        RECT 312.505 -102.855 312.735 -101.855 ;
        RECT 312.995 -102.995 313.225 -101.855 ;
        RECT 314.180 -102.585 314.450 -101.135 ;
        RECT 315.900 -102.465 316.130 -100.970 ;
        RECT 316.390 -102.465 316.620 -100.965 ;
        RECT 316.880 -102.465 317.110 -100.785 ;
        RECT 314.180 -102.855 315.820 -102.585 ;
        RECT 311.525 -103.225 314.710 -102.995 ;
        RECT 315.550 -103.130 315.820 -102.855 ;
        RECT 310.345 -110.355 310.615 -103.335 ;
        RECT 311.525 -104.505 311.755 -103.225 ;
        RECT 312.015 -103.235 313.225 -103.225 ;
        RECT 312.505 -104.505 312.735 -103.235 ;
        RECT 313.485 -104.505 313.715 -103.225 ;
        RECT 315.420 -103.420 316.215 -103.130 ;
        RECT 316.390 -105.150 316.620 -103.650 ;
        RECT 317.370 -105.150 317.600 -100.965 ;
        RECT 317.860 -102.465 318.090 -100.785 ;
        RECT 321.370 -103.325 324.910 -102.760 ;
        RECT 319.435 -104.000 319.665 -103.500 ;
        RECT 319.925 -104.145 320.155 -103.500 ;
        RECT 320.415 -104.000 320.645 -103.500 ;
        RECT 320.905 -104.145 321.135 -103.500 ;
        RECT 319.435 -104.375 322.620 -104.145 ;
        RECT 319.435 -105.155 319.665 -104.375 ;
        RECT 319.925 -104.385 321.135 -104.375 ;
        RECT 320.415 -105.155 320.645 -104.385 ;
        RECT 321.395 -105.155 321.625 -104.375 ;
        RECT 311.395 -109.650 311.625 -108.150 ;
        RECT 309.630 -110.625 310.615 -110.355 ;
        RECT 310.905 -112.330 311.135 -110.835 ;
        RECT 310.900 -112.515 311.135 -112.330 ;
        RECT 311.395 -112.335 311.625 -110.835 ;
        RECT 311.885 -112.515 312.115 -110.835 ;
        RECT 312.375 -112.335 312.605 -108.150 ;
        RECT 314.440 -108.925 314.670 -108.145 ;
        RECT 315.420 -108.915 315.650 -108.145 ;
        RECT 314.930 -108.925 316.140 -108.915 ;
        RECT 316.400 -108.925 316.630 -108.145 ;
        RECT 314.440 -109.155 317.625 -108.925 ;
        RECT 314.440 -109.800 314.670 -109.300 ;
        RECT 314.930 -109.800 315.160 -109.155 ;
        RECT 315.420 -109.800 315.650 -109.300 ;
        RECT 315.910 -109.800 316.140 -109.155 ;
        RECT 318.630 -110.705 318.860 -107.705 ;
        RECT 319.685 -110.705 319.915 -107.705 ;
        RECT 320.175 -110.705 320.405 -107.705 ;
        RECT 320.665 -110.705 320.895 -107.705 ;
        RECT 321.725 -110.705 321.955 -107.705 ;
        RECT 312.865 -112.515 313.095 -110.835 ;
        RECT 322.880 -111.360 323.405 -111.000 ;
        RECT 322.910 -111.775 323.235 -111.360 ;
        RECT 318.135 -112.100 323.235 -111.775 ;
        RECT 310.900 -112.750 313.095 -112.515 ;
        RECT 318.630 -113.765 318.860 -112.265 ;
        RECT 319.120 -113.765 319.350 -112.265 ;
        RECT 319.610 -113.765 319.840 -112.265 ;
        RECT 320.820 -113.765 321.050 -112.265 ;
        RECT 321.310 -113.765 321.540 -112.265 ;
        RECT 322.475 -114.305 323.040 -114.300 ;
        RECT 324.345 -114.305 324.910 -103.325 ;
        RECT 328.590 -109.495 328.820 -106.995 ;
        RECT 329.935 -109.495 330.165 -106.995 ;
        RECT 330.425 -109.495 330.655 -106.995 ;
        RECT 330.915 -109.495 331.145 -106.995 ;
        RECT 331.565 -109.495 331.795 -106.995 ;
        RECT 333.195 -109.495 333.425 -106.995 ;
        RECT 334.335 -108.495 334.565 -106.995 ;
        RECT 327.435 -110.295 328.125 -110.275 ;
        RECT 331.465 -110.295 332.155 -110.275 ;
        RECT 333.390 -110.295 333.660 -109.930 ;
        RECT 327.435 -110.515 333.660 -110.295 ;
        RECT 327.435 -110.545 328.125 -110.515 ;
        RECT 331.465 -110.545 332.155 -110.515 ;
        RECT 333.390 -110.620 333.660 -110.515 ;
        RECT 334.250 -110.695 334.580 -110.635 ;
        RECT 340.960 -110.695 342.150 -99.840 ;
        RECT 343.735 -100.050 344.620 -84.140 ;
        RECT 346.160 -99.880 388.100 -98.380 ;
        RECT 343.335 -101.505 345.025 -100.050 ;
        RECT 326.630 -112.230 327.145 -111.775 ;
        RECT 321.525 -114.870 324.910 -114.305 ;
        RECT 302.230 -118.130 307.910 -117.460 ;
        RECT 315.855 -118.050 318.050 -117.815 ;
        RECT 302.230 -118.400 314.410 -118.130 ;
        RECT 315.855 -118.235 316.090 -118.050 ;
        RECT 302.230 -118.650 307.910 -118.400 ;
        RECT 310.055 -120.600 310.705 -119.850 ;
        RECT 311.485 -120.120 311.715 -119.120 ;
        RECT 311.975 -120.260 312.205 -119.120 ;
        RECT 312.465 -120.120 312.695 -119.120 ;
        RECT 312.955 -120.260 313.185 -119.120 ;
        RECT 314.140 -119.850 314.410 -118.400 ;
        RECT 315.860 -119.730 316.090 -118.235 ;
        RECT 316.350 -119.730 316.580 -118.230 ;
        RECT 316.840 -119.730 317.070 -118.050 ;
        RECT 314.140 -120.120 315.780 -119.850 ;
        RECT 311.485 -120.490 314.670 -120.260 ;
        RECT 315.510 -120.395 315.780 -120.120 ;
        RECT 310.305 -127.620 310.575 -120.600 ;
        RECT 311.485 -121.770 311.715 -120.490 ;
        RECT 311.975 -120.500 313.185 -120.490 ;
        RECT 312.465 -121.770 312.695 -120.500 ;
        RECT 313.445 -121.770 313.675 -120.490 ;
        RECT 315.380 -120.685 316.175 -120.395 ;
        RECT 316.350 -122.415 316.580 -120.915 ;
        RECT 317.330 -122.415 317.560 -118.230 ;
        RECT 317.820 -119.730 318.050 -118.050 ;
        RECT 322.475 -120.025 323.040 -114.870 ;
        RECT 326.690 -115.395 327.085 -112.230 ;
        RECT 328.100 -113.475 328.330 -111.975 ;
        RECT 328.590 -113.475 328.820 -111.975 ;
        RECT 330.450 -113.475 330.680 -110.975 ;
        RECT 330.940 -113.475 331.170 -110.975 ;
        RECT 331.565 -113.475 331.795 -110.975 ;
        RECT 332.055 -113.475 332.285 -110.975 ;
        RECT 332.705 -113.475 332.935 -110.975 ;
        RECT 333.195 -113.475 333.425 -110.975 ;
        RECT 333.685 -113.475 333.915 -110.975 ;
        RECT 334.250 -111.005 342.360 -110.695 ;
        RECT 334.250 -111.050 334.580 -111.005 ;
        RECT 334.335 -113.475 334.565 -111.975 ;
        RECT 334.825 -113.475 335.055 -111.975 ;
        RECT 324.190 -115.790 327.085 -115.395 ;
        RECT 324.190 -117.565 324.585 -115.790 ;
        RECT 324.060 -118.050 324.640 -117.565 ;
        RECT 334.195 -118.205 336.390 -117.970 ;
        RECT 327.205 -118.285 327.690 -118.255 ;
        RECT 327.205 -118.555 332.750 -118.285 ;
        RECT 334.195 -118.390 334.430 -118.205 ;
        RECT 327.205 -118.585 327.690 -118.555 ;
        RECT 321.330 -120.590 324.870 -120.025 ;
        RECT 319.395 -121.265 319.625 -120.765 ;
        RECT 319.885 -121.410 320.115 -120.765 ;
        RECT 320.375 -121.265 320.605 -120.765 ;
        RECT 320.865 -121.410 321.095 -120.765 ;
        RECT 319.395 -121.640 322.580 -121.410 ;
        RECT 319.395 -122.420 319.625 -121.640 ;
        RECT 319.885 -121.650 321.095 -121.640 ;
        RECT 320.375 -122.420 320.605 -121.650 ;
        RECT 321.355 -122.420 321.585 -121.640 ;
        RECT 311.355 -126.915 311.585 -125.415 ;
        RECT 309.590 -127.890 310.575 -127.620 ;
        RECT 299.700 -130.275 301.160 -128.780 ;
        RECT 310.865 -129.595 311.095 -128.100 ;
        RECT 310.860 -129.780 311.095 -129.595 ;
        RECT 311.355 -129.600 311.585 -128.100 ;
        RECT 311.845 -129.780 312.075 -128.100 ;
        RECT 312.335 -129.600 312.565 -125.415 ;
        RECT 314.400 -126.190 314.630 -125.410 ;
        RECT 315.380 -126.180 315.610 -125.410 ;
        RECT 314.890 -126.190 316.100 -126.180 ;
        RECT 316.360 -126.190 316.590 -125.410 ;
        RECT 314.400 -126.420 317.585 -126.190 ;
        RECT 314.400 -127.065 314.630 -126.565 ;
        RECT 314.890 -127.065 315.120 -126.420 ;
        RECT 315.380 -127.065 315.610 -126.565 ;
        RECT 315.870 -127.065 316.100 -126.420 ;
        RECT 318.590 -127.970 318.820 -124.970 ;
        RECT 319.645 -127.970 319.875 -124.970 ;
        RECT 320.135 -127.970 320.365 -124.970 ;
        RECT 320.625 -127.970 320.855 -124.970 ;
        RECT 321.685 -127.970 321.915 -124.970 ;
        RECT 312.825 -129.780 313.055 -128.100 ;
        RECT 322.840 -128.625 323.365 -128.265 ;
        RECT 322.870 -129.040 323.195 -128.625 ;
        RECT 318.095 -129.365 323.195 -129.040 ;
        RECT 310.860 -130.015 313.055 -129.780 ;
        RECT 318.590 -131.030 318.820 -129.530 ;
        RECT 319.080 -131.030 319.310 -129.530 ;
        RECT 319.570 -131.030 319.800 -129.530 ;
        RECT 320.780 -131.030 321.010 -129.530 ;
        RECT 321.270 -131.030 321.500 -129.530 ;
        RECT 324.305 -131.570 324.870 -120.590 ;
        RECT 328.395 -120.755 329.045 -120.005 ;
        RECT 329.825 -120.275 330.055 -119.275 ;
        RECT 330.315 -120.415 330.545 -119.275 ;
        RECT 330.805 -120.275 331.035 -119.275 ;
        RECT 331.295 -120.415 331.525 -119.275 ;
        RECT 332.480 -120.005 332.750 -118.555 ;
        RECT 334.200 -119.885 334.430 -118.390 ;
        RECT 334.690 -119.885 334.920 -118.385 ;
        RECT 335.180 -119.885 335.410 -118.205 ;
        RECT 332.480 -120.275 334.120 -120.005 ;
        RECT 329.825 -120.645 333.010 -120.415 ;
        RECT 333.850 -120.550 334.120 -120.275 ;
        RECT 328.645 -127.775 328.915 -120.755 ;
        RECT 329.825 -121.925 330.055 -120.645 ;
        RECT 330.315 -120.655 331.525 -120.645 ;
        RECT 330.805 -121.925 331.035 -120.655 ;
        RECT 331.785 -121.925 332.015 -120.645 ;
        RECT 333.720 -120.840 334.515 -120.550 ;
        RECT 334.690 -122.570 334.920 -121.070 ;
        RECT 335.670 -122.570 335.900 -118.385 ;
        RECT 336.160 -119.885 336.390 -118.205 ;
        RECT 339.670 -120.745 343.210 -120.180 ;
        RECT 337.735 -121.420 337.965 -120.920 ;
        RECT 338.225 -121.565 338.455 -120.920 ;
        RECT 338.715 -121.420 338.945 -120.920 ;
        RECT 339.205 -121.565 339.435 -120.920 ;
        RECT 337.735 -121.795 340.920 -121.565 ;
        RECT 337.735 -122.575 337.965 -121.795 ;
        RECT 338.225 -121.805 339.435 -121.795 ;
        RECT 338.715 -122.575 338.945 -121.805 ;
        RECT 339.695 -122.575 339.925 -121.795 ;
        RECT 329.695 -127.070 329.925 -125.570 ;
        RECT 327.930 -128.045 328.915 -127.775 ;
        RECT 329.205 -129.750 329.435 -128.255 ;
        RECT 329.200 -129.935 329.435 -129.750 ;
        RECT 329.695 -129.755 329.925 -128.255 ;
        RECT 330.185 -129.935 330.415 -128.255 ;
        RECT 330.675 -129.755 330.905 -125.570 ;
        RECT 332.740 -126.345 332.970 -125.565 ;
        RECT 333.720 -126.335 333.950 -125.565 ;
        RECT 333.230 -126.345 334.440 -126.335 ;
        RECT 334.700 -126.345 334.930 -125.565 ;
        RECT 332.740 -126.575 335.925 -126.345 ;
        RECT 332.740 -127.220 332.970 -126.720 ;
        RECT 333.230 -127.220 333.460 -126.575 ;
        RECT 333.720 -127.220 333.950 -126.720 ;
        RECT 334.210 -127.220 334.440 -126.575 ;
        RECT 336.930 -128.125 337.160 -125.125 ;
        RECT 337.985 -128.125 338.215 -125.125 ;
        RECT 338.475 -128.125 338.705 -125.125 ;
        RECT 338.965 -128.125 339.195 -125.125 ;
        RECT 340.025 -128.125 340.255 -125.125 ;
        RECT 331.165 -129.935 331.395 -128.255 ;
        RECT 341.180 -128.780 341.705 -128.420 ;
        RECT 341.210 -129.195 341.535 -128.780 ;
        RECT 336.435 -129.520 341.535 -129.195 ;
        RECT 329.200 -130.170 331.395 -129.935 ;
        RECT 336.930 -131.185 337.160 -129.685 ;
        RECT 337.420 -131.185 337.650 -129.685 ;
        RECT 337.910 -131.185 338.140 -129.685 ;
        RECT 339.120 -131.185 339.350 -129.685 ;
        RECT 339.610 -131.185 339.840 -129.685 ;
        RECT 277.715 -132.465 299.440 -132.055 ;
        RECT 321.485 -131.725 324.870 -131.570 ;
        RECT 342.645 -131.725 343.210 -120.745 ;
        RECT 343.735 -128.490 344.620 -101.505 ;
        RECT 346.160 -117.130 347.660 -99.880 ;
        RECT 353.275 -100.780 354.615 -100.325 ;
        RECT 361.660 -100.700 363.855 -100.465 ;
        RECT 353.275 -101.050 360.215 -100.780 ;
        RECT 361.660 -100.885 361.895 -100.700 ;
        RECT 353.275 -101.525 354.615 -101.050 ;
        RECT 355.860 -103.250 356.510 -102.500 ;
        RECT 357.290 -102.770 357.520 -101.770 ;
        RECT 357.780 -102.910 358.010 -101.770 ;
        RECT 358.270 -102.770 358.500 -101.770 ;
        RECT 358.760 -102.910 358.990 -101.770 ;
        RECT 359.945 -102.500 360.215 -101.050 ;
        RECT 361.665 -102.380 361.895 -100.885 ;
        RECT 362.155 -102.380 362.385 -100.880 ;
        RECT 362.645 -102.380 362.875 -100.700 ;
        RECT 359.945 -102.770 361.585 -102.500 ;
        RECT 357.290 -103.140 360.475 -102.910 ;
        RECT 361.315 -103.045 361.585 -102.770 ;
        RECT 356.110 -110.270 356.380 -103.250 ;
        RECT 357.290 -104.420 357.520 -103.140 ;
        RECT 357.780 -103.150 358.990 -103.140 ;
        RECT 358.270 -104.420 358.500 -103.150 ;
        RECT 359.250 -104.420 359.480 -103.140 ;
        RECT 361.185 -103.335 361.980 -103.045 ;
        RECT 362.155 -105.065 362.385 -103.565 ;
        RECT 363.135 -105.065 363.365 -100.880 ;
        RECT 363.625 -102.380 363.855 -100.700 ;
        RECT 367.135 -103.240 370.675 -102.675 ;
        RECT 365.200 -103.915 365.430 -103.415 ;
        RECT 365.690 -104.060 365.920 -103.415 ;
        RECT 366.180 -103.915 366.410 -103.415 ;
        RECT 366.670 -104.060 366.900 -103.415 ;
        RECT 365.200 -104.290 368.385 -104.060 ;
        RECT 365.200 -105.070 365.430 -104.290 ;
        RECT 365.690 -104.300 366.900 -104.290 ;
        RECT 366.180 -105.070 366.410 -104.300 ;
        RECT 367.160 -105.070 367.390 -104.290 ;
        RECT 357.160 -109.565 357.390 -108.065 ;
        RECT 355.395 -110.540 356.380 -110.270 ;
        RECT 356.670 -112.245 356.900 -110.750 ;
        RECT 356.665 -112.430 356.900 -112.245 ;
        RECT 357.160 -112.250 357.390 -110.750 ;
        RECT 357.650 -112.430 357.880 -110.750 ;
        RECT 358.140 -112.250 358.370 -108.065 ;
        RECT 360.205 -108.840 360.435 -108.060 ;
        RECT 361.185 -108.830 361.415 -108.060 ;
        RECT 360.695 -108.840 361.905 -108.830 ;
        RECT 362.165 -108.840 362.395 -108.060 ;
        RECT 360.205 -109.070 363.390 -108.840 ;
        RECT 360.205 -109.715 360.435 -109.215 ;
        RECT 360.695 -109.715 360.925 -109.070 ;
        RECT 361.185 -109.715 361.415 -109.215 ;
        RECT 361.675 -109.715 361.905 -109.070 ;
        RECT 364.395 -110.620 364.625 -107.620 ;
        RECT 365.450 -110.620 365.680 -107.620 ;
        RECT 365.940 -110.620 366.170 -107.620 ;
        RECT 366.430 -110.620 366.660 -107.620 ;
        RECT 367.490 -110.620 367.720 -107.620 ;
        RECT 358.630 -112.430 358.860 -110.750 ;
        RECT 368.645 -111.275 369.170 -110.915 ;
        RECT 368.675 -111.690 369.000 -111.275 ;
        RECT 363.900 -112.015 369.000 -111.690 ;
        RECT 356.665 -112.665 358.860 -112.430 ;
        RECT 364.395 -113.680 364.625 -112.180 ;
        RECT 364.885 -113.680 365.115 -112.180 ;
        RECT 365.375 -113.680 365.605 -112.180 ;
        RECT 366.585 -113.680 366.815 -112.180 ;
        RECT 367.075 -113.680 367.305 -112.180 ;
        RECT 368.240 -114.220 368.805 -114.215 ;
        RECT 370.110 -114.220 370.675 -103.240 ;
        RECT 374.355 -109.410 374.585 -106.910 ;
        RECT 375.700 -109.410 375.930 -106.910 ;
        RECT 376.190 -109.410 376.420 -106.910 ;
        RECT 376.680 -109.410 376.910 -106.910 ;
        RECT 377.330 -109.410 377.560 -106.910 ;
        RECT 378.960 -109.410 379.190 -106.910 ;
        RECT 380.100 -108.410 380.330 -106.910 ;
        RECT 373.200 -110.210 373.890 -110.190 ;
        RECT 377.230 -110.210 377.920 -110.190 ;
        RECT 379.155 -110.210 379.425 -109.845 ;
        RECT 373.200 -110.430 379.425 -110.210 ;
        RECT 373.200 -110.460 373.890 -110.430 ;
        RECT 377.230 -110.460 377.920 -110.430 ;
        RECT 379.155 -110.535 379.425 -110.430 ;
        RECT 380.015 -110.610 380.345 -110.550 ;
        RECT 386.565 -110.610 388.100 -99.880 ;
        RECT 372.395 -112.145 372.910 -111.690 ;
        RECT 367.290 -114.785 370.675 -114.220 ;
        RECT 346.160 -118.045 353.610 -117.130 ;
        RECT 361.620 -117.965 363.815 -117.730 ;
        RECT 346.160 -118.315 360.175 -118.045 ;
        RECT 361.620 -118.150 361.855 -117.965 ;
        RECT 346.160 -118.630 353.610 -118.315 ;
        RECT 355.820 -120.515 356.470 -119.765 ;
        RECT 357.250 -120.035 357.480 -119.035 ;
        RECT 357.740 -120.175 357.970 -119.035 ;
        RECT 358.230 -120.035 358.460 -119.035 ;
        RECT 358.720 -120.175 358.950 -119.035 ;
        RECT 359.905 -119.765 360.175 -118.315 ;
        RECT 361.625 -119.645 361.855 -118.150 ;
        RECT 362.115 -119.645 362.345 -118.145 ;
        RECT 362.605 -119.645 362.835 -117.965 ;
        RECT 359.905 -120.035 361.545 -119.765 ;
        RECT 357.250 -120.405 360.435 -120.175 ;
        RECT 361.275 -120.310 361.545 -120.035 ;
        RECT 356.070 -127.535 356.340 -120.515 ;
        RECT 357.250 -121.685 357.480 -120.405 ;
        RECT 357.740 -120.415 358.950 -120.405 ;
        RECT 358.230 -121.685 358.460 -120.415 ;
        RECT 359.210 -121.685 359.440 -120.405 ;
        RECT 361.145 -120.600 361.940 -120.310 ;
        RECT 362.115 -122.330 362.345 -120.830 ;
        RECT 363.095 -122.330 363.325 -118.145 ;
        RECT 363.585 -119.645 363.815 -117.965 ;
        RECT 368.240 -119.940 368.805 -114.785 ;
        RECT 372.455 -115.310 372.850 -112.145 ;
        RECT 373.865 -113.390 374.095 -111.890 ;
        RECT 374.355 -113.390 374.585 -111.890 ;
        RECT 376.215 -113.390 376.445 -110.890 ;
        RECT 376.705 -113.390 376.935 -110.890 ;
        RECT 377.330 -113.390 377.560 -110.890 ;
        RECT 377.820 -113.390 378.050 -110.890 ;
        RECT 378.470 -113.390 378.700 -110.890 ;
        RECT 378.960 -113.390 379.190 -110.890 ;
        RECT 379.450 -113.390 379.680 -110.890 ;
        RECT 380.015 -110.920 388.125 -110.610 ;
        RECT 380.015 -110.965 380.345 -110.920 ;
        RECT 380.100 -113.390 380.330 -111.890 ;
        RECT 380.590 -113.390 380.820 -111.890 ;
        RECT 369.955 -115.705 372.850 -115.310 ;
        RECT 369.955 -117.480 370.350 -115.705 ;
        RECT 369.825 -117.965 370.405 -117.480 ;
        RECT 379.960 -118.120 382.155 -117.885 ;
        RECT 372.970 -118.200 373.455 -118.170 ;
        RECT 372.970 -118.470 378.515 -118.200 ;
        RECT 379.960 -118.305 380.195 -118.120 ;
        RECT 372.970 -118.500 373.455 -118.470 ;
        RECT 367.095 -120.505 370.635 -119.940 ;
        RECT 365.160 -121.180 365.390 -120.680 ;
        RECT 365.650 -121.325 365.880 -120.680 ;
        RECT 366.140 -121.180 366.370 -120.680 ;
        RECT 366.630 -121.325 366.860 -120.680 ;
        RECT 365.160 -121.555 368.345 -121.325 ;
        RECT 365.160 -122.335 365.390 -121.555 ;
        RECT 365.650 -121.565 366.860 -121.555 ;
        RECT 366.140 -122.335 366.370 -121.565 ;
        RECT 367.120 -122.335 367.350 -121.555 ;
        RECT 357.120 -126.830 357.350 -125.330 ;
        RECT 355.355 -127.805 356.340 -127.535 ;
        RECT 343.525 -130.010 344.830 -128.490 ;
        RECT 356.630 -129.510 356.860 -128.015 ;
        RECT 356.625 -129.695 356.860 -129.510 ;
        RECT 357.120 -129.515 357.350 -128.015 ;
        RECT 357.610 -129.695 357.840 -128.015 ;
        RECT 358.100 -129.515 358.330 -125.330 ;
        RECT 360.165 -126.105 360.395 -125.325 ;
        RECT 361.145 -126.095 361.375 -125.325 ;
        RECT 360.655 -126.105 361.865 -126.095 ;
        RECT 362.125 -126.105 362.355 -125.325 ;
        RECT 360.165 -126.335 363.350 -126.105 ;
        RECT 360.165 -126.980 360.395 -126.480 ;
        RECT 360.655 -126.980 360.885 -126.335 ;
        RECT 361.145 -126.980 361.375 -126.480 ;
        RECT 361.635 -126.980 361.865 -126.335 ;
        RECT 364.355 -127.885 364.585 -124.885 ;
        RECT 365.410 -127.885 365.640 -124.885 ;
        RECT 365.900 -127.885 366.130 -124.885 ;
        RECT 366.390 -127.885 366.620 -124.885 ;
        RECT 367.450 -127.885 367.680 -124.885 ;
        RECT 358.590 -129.695 358.820 -128.015 ;
        RECT 368.605 -128.540 369.130 -128.180 ;
        RECT 368.635 -128.955 368.960 -128.540 ;
        RECT 363.860 -129.280 368.960 -128.955 ;
        RECT 356.625 -129.930 358.820 -129.695 ;
        RECT 364.355 -130.945 364.585 -129.445 ;
        RECT 364.845 -130.945 365.075 -129.445 ;
        RECT 365.335 -130.945 365.565 -129.445 ;
        RECT 366.545 -130.945 366.775 -129.445 ;
        RECT 367.035 -130.945 367.265 -129.445 ;
        RECT 370.070 -131.485 370.635 -120.505 ;
        RECT 374.160 -120.670 374.810 -119.920 ;
        RECT 375.590 -120.190 375.820 -119.190 ;
        RECT 376.080 -120.330 376.310 -119.190 ;
        RECT 376.570 -120.190 376.800 -119.190 ;
        RECT 377.060 -120.330 377.290 -119.190 ;
        RECT 378.245 -119.920 378.515 -118.470 ;
        RECT 379.965 -119.800 380.195 -118.305 ;
        RECT 380.455 -119.800 380.685 -118.300 ;
        RECT 380.945 -119.800 381.175 -118.120 ;
        RECT 378.245 -120.190 379.885 -119.920 ;
        RECT 375.590 -120.560 378.775 -120.330 ;
        RECT 379.615 -120.465 379.885 -120.190 ;
        RECT 374.410 -127.690 374.680 -120.670 ;
        RECT 375.590 -121.840 375.820 -120.560 ;
        RECT 376.080 -120.570 377.290 -120.560 ;
        RECT 376.570 -121.840 376.800 -120.570 ;
        RECT 377.550 -121.840 377.780 -120.560 ;
        RECT 379.485 -120.755 380.280 -120.465 ;
        RECT 380.455 -122.485 380.685 -120.985 ;
        RECT 381.435 -122.485 381.665 -118.300 ;
        RECT 381.925 -119.800 382.155 -118.120 ;
        RECT 385.435 -120.660 388.975 -120.095 ;
        RECT 383.500 -121.335 383.730 -120.835 ;
        RECT 383.990 -121.480 384.220 -120.835 ;
        RECT 384.480 -121.335 384.710 -120.835 ;
        RECT 384.970 -121.480 385.200 -120.835 ;
        RECT 383.500 -121.710 386.685 -121.480 ;
        RECT 383.500 -122.490 383.730 -121.710 ;
        RECT 383.990 -121.720 385.200 -121.710 ;
        RECT 384.480 -122.490 384.710 -121.720 ;
        RECT 385.460 -122.490 385.690 -121.710 ;
        RECT 375.460 -126.985 375.690 -125.485 ;
        RECT 373.695 -127.960 374.680 -127.690 ;
        RECT 374.970 -129.665 375.200 -128.170 ;
        RECT 374.965 -129.850 375.200 -129.665 ;
        RECT 375.460 -129.670 375.690 -128.170 ;
        RECT 375.950 -129.850 376.180 -128.170 ;
        RECT 376.440 -129.670 376.670 -125.485 ;
        RECT 378.505 -126.260 378.735 -125.480 ;
        RECT 379.485 -126.250 379.715 -125.480 ;
        RECT 378.995 -126.260 380.205 -126.250 ;
        RECT 380.465 -126.260 380.695 -125.480 ;
        RECT 378.505 -126.490 381.690 -126.260 ;
        RECT 378.505 -127.135 378.735 -126.635 ;
        RECT 378.995 -127.135 379.225 -126.490 ;
        RECT 379.485 -127.135 379.715 -126.635 ;
        RECT 379.975 -127.135 380.205 -126.490 ;
        RECT 382.695 -128.040 382.925 -125.040 ;
        RECT 383.750 -128.040 383.980 -125.040 ;
        RECT 384.240 -128.040 384.470 -125.040 ;
        RECT 384.730 -128.040 384.960 -125.040 ;
        RECT 385.790 -128.040 386.020 -125.040 ;
        RECT 376.930 -129.850 377.160 -128.170 ;
        RECT 386.945 -128.695 387.470 -128.335 ;
        RECT 386.975 -129.110 387.300 -128.695 ;
        RECT 382.200 -129.435 387.300 -129.110 ;
        RECT 374.965 -130.085 377.160 -129.850 ;
        RECT 382.695 -131.100 382.925 -129.600 ;
        RECT 383.185 -131.100 383.415 -129.600 ;
        RECT 383.675 -131.100 383.905 -129.600 ;
        RECT 384.885 -131.100 385.115 -129.600 ;
        RECT 385.375 -131.100 385.605 -129.600 ;
        RECT 321.485 -132.135 343.210 -131.725 ;
        RECT 367.250 -131.640 370.635 -131.485 ;
        RECT 388.410 -131.640 388.975 -120.660 ;
        RECT 389.405 -130.110 390.960 -81.890 ;
        RECT 392.285 -99.470 434.880 -98.375 ;
        RECT 392.285 -117.660 393.380 -99.470 ;
        RECT 399.550 -100.590 401.025 -100.015 ;
        RECT 408.480 -100.510 410.675 -100.275 ;
        RECT 399.550 -100.860 407.035 -100.590 ;
        RECT 408.480 -100.695 408.715 -100.510 ;
        RECT 399.550 -101.380 401.025 -100.860 ;
        RECT 402.680 -103.060 403.330 -102.310 ;
        RECT 404.110 -102.580 404.340 -101.580 ;
        RECT 404.600 -102.720 404.830 -101.580 ;
        RECT 405.090 -102.580 405.320 -101.580 ;
        RECT 405.580 -102.720 405.810 -101.580 ;
        RECT 406.765 -102.310 407.035 -100.860 ;
        RECT 408.485 -102.190 408.715 -100.695 ;
        RECT 408.975 -102.190 409.205 -100.690 ;
        RECT 409.465 -102.190 409.695 -100.510 ;
        RECT 406.765 -102.580 408.405 -102.310 ;
        RECT 404.110 -102.950 407.295 -102.720 ;
        RECT 408.135 -102.855 408.405 -102.580 ;
        RECT 402.930 -110.080 403.200 -103.060 ;
        RECT 404.110 -104.230 404.340 -102.950 ;
        RECT 404.600 -102.960 405.810 -102.950 ;
        RECT 405.090 -104.230 405.320 -102.960 ;
        RECT 406.070 -104.230 406.300 -102.950 ;
        RECT 408.005 -103.145 408.800 -102.855 ;
        RECT 408.975 -104.875 409.205 -103.375 ;
        RECT 409.955 -104.875 410.185 -100.690 ;
        RECT 410.445 -102.190 410.675 -100.510 ;
        RECT 413.955 -103.050 417.495 -102.485 ;
        RECT 412.020 -103.725 412.250 -103.225 ;
        RECT 412.510 -103.870 412.740 -103.225 ;
        RECT 413.000 -103.725 413.230 -103.225 ;
        RECT 413.490 -103.870 413.720 -103.225 ;
        RECT 412.020 -104.100 415.205 -103.870 ;
        RECT 412.020 -104.880 412.250 -104.100 ;
        RECT 412.510 -104.110 413.720 -104.100 ;
        RECT 413.000 -104.880 413.230 -104.110 ;
        RECT 413.980 -104.880 414.210 -104.100 ;
        RECT 403.980 -109.375 404.210 -107.875 ;
        RECT 402.215 -110.350 403.200 -110.080 ;
        RECT 403.490 -112.055 403.720 -110.560 ;
        RECT 403.485 -112.240 403.720 -112.055 ;
        RECT 403.980 -112.060 404.210 -110.560 ;
        RECT 404.470 -112.240 404.700 -110.560 ;
        RECT 404.960 -112.060 405.190 -107.875 ;
        RECT 407.025 -108.650 407.255 -107.870 ;
        RECT 408.005 -108.640 408.235 -107.870 ;
        RECT 407.515 -108.650 408.725 -108.640 ;
        RECT 408.985 -108.650 409.215 -107.870 ;
        RECT 407.025 -108.880 410.210 -108.650 ;
        RECT 407.025 -109.525 407.255 -109.025 ;
        RECT 407.515 -109.525 407.745 -108.880 ;
        RECT 408.005 -109.525 408.235 -109.025 ;
        RECT 408.495 -109.525 408.725 -108.880 ;
        RECT 411.215 -110.430 411.445 -107.430 ;
        RECT 412.270 -110.430 412.500 -107.430 ;
        RECT 412.760 -110.430 412.990 -107.430 ;
        RECT 413.250 -110.430 413.480 -107.430 ;
        RECT 414.310 -110.430 414.540 -107.430 ;
        RECT 405.450 -112.240 405.680 -110.560 ;
        RECT 415.465 -111.085 415.990 -110.725 ;
        RECT 415.495 -111.500 415.820 -111.085 ;
        RECT 410.720 -111.825 415.820 -111.500 ;
        RECT 403.485 -112.475 405.680 -112.240 ;
        RECT 411.215 -113.490 411.445 -111.990 ;
        RECT 411.705 -113.490 411.935 -111.990 ;
        RECT 412.195 -113.490 412.425 -111.990 ;
        RECT 413.405 -113.490 413.635 -111.990 ;
        RECT 413.895 -113.490 414.125 -111.990 ;
        RECT 415.060 -114.030 415.625 -114.025 ;
        RECT 416.930 -114.030 417.495 -103.050 ;
        RECT 421.175 -109.220 421.405 -106.720 ;
        RECT 422.520 -109.220 422.750 -106.720 ;
        RECT 423.010 -109.220 423.240 -106.720 ;
        RECT 423.500 -109.220 423.730 -106.720 ;
        RECT 424.150 -109.220 424.380 -106.720 ;
        RECT 425.780 -109.220 426.010 -106.720 ;
        RECT 426.920 -108.220 427.150 -106.720 ;
        RECT 420.020 -110.020 420.710 -110.000 ;
        RECT 424.050 -110.020 424.740 -110.000 ;
        RECT 425.975 -110.020 426.245 -109.655 ;
        RECT 420.020 -110.240 426.245 -110.020 ;
        RECT 420.020 -110.270 420.710 -110.240 ;
        RECT 424.050 -110.270 424.740 -110.240 ;
        RECT 425.975 -110.345 426.245 -110.240 ;
        RECT 426.835 -110.420 427.165 -110.360 ;
        RECT 433.785 -110.420 434.880 -99.470 ;
        RECT 419.215 -111.955 419.730 -111.500 ;
        RECT 414.110 -114.595 417.495 -114.030 ;
        RECT 392.285 -117.855 401.180 -117.660 ;
        RECT 408.440 -117.775 410.635 -117.540 ;
        RECT 392.285 -118.125 406.995 -117.855 ;
        RECT 408.440 -117.960 408.675 -117.775 ;
        RECT 392.285 -118.755 401.180 -118.125 ;
        RECT 402.640 -120.325 403.290 -119.575 ;
        RECT 404.070 -119.845 404.300 -118.845 ;
        RECT 404.560 -119.985 404.790 -118.845 ;
        RECT 405.050 -119.845 405.280 -118.845 ;
        RECT 405.540 -119.985 405.770 -118.845 ;
        RECT 406.725 -119.575 406.995 -118.125 ;
        RECT 408.445 -119.455 408.675 -117.960 ;
        RECT 408.935 -119.455 409.165 -117.955 ;
        RECT 409.425 -119.455 409.655 -117.775 ;
        RECT 406.725 -119.845 408.365 -119.575 ;
        RECT 404.070 -120.215 407.255 -119.985 ;
        RECT 408.095 -120.120 408.365 -119.845 ;
        RECT 402.890 -127.345 403.160 -120.325 ;
        RECT 404.070 -121.495 404.300 -120.215 ;
        RECT 404.560 -120.225 405.770 -120.215 ;
        RECT 405.050 -121.495 405.280 -120.225 ;
        RECT 406.030 -121.495 406.260 -120.215 ;
        RECT 407.965 -120.410 408.760 -120.120 ;
        RECT 408.935 -122.140 409.165 -120.640 ;
        RECT 409.915 -122.140 410.145 -117.955 ;
        RECT 410.405 -119.455 410.635 -117.775 ;
        RECT 415.060 -119.750 415.625 -114.595 ;
        RECT 419.275 -115.120 419.670 -111.955 ;
        RECT 420.685 -113.200 420.915 -111.700 ;
        RECT 421.175 -113.200 421.405 -111.700 ;
        RECT 423.035 -113.200 423.265 -110.700 ;
        RECT 423.525 -113.200 423.755 -110.700 ;
        RECT 424.150 -113.200 424.380 -110.700 ;
        RECT 424.640 -113.200 424.870 -110.700 ;
        RECT 425.290 -113.200 425.520 -110.700 ;
        RECT 425.780 -113.200 426.010 -110.700 ;
        RECT 426.270 -113.200 426.500 -110.700 ;
        RECT 426.835 -110.730 434.945 -110.420 ;
        RECT 426.835 -110.775 427.165 -110.730 ;
        RECT 426.920 -113.200 427.150 -111.700 ;
        RECT 427.410 -113.200 427.640 -111.700 ;
        RECT 416.775 -115.515 419.670 -115.120 ;
        RECT 416.775 -117.290 417.170 -115.515 ;
        RECT 416.645 -117.775 417.225 -117.290 ;
        RECT 426.780 -117.930 428.975 -117.695 ;
        RECT 419.790 -118.010 420.275 -117.980 ;
        RECT 419.790 -118.280 425.335 -118.010 ;
        RECT 426.780 -118.115 427.015 -117.930 ;
        RECT 419.790 -118.310 420.275 -118.280 ;
        RECT 413.915 -120.315 417.455 -119.750 ;
        RECT 411.980 -120.990 412.210 -120.490 ;
        RECT 412.470 -121.135 412.700 -120.490 ;
        RECT 412.960 -120.990 413.190 -120.490 ;
        RECT 413.450 -121.135 413.680 -120.490 ;
        RECT 411.980 -121.365 415.165 -121.135 ;
        RECT 411.980 -122.145 412.210 -121.365 ;
        RECT 412.470 -121.375 413.680 -121.365 ;
        RECT 412.960 -122.145 413.190 -121.375 ;
        RECT 413.940 -122.145 414.170 -121.365 ;
        RECT 403.940 -126.640 404.170 -125.140 ;
        RECT 402.175 -127.615 403.160 -127.345 ;
        RECT 403.450 -129.320 403.680 -127.825 ;
        RECT 403.445 -129.505 403.680 -129.320 ;
        RECT 403.940 -129.325 404.170 -127.825 ;
        RECT 404.430 -129.505 404.660 -127.825 ;
        RECT 404.920 -129.325 405.150 -125.140 ;
        RECT 406.985 -125.915 407.215 -125.135 ;
        RECT 407.965 -125.905 408.195 -125.135 ;
        RECT 407.475 -125.915 408.685 -125.905 ;
        RECT 408.945 -125.915 409.175 -125.135 ;
        RECT 406.985 -126.145 410.170 -125.915 ;
        RECT 406.985 -126.790 407.215 -126.290 ;
        RECT 407.475 -126.790 407.705 -126.145 ;
        RECT 407.965 -126.790 408.195 -126.290 ;
        RECT 408.455 -126.790 408.685 -126.145 ;
        RECT 411.175 -127.695 411.405 -124.695 ;
        RECT 412.230 -127.695 412.460 -124.695 ;
        RECT 412.720 -127.695 412.950 -124.695 ;
        RECT 413.210 -127.695 413.440 -124.695 ;
        RECT 414.270 -127.695 414.500 -124.695 ;
        RECT 405.410 -129.505 405.640 -127.825 ;
        RECT 415.425 -128.350 415.950 -127.990 ;
        RECT 415.455 -128.765 415.780 -128.350 ;
        RECT 410.680 -129.090 415.780 -128.765 ;
        RECT 403.445 -129.740 405.640 -129.505 ;
        RECT 411.175 -130.755 411.405 -129.255 ;
        RECT 411.665 -130.755 411.895 -129.255 ;
        RECT 412.155 -130.755 412.385 -129.255 ;
        RECT 413.365 -130.755 413.595 -129.255 ;
        RECT 413.855 -130.755 414.085 -129.255 ;
        RECT 416.890 -131.295 417.455 -120.315 ;
        RECT 420.980 -120.480 421.630 -119.730 ;
        RECT 422.410 -120.000 422.640 -119.000 ;
        RECT 422.900 -120.140 423.130 -119.000 ;
        RECT 423.390 -120.000 423.620 -119.000 ;
        RECT 423.880 -120.140 424.110 -119.000 ;
        RECT 425.065 -119.730 425.335 -118.280 ;
        RECT 426.785 -119.610 427.015 -118.115 ;
        RECT 427.275 -119.610 427.505 -118.110 ;
        RECT 427.765 -119.610 427.995 -117.930 ;
        RECT 425.065 -120.000 426.705 -119.730 ;
        RECT 422.410 -120.370 425.595 -120.140 ;
        RECT 426.435 -120.275 426.705 -120.000 ;
        RECT 421.230 -127.500 421.500 -120.480 ;
        RECT 422.410 -121.650 422.640 -120.370 ;
        RECT 422.900 -120.380 424.110 -120.370 ;
        RECT 423.390 -121.650 423.620 -120.380 ;
        RECT 424.370 -121.650 424.600 -120.370 ;
        RECT 426.305 -120.565 427.100 -120.275 ;
        RECT 427.275 -122.295 427.505 -120.795 ;
        RECT 428.255 -122.295 428.485 -118.110 ;
        RECT 428.745 -119.610 428.975 -117.930 ;
        RECT 432.255 -120.470 435.795 -119.905 ;
        RECT 430.320 -121.145 430.550 -120.645 ;
        RECT 430.810 -121.290 431.040 -120.645 ;
        RECT 431.300 -121.145 431.530 -120.645 ;
        RECT 431.790 -121.290 432.020 -120.645 ;
        RECT 430.320 -121.520 433.505 -121.290 ;
        RECT 430.320 -122.300 430.550 -121.520 ;
        RECT 430.810 -121.530 432.020 -121.520 ;
        RECT 431.300 -122.300 431.530 -121.530 ;
        RECT 432.280 -122.300 432.510 -121.520 ;
        RECT 422.280 -126.795 422.510 -125.295 ;
        RECT 420.515 -127.770 421.500 -127.500 ;
        RECT 421.790 -129.475 422.020 -127.980 ;
        RECT 421.785 -129.660 422.020 -129.475 ;
        RECT 422.280 -129.480 422.510 -127.980 ;
        RECT 422.770 -129.660 423.000 -127.980 ;
        RECT 423.260 -129.480 423.490 -125.295 ;
        RECT 425.325 -126.070 425.555 -125.290 ;
        RECT 426.305 -126.060 426.535 -125.290 ;
        RECT 425.815 -126.070 427.025 -126.060 ;
        RECT 427.285 -126.070 427.515 -125.290 ;
        RECT 425.325 -126.300 428.510 -126.070 ;
        RECT 425.325 -126.945 425.555 -126.445 ;
        RECT 425.815 -126.945 426.045 -126.300 ;
        RECT 426.305 -126.945 426.535 -126.445 ;
        RECT 426.795 -126.945 427.025 -126.300 ;
        RECT 429.515 -127.850 429.745 -124.850 ;
        RECT 430.570 -127.850 430.800 -124.850 ;
        RECT 431.060 -127.850 431.290 -124.850 ;
        RECT 431.550 -127.850 431.780 -124.850 ;
        RECT 432.610 -127.850 432.840 -124.850 ;
        RECT 423.750 -129.660 423.980 -127.980 ;
        RECT 433.765 -128.505 434.290 -128.145 ;
        RECT 433.795 -128.920 434.120 -128.505 ;
        RECT 429.020 -129.245 434.120 -128.920 ;
        RECT 421.785 -129.895 423.980 -129.660 ;
        RECT 429.515 -130.910 429.745 -129.410 ;
        RECT 430.005 -130.910 430.235 -129.410 ;
        RECT 430.495 -130.910 430.725 -129.410 ;
        RECT 431.705 -130.910 431.935 -129.410 ;
        RECT 432.195 -130.910 432.425 -129.410 ;
        RECT 367.250 -132.050 388.975 -131.640 ;
        RECT 414.070 -131.450 417.455 -131.295 ;
        RECT 435.230 -131.450 435.795 -120.470 ;
        RECT 437.060 -128.270 438.480 -77.225 ;
        RECT 436.910 -129.985 438.705 -128.270 ;
        RECT 414.070 -131.860 435.795 -131.450 ;
        RECT 414.090 -132.015 435.795 -131.860 ;
        RECT 321.505 -132.290 343.210 -132.135 ;
        RECT 367.270 -132.205 388.975 -132.050 ;
        RECT 277.735 -132.620 299.440 -132.465 ;
        RECT 231.745 -132.790 253.450 -132.635 ;
        RECT 439.580 -134.715 440.805 -17.905 ;
        RECT 207.885 -135.660 209.470 -135.245 ;
        RECT 129.385 -136.565 173.385 -135.660 ;
        RECT 207.885 -136.565 406.635 -135.660 ;
        RECT 420.200 -135.940 440.805 -134.715 ;
        RECT 207.885 -136.700 209.470 -136.565 ;
        RECT 423.060 -137.410 424.285 -135.940 ;
        RECT 126.645 -138.635 424.285 -137.410 ;
        RECT 207.670 -141.160 209.515 -139.275 ;
        RECT 214.270 -140.765 406.635 -139.340 ;
        RECT 207.715 -150.100 209.215 -141.160 ;
        RECT 120.325 -151.600 209.215 -150.100 ;
        RECT 214.270 -152.815 215.695 -140.765 ;
        RECT 119.300 -153.110 215.695 -152.815 ;
        RECT 117.985 -153.715 215.695 -153.110 ;
        RECT 119.300 -154.240 215.695 -153.715 ;
        RECT 63.865 -160.180 441.970 -158.760 ;
        RECT -134.100 -170.785 -132.100 -170.555 ;
        RECT -134.100 -171.375 -132.100 -171.145 ;
        RECT -134.100 -171.965 -132.100 -171.735 ;
        RECT -134.100 -172.555 -132.100 -172.325 ;
        RECT -134.100 -173.145 -132.100 -172.915 ;
        RECT -134.100 -173.735 -132.100 -173.505 ;
        RECT -79.530 -173.630 42.510 -172.680 ;
        RECT -134.100 -174.325 -132.100 -174.095 ;
        RECT -134.100 -174.915 -132.100 -174.685 ;
        RECT -134.100 -175.505 -132.100 -175.275 ;
        RECT -134.100 -176.095 -132.100 -175.865 ;
        RECT -134.100 -176.685 -132.100 -176.455 ;
        RECT -134.100 -177.275 -132.100 -177.045 ;
        RECT -134.100 -177.865 -132.100 -177.635 ;
        RECT -134.100 -178.455 -132.100 -178.225 ;
        RECT -134.100 -179.045 -132.100 -178.815 ;
        RECT -134.100 -179.635 -132.100 -179.405 ;
        RECT -109.740 -179.875 -109.510 -178.875 ;
        RECT -108.760 -179.875 -108.530 -178.875 ;
        RECT -107.780 -179.875 -107.550 -178.875 ;
        RECT -104.090 -179.875 -103.860 -178.875 ;
        RECT -79.530 -179.075 -78.580 -173.630 ;
        RECT -71.745 -175.940 -71.515 -174.940 ;
        RECT -70.765 -175.940 -70.535 -174.940 ;
        RECT -69.785 -175.940 -69.555 -174.940 ;
        RECT -68.635 -176.205 -68.350 -175.030 ;
        RECT -67.560 -175.940 -67.330 -174.940 ;
        RECT -66.580 -175.940 -66.350 -174.940 ;
        RECT -65.600 -175.940 -65.370 -174.940 ;
        RECT -64.505 -175.515 -64.275 -175.015 ;
        RECT -64.015 -175.515 -63.785 -175.015 ;
        RECT -63.525 -175.515 -63.295 -175.015 ;
        RECT -63.035 -175.515 -62.805 -175.015 ;
        RECT -62.545 -175.515 -62.315 -175.015 ;
        RECT -62.055 -175.515 -61.825 -175.015 ;
        RECT -61.565 -175.515 -61.335 -175.015 ;
        RECT -61.075 -175.515 -60.845 -175.015 ;
        RECT -58.245 -175.940 -58.015 -174.940 ;
        RECT -57.265 -175.940 -57.035 -174.940 ;
        RECT -56.285 -175.940 -56.055 -174.940 ;
        RECT -64.490 -176.205 -63.645 -176.155 ;
        RECT -68.635 -176.490 -63.645 -176.205 ;
        RECT -55.135 -176.205 -54.850 -175.030 ;
        RECT -54.060 -175.940 -53.830 -174.940 ;
        RECT -53.080 -175.940 -52.850 -174.940 ;
        RECT -52.100 -175.940 -51.870 -174.940 ;
        RECT -51.005 -175.515 -50.775 -175.015 ;
        RECT -50.515 -175.515 -50.285 -175.015 ;
        RECT -50.025 -175.515 -49.795 -175.015 ;
        RECT -49.535 -175.515 -49.305 -175.015 ;
        RECT -49.045 -175.515 -48.815 -175.015 ;
        RECT -48.555 -175.515 -48.325 -175.015 ;
        RECT -48.065 -175.515 -47.835 -175.015 ;
        RECT -47.575 -175.515 -47.345 -175.015 ;
        RECT -50.990 -176.205 -50.145 -176.155 ;
        RECT -59.430 -176.315 -59.130 -176.285 ;
        RECT -60.605 -176.420 -60.400 -176.415 ;
        RECT -64.490 -176.525 -63.645 -176.490 ;
        RECT -72.235 -177.340 -72.005 -176.840 ;
        RECT -71.745 -177.340 -71.515 -176.840 ;
        RECT -71.255 -177.340 -71.025 -176.840 ;
        RECT -70.765 -177.340 -70.535 -176.840 ;
        RECT -70.275 -177.340 -70.045 -176.840 ;
        RECT -69.785 -177.340 -69.555 -176.840 ;
        RECT -71.065 -178.455 -70.380 -178.155 ;
        RECT -72.805 -178.745 -72.505 -178.510 ;
        RECT -74.115 -179.065 -72.505 -178.745 ;
        RECT -134.100 -180.225 -132.100 -179.995 ;
        RECT -134.100 -180.815 -132.100 -180.585 ;
        RECT -99.745 -180.985 -99.515 -179.485 ;
        RECT -134.100 -181.405 -132.100 -181.175 ;
        RECT -101.780 -181.260 -101.095 -181.175 ;
        RECT -101.920 -181.465 -101.095 -181.260 ;
        RECT -134.100 -181.995 -132.100 -181.765 ;
        RECT -134.100 -182.585 -132.100 -182.355 ;
        RECT -134.100 -183.175 -132.100 -182.945 ;
        RECT -110.230 -183.410 -110.000 -181.910 ;
        RECT -109.740 -183.410 -109.510 -181.910 ;
        RECT -109.250 -183.410 -109.020 -181.910 ;
        RECT -108.680 -183.415 -108.450 -181.915 ;
        RECT -108.190 -183.415 -107.960 -181.915 ;
        RECT -107.700 -183.415 -107.470 -181.915 ;
        RECT -107.135 -183.415 -106.905 -181.915 ;
        RECT -106.645 -183.415 -106.415 -181.915 ;
        RECT -106.155 -183.415 -105.925 -181.915 ;
        RECT -104.580 -183.415 -104.350 -182.415 ;
        RECT -104.090 -182.995 -103.860 -182.415 ;
        RECT -104.090 -183.170 -102.295 -182.995 ;
        RECT -104.090 -183.415 -103.860 -183.170 ;
        RECT -134.100 -183.765 -132.100 -183.535 ;
        RECT -134.100 -184.355 -132.100 -184.125 ;
        RECT -134.100 -184.945 -132.100 -184.715 ;
        RECT -134.100 -185.535 -132.100 -185.305 ;
        RECT -134.100 -186.125 -132.100 -185.895 ;
        RECT -134.100 -186.715 -132.100 -186.485 ;
        RECT -134.100 -187.305 -132.100 -187.075 ;
        RECT -134.100 -187.895 -132.100 -187.665 ;
        RECT -134.100 -188.485 -132.100 -188.255 ;
        RECT -134.100 -189.665 -132.100 -189.435 ;
        RECT -130.785 -190.185 -130.415 -189.610 ;
        RECT -130.785 -190.415 -128.060 -190.185 ;
        RECT -134.100 -190.845 -132.100 -190.615 ;
        RECT -130.785 -191.365 -130.415 -190.415 ;
        RECT -130.785 -191.595 -128.060 -191.365 ;
        RECT -134.100 -192.025 -132.100 -191.795 ;
        RECT -130.785 -192.545 -130.415 -191.595 ;
        RECT -130.785 -192.775 -128.060 -192.545 ;
        RECT -134.100 -193.205 -132.100 -192.975 ;
        RECT -130.785 -193.725 -130.415 -192.775 ;
        RECT -130.785 -193.955 -128.060 -193.725 ;
        RECT -134.100 -194.385 -132.100 -194.155 ;
        RECT -130.785 -194.905 -130.415 -193.955 ;
        RECT -130.785 -195.135 -128.060 -194.905 ;
        RECT -134.100 -195.565 -132.100 -195.335 ;
        RECT -130.785 -196.085 -130.415 -195.135 ;
        RECT -130.785 -196.315 -128.060 -196.085 ;
        RECT -134.100 -196.745 -132.100 -196.515 ;
        RECT -130.785 -197.265 -130.415 -196.315 ;
        RECT -130.785 -197.495 -128.060 -197.265 ;
        RECT -134.100 -197.925 -132.100 -197.695 ;
        RECT -134.100 -198.480 -131.425 -198.285 ;
        RECT -130.785 -198.445 -130.415 -197.495 ;
        RECT -130.785 -198.480 -128.060 -198.445 ;
        RECT -134.100 -198.515 -128.060 -198.480 ;
        RECT -131.655 -198.675 -128.060 -198.515 ;
        RECT -131.655 -198.710 -130.415 -198.675 ;
        RECT -134.100 -199.105 -132.100 -198.875 ;
        RECT -131.655 -199.465 -131.425 -198.710 ;
        RECT -130.785 -199.335 -130.415 -198.710 ;
        RECT -134.100 -199.695 -131.425 -199.465 ;
        RECT -134.100 -200.285 -132.100 -200.055 ;
        RECT -131.655 -200.645 -131.425 -199.695 ;
        RECT -134.100 -200.875 -131.425 -200.645 ;
        RECT -134.100 -201.465 -132.100 -201.235 ;
        RECT -131.655 -201.825 -131.425 -200.875 ;
        RECT -134.100 -202.055 -131.425 -201.825 ;
        RECT -130.785 -200.275 -130.415 -199.640 ;
        RECT -130.785 -200.505 -128.060 -200.275 ;
        RECT -130.785 -201.455 -130.415 -200.505 ;
        RECT -130.785 -201.685 -128.060 -201.455 ;
        RECT -134.100 -202.645 -132.100 -202.415 ;
        RECT -130.785 -202.635 -130.415 -201.685 ;
        RECT -130.785 -202.865 -128.060 -202.635 ;
        RECT -134.100 -203.235 -131.485 -203.005 ;
        RECT -131.715 -203.390 -131.485 -203.235 ;
        RECT -130.785 -203.390 -130.415 -202.865 ;
        RECT -134.100 -203.825 -132.100 -203.595 ;
        RECT -131.715 -203.620 -130.415 -203.390 ;
        RECT -131.715 -204.185 -131.485 -203.620 ;
        RECT -134.100 -204.415 -131.485 -204.185 ;
        RECT -130.785 -203.815 -130.415 -203.620 ;
        RECT -130.785 -204.045 -128.060 -203.815 ;
        RECT -130.785 -204.690 -130.415 -204.045 ;
        RECT -134.100 -205.005 -132.100 -204.775 ;
        RECT -130.785 -205.365 -130.415 -204.995 ;
        RECT -134.100 -205.595 -130.415 -205.365 ;
        RECT -130.785 -205.645 -130.415 -205.595 ;
        RECT -130.785 -205.875 -128.060 -205.645 ;
        RECT -134.100 -206.185 -132.100 -205.955 ;
        RECT -130.785 -206.825 -130.415 -205.875 ;
        RECT -130.785 -207.055 -128.060 -206.825 ;
        RECT -130.785 -207.080 -130.415 -207.055 ;
        RECT -129.885 -214.280 -128.195 -213.945 ;
        RECT -139.045 -215.235 -128.195 -214.280 ;
        RECT -139.045 -216.755 -136.285 -215.235 ;
        RECT -129.885 -215.635 -128.195 -215.235 ;
        RECT -113.370 -227.440 -113.065 -184.605 ;
        RECT -113.715 -227.445 -113.065 -227.440 ;
        RECT -113.715 -227.610 -113.060 -227.445 ;
        RECT -113.710 -228.035 -113.060 -227.610 ;
        RECT -112.800 -228.080 -112.480 -191.965 ;
        RECT -112.810 -228.940 -112.480 -228.080 ;
        RECT -112.915 -228.945 -112.480 -228.940 ;
        RECT -112.075 -214.320 -111.775 -189.810 ;
        RECT -109.455 -190.530 -109.225 -189.030 ;
        RECT -109.945 -193.210 -109.715 -191.715 ;
        RECT -109.950 -193.395 -109.715 -193.210 ;
        RECT -109.455 -193.215 -109.225 -191.715 ;
        RECT -108.965 -193.395 -108.735 -191.715 ;
        RECT -108.475 -193.215 -108.245 -189.030 ;
        RECT -106.410 -189.805 -106.180 -189.025 ;
        RECT -105.430 -189.795 -105.200 -189.025 ;
        RECT -105.920 -189.805 -104.710 -189.795 ;
        RECT -104.450 -189.805 -104.220 -189.025 ;
        RECT -106.410 -190.035 -103.225 -189.805 ;
        RECT -106.410 -190.680 -106.180 -190.180 ;
        RECT -105.920 -190.680 -105.690 -190.035 ;
        RECT -105.430 -190.680 -105.200 -190.180 ;
        RECT -104.940 -190.680 -104.710 -190.035 ;
        RECT -102.470 -190.840 -102.295 -183.170 ;
        RECT -101.920 -185.015 -101.740 -181.465 ;
        RECT -100.235 -183.665 -100.005 -182.170 ;
        RECT -100.240 -183.850 -100.005 -183.665 ;
        RECT -99.745 -183.670 -99.515 -182.170 ;
        RECT -99.255 -183.850 -99.025 -182.170 ;
        RECT -98.765 -183.670 -98.535 -179.485 ;
        RECT -96.700 -180.260 -96.470 -179.480 ;
        RECT -95.720 -180.250 -95.490 -179.480 ;
        RECT -96.210 -180.260 -95.000 -180.250 ;
        RECT -94.740 -180.260 -94.510 -179.480 ;
        RECT -81.435 -179.640 -78.050 -179.075 ;
        RECT -96.700 -180.490 -93.515 -180.260 ;
        RECT -96.700 -181.135 -96.470 -180.635 ;
        RECT -96.210 -181.135 -95.980 -180.490 ;
        RECT -95.720 -181.135 -95.490 -180.635 ;
        RECT -95.230 -181.135 -95.000 -180.490 ;
        RECT -93.100 -180.615 -92.370 -180.325 ;
        RECT -93.100 -180.745 -92.695 -180.615 ;
        RECT -94.660 -180.920 -92.695 -180.745 ;
        RECT -98.275 -183.850 -98.045 -182.170 ;
        RECT -100.240 -184.085 -98.045 -183.850 ;
        RECT -101.930 -185.675 -101.665 -185.015 ;
        RECT -94.660 -186.270 -94.485 -180.920 ;
        RECT -92.060 -181.430 -89.865 -181.195 ;
        RECT -92.060 -181.615 -91.825 -181.430 ;
        RECT -92.055 -183.110 -91.825 -181.615 ;
        RECT -91.565 -183.110 -91.335 -181.610 ;
        RECT -91.075 -183.110 -90.845 -181.430 ;
        RECT -93.330 -183.590 -92.345 -183.320 ;
        RECT -102.140 -186.445 -94.485 -186.270 ;
        RECT -102.140 -190.185 -101.965 -186.445 ;
        RECT -100.590 -189.555 -100.360 -188.555 ;
        RECT -99.610 -189.555 -99.380 -188.555 ;
        RECT -98.630 -189.555 -98.400 -188.555 ;
        RECT -94.940 -189.555 -94.710 -188.555 ;
        RECT -102.140 -190.415 -101.720 -190.185 ;
        RECT -107.985 -193.395 -107.755 -191.715 ;
        RECT -103.565 -192.010 -103.275 -191.325 ;
        RECT -102.495 -191.525 -102.205 -190.840 ;
        RECT -102.010 -190.870 -101.720 -190.415 ;
        RECT -92.615 -190.610 -92.345 -183.590 ;
        RECT -91.565 -185.795 -91.335 -184.295 ;
        RECT -90.585 -185.795 -90.355 -181.610 ;
        RECT -90.095 -183.110 -89.865 -181.430 ;
        RECT -84.330 -181.680 -84.100 -180.180 ;
        RECT -83.840 -181.680 -83.610 -180.180 ;
        RECT -83.350 -181.680 -83.120 -180.180 ;
        RECT -82.140 -181.680 -81.910 -180.180 ;
        RECT -81.650 -181.680 -81.420 -180.180 ;
        RECT -84.825 -182.170 -79.725 -181.845 ;
        RECT -80.050 -182.585 -79.725 -182.170 ;
        RECT -80.080 -182.945 -79.555 -182.585 ;
        RECT -88.520 -184.645 -88.290 -184.145 ;
        RECT -88.030 -184.790 -87.800 -184.145 ;
        RECT -87.540 -184.645 -87.310 -184.145 ;
        RECT -87.050 -184.790 -86.820 -184.145 ;
        RECT -88.520 -185.020 -85.335 -184.790 ;
        RECT -88.520 -185.800 -88.290 -185.020 ;
        RECT -88.030 -185.030 -86.820 -185.020 ;
        RECT -87.540 -185.800 -87.310 -185.030 ;
        RECT -86.560 -185.800 -86.330 -185.020 ;
        RECT -84.330 -186.240 -84.100 -183.240 ;
        RECT -83.275 -186.240 -83.045 -183.240 ;
        RECT -82.785 -186.240 -82.555 -183.240 ;
        RECT -82.295 -186.240 -82.065 -183.240 ;
        RECT -81.235 -186.240 -81.005 -183.240 ;
        RECT -92.865 -191.360 -92.215 -190.610 ;
        RECT -91.435 -190.720 -91.205 -189.440 ;
        RECT -90.455 -190.710 -90.225 -189.440 ;
        RECT -90.945 -190.720 -89.735 -190.710 ;
        RECT -89.475 -190.720 -89.245 -189.440 ;
        RECT -86.570 -190.295 -86.340 -188.795 ;
        RECT -91.435 -190.950 -88.250 -190.720 ;
        RECT -87.540 -190.815 -86.745 -190.525 ;
        RECT -101.080 -193.090 -100.850 -191.590 ;
        RECT -100.590 -193.090 -100.360 -191.590 ;
        RECT -100.100 -193.090 -99.870 -191.590 ;
        RECT -99.530 -193.095 -99.300 -191.595 ;
        RECT -99.040 -193.095 -98.810 -191.595 ;
        RECT -98.550 -193.095 -98.320 -191.595 ;
        RECT -97.985 -193.095 -97.755 -191.595 ;
        RECT -97.495 -193.095 -97.265 -191.595 ;
        RECT -97.005 -193.095 -96.775 -191.595 ;
        RECT -91.435 -192.090 -91.205 -191.090 ;
        RECT -90.945 -192.090 -90.715 -190.950 ;
        RECT -90.455 -192.090 -90.225 -191.090 ;
        RECT -89.965 -192.090 -89.735 -190.950 ;
        RECT -87.410 -191.090 -87.140 -190.815 ;
        RECT -88.780 -191.360 -87.140 -191.090 ;
        RECT -95.430 -193.095 -95.200 -192.095 ;
        RECT -94.940 -193.095 -94.710 -192.095 ;
        RECT -88.780 -192.810 -88.510 -191.360 ;
        RECT -93.995 -193.080 -88.510 -192.810 ;
        RECT -87.060 -192.975 -86.830 -191.480 ;
        RECT -109.950 -193.630 -107.755 -193.395 ;
        RECT -93.935 -196.650 -92.735 -193.080 ;
        RECT -87.065 -193.160 -86.830 -192.975 ;
        RECT -86.570 -192.980 -86.340 -191.480 ;
        RECT -86.080 -193.160 -85.850 -191.480 ;
        RECT -85.590 -192.980 -85.360 -188.795 ;
        RECT -83.525 -189.570 -83.295 -188.790 ;
        RECT -82.545 -189.560 -82.315 -188.790 ;
        RECT -83.035 -189.570 -81.825 -189.560 ;
        RECT -81.565 -189.570 -81.335 -188.790 ;
        RECT -83.525 -189.800 -80.340 -189.570 ;
        RECT -83.525 -190.445 -83.295 -189.945 ;
        RECT -83.035 -190.445 -82.805 -189.800 ;
        RECT -82.545 -190.445 -82.315 -189.945 ;
        RECT -82.055 -190.445 -81.825 -189.800 ;
        RECT -78.615 -190.620 -78.050 -179.640 ;
        RECT -74.115 -188.645 -73.795 -179.065 ;
        RECT -72.805 -179.195 -72.505 -179.065 ;
        RECT -70.990 -179.545 -70.515 -178.455 ;
        RECT -68.940 -179.045 -68.640 -176.710 ;
        RECT -61.080 -176.720 -60.395 -176.420 ;
        RECT -59.430 -176.615 -58.715 -176.315 ;
        RECT -55.135 -176.490 -50.145 -176.205 ;
        RECT -50.990 -176.525 -50.145 -176.490 ;
        RECT -68.050 -177.340 -67.820 -176.840 ;
        RECT -67.560 -177.340 -67.330 -176.840 ;
        RECT -67.070 -177.340 -66.840 -176.840 ;
        RECT -66.580 -177.340 -66.350 -176.840 ;
        RECT -66.090 -177.340 -65.860 -176.840 ;
        RECT -65.600 -177.340 -65.370 -176.840 ;
        RECT -64.505 -177.590 -64.275 -177.090 ;
        RECT -64.015 -177.590 -63.785 -177.090 ;
        RECT -63.525 -177.590 -63.295 -177.090 ;
        RECT -63.035 -177.590 -62.805 -177.090 ;
        RECT -62.545 -177.590 -62.315 -177.090 ;
        RECT -62.055 -177.590 -61.825 -177.090 ;
        RECT -61.565 -177.590 -61.335 -177.090 ;
        RECT -61.075 -177.590 -60.845 -177.090 ;
        RECT -69.120 -179.345 -68.460 -179.045 ;
        RECT -60.605 -179.145 -60.400 -176.720 ;
        RECT -60.255 -178.900 -59.570 -178.600 ;
        RECT -68.055 -179.385 -60.400 -179.145 ;
        RECT -71.110 -179.845 -70.450 -179.545 ;
        RECT -72.235 -180.630 -72.005 -180.130 ;
        RECT -71.745 -180.630 -71.515 -180.130 ;
        RECT -71.255 -180.630 -71.025 -180.130 ;
        RECT -70.765 -180.630 -70.535 -180.130 ;
        RECT -70.275 -180.630 -70.045 -180.130 ;
        RECT -69.785 -180.630 -69.555 -180.130 ;
        RECT -68.055 -180.155 -67.815 -179.385 ;
        RECT -68.045 -180.380 -67.815 -180.155 ;
        RECT -67.555 -180.380 -67.325 -179.880 ;
        RECT -67.095 -179.975 -66.790 -179.385 ;
        RECT -67.065 -180.380 -66.835 -179.975 ;
        RECT -66.575 -180.380 -66.345 -179.880 ;
        RECT -66.115 -179.985 -65.810 -179.385 ;
        RECT -66.085 -180.380 -65.855 -179.985 ;
        RECT -65.595 -180.380 -65.365 -179.880 ;
        RECT -65.160 -179.975 -64.855 -179.385 ;
        RECT -65.105 -180.380 -64.875 -179.975 ;
        RECT -64.615 -180.380 -64.385 -179.880 ;
        RECT -63.520 -180.630 -63.290 -180.130 ;
        RECT -63.030 -180.630 -62.800 -180.130 ;
        RECT -62.540 -180.630 -62.310 -180.130 ;
        RECT -62.050 -180.630 -61.820 -180.130 ;
        RECT -61.560 -180.630 -61.330 -180.130 ;
        RECT -61.070 -180.630 -60.840 -180.130 ;
        RECT -65.245 -180.980 -64.400 -180.945 ;
        RECT -65.245 -181.265 -60.255 -180.980 ;
        RECT -60.010 -181.140 -59.710 -178.900 ;
        RECT -59.430 -180.355 -59.130 -176.615 ;
        RECT -47.635 -176.730 -46.865 -176.430 ;
        RECT -58.735 -177.340 -58.505 -176.840 ;
        RECT -58.245 -177.340 -58.015 -176.840 ;
        RECT -57.755 -177.340 -57.525 -176.840 ;
        RECT -57.265 -177.340 -57.035 -176.840 ;
        RECT -56.775 -177.340 -56.545 -176.840 ;
        RECT -56.285 -177.340 -56.055 -176.840 ;
        RECT -58.080 -178.485 -57.395 -178.185 ;
        RECT -58.025 -179.525 -57.550 -178.485 ;
        RECT -55.380 -178.605 -55.080 -176.785 ;
        RECT -54.550 -177.340 -54.320 -176.840 ;
        RECT -54.060 -177.340 -53.830 -176.840 ;
        RECT -53.570 -177.340 -53.340 -176.840 ;
        RECT -53.080 -177.340 -52.850 -176.840 ;
        RECT -52.590 -177.340 -52.360 -176.840 ;
        RECT -52.100 -177.340 -51.870 -176.840 ;
        RECT -51.005 -177.590 -50.775 -177.090 ;
        RECT -50.515 -177.590 -50.285 -177.090 ;
        RECT -50.025 -177.590 -49.795 -177.090 ;
        RECT -49.535 -177.590 -49.305 -177.090 ;
        RECT -49.045 -177.590 -48.815 -177.090 ;
        RECT -48.555 -177.590 -48.325 -177.090 ;
        RECT -48.065 -177.590 -47.835 -177.090 ;
        RECT -47.575 -177.590 -47.345 -177.090 ;
        RECT -47.095 -178.105 -46.865 -176.730 ;
        RECT -50.960 -178.330 -46.865 -178.105 ;
        RECT -50.960 -178.335 -46.905 -178.330 ;
        RECT -55.525 -178.905 -54.865 -178.605 ;
        RECT -50.960 -179.165 -50.730 -178.335 ;
        RECT -44.890 -178.485 -44.230 -178.185 ;
        RECT -44.805 -178.810 -44.330 -178.485 ;
        RECT -42.130 -178.810 -41.655 -173.630 ;
        RECT -40.915 -177.990 -40.685 -174.990 ;
        RECT -39.855 -177.990 -39.625 -174.990 ;
        RECT -39.365 -177.990 -39.135 -174.990 ;
        RECT -38.875 -177.990 -38.645 -174.990 ;
        RECT -37.820 -177.990 -37.590 -174.990 ;
        RECT -33.765 -176.970 -33.535 -175.970 ;
        RECT -33.275 -176.970 -33.045 -175.970 ;
        RECT -32.785 -176.970 -32.555 -175.970 ;
        RECT -32.185 -176.970 -31.955 -175.970 ;
        RECT -31.695 -176.970 -31.465 -175.970 ;
        RECT -31.205 -176.970 -30.975 -175.970 ;
        RECT -29.395 -176.970 -29.165 -175.970 ;
        RECT -28.415 -176.970 -28.185 -175.970 ;
        RECT -26.865 -176.970 -26.635 -175.970 ;
        RECT -25.320 -176.970 -25.090 -175.970 ;
        RECT -21.265 -176.970 -21.035 -175.970 ;
        RECT -20.775 -176.970 -20.545 -175.970 ;
        RECT -20.285 -176.970 -20.055 -175.970 ;
        RECT -19.685 -176.970 -19.455 -175.970 ;
        RECT -19.195 -176.970 -18.965 -175.970 ;
        RECT -18.705 -176.970 -18.475 -175.970 ;
        RECT -16.895 -176.970 -16.665 -175.970 ;
        RECT -15.915 -176.970 -15.685 -175.970 ;
        RECT -14.365 -176.970 -14.135 -175.970 ;
        RECT -12.820 -176.970 -12.590 -175.970 ;
        RECT -8.765 -176.970 -8.535 -175.970 ;
        RECT -8.275 -176.970 -8.045 -175.970 ;
        RECT -7.785 -176.970 -7.555 -175.970 ;
        RECT -7.185 -176.970 -6.955 -175.970 ;
        RECT -6.695 -176.970 -6.465 -175.970 ;
        RECT -6.205 -176.970 -5.975 -175.970 ;
        RECT -4.395 -176.970 -4.165 -175.970 ;
        RECT -3.415 -176.970 -3.185 -175.970 ;
        RECT -1.865 -176.970 -1.635 -175.970 ;
        RECT -0.320 -176.970 -0.090 -175.970 ;
        RECT 3.735 -176.970 3.965 -175.970 ;
        RECT 4.225 -176.970 4.455 -175.970 ;
        RECT 4.715 -176.970 4.945 -175.970 ;
        RECT 5.315 -176.970 5.545 -175.970 ;
        RECT 5.805 -176.970 6.035 -175.970 ;
        RECT 6.295 -176.970 6.525 -175.970 ;
        RECT 8.105 -176.970 8.335 -175.970 ;
        RECT 9.085 -176.970 9.315 -175.970 ;
        RECT 10.635 -176.970 10.865 -175.970 ;
        RECT 12.180 -176.970 12.410 -175.970 ;
        RECT 16.235 -176.970 16.465 -175.970 ;
        RECT 16.725 -176.970 16.955 -175.970 ;
        RECT 17.215 -176.970 17.445 -175.970 ;
        RECT 17.815 -176.970 18.045 -175.970 ;
        RECT 18.305 -176.970 18.535 -175.970 ;
        RECT 18.795 -176.970 19.025 -175.970 ;
        RECT 20.605 -176.970 20.835 -175.970 ;
        RECT 21.585 -176.970 21.815 -175.970 ;
        RECT 23.135 -176.970 23.365 -175.970 ;
        RECT 24.680 -176.970 24.910 -175.970 ;
        RECT 31.235 -176.970 31.465 -175.970 ;
        RECT 31.725 -176.970 31.955 -175.970 ;
        RECT 32.215 -176.970 32.445 -175.970 ;
        RECT 32.815 -176.970 33.045 -175.970 ;
        RECT 33.305 -176.970 33.535 -175.970 ;
        RECT 33.795 -176.970 34.025 -175.970 ;
        RECT 35.605 -176.970 35.835 -175.970 ;
        RECT 36.585 -176.970 36.815 -175.970 ;
        RECT 38.135 -176.970 38.365 -175.970 ;
        RECT 39.680 -176.970 39.910 -175.970 ;
        RECT -27.950 -177.610 -27.255 -177.520 ;
        RECT -24.875 -177.610 -24.180 -177.550 ;
        RECT -15.450 -177.610 -14.755 -177.520 ;
        RECT -12.375 -177.610 -11.680 -177.550 ;
        RECT -2.950 -177.610 -2.255 -177.520 ;
        RECT 0.125 -177.610 0.820 -177.550 ;
        RECT 9.550 -177.610 10.245 -177.520 ;
        RECT 12.625 -177.610 13.320 -177.550 ;
        RECT 22.050 -177.610 22.745 -177.520 ;
        RECT 25.125 -177.610 25.820 -177.550 ;
        RECT 37.050 -177.610 37.745 -177.520 ;
        RECT 40.125 -177.610 40.820 -177.550 ;
        RECT 43.630 -177.610 44.630 -175.850 ;
        RECT -33.740 -177.805 -33.045 -177.740 ;
        RECT -27.950 -177.750 -23.425 -177.610 ;
        RECT -27.950 -177.790 -27.255 -177.750 ;
        RECT -33.740 -177.945 -31.970 -177.805 ;
        RECT -24.875 -177.820 -24.180 -177.750 ;
        RECT -33.740 -178.010 -33.045 -177.945 ;
        RECT -54.530 -179.395 -50.730 -179.165 ;
        RECT -46.505 -179.335 -45.845 -179.035 ;
        RECT -44.805 -179.285 -41.655 -178.810 ;
        RECT -58.115 -179.825 -57.430 -179.525 ;
        RECT -54.530 -179.880 -54.300 -179.395 ;
        RECT -53.555 -179.880 -53.345 -179.395 ;
        RECT -52.580 -179.880 -52.370 -179.395 ;
        RECT -51.600 -179.880 -51.390 -179.395 ;
        RECT -59.435 -180.580 -59.130 -180.355 ;
        RECT -59.435 -181.015 -59.135 -180.580 ;
        RECT -58.735 -180.630 -58.505 -180.130 ;
        RECT -58.245 -180.630 -58.015 -180.130 ;
        RECT -57.755 -180.630 -57.525 -180.130 ;
        RECT -57.265 -180.630 -57.035 -180.130 ;
        RECT -56.775 -180.630 -56.545 -180.130 ;
        RECT -56.285 -180.630 -56.055 -180.130 ;
        RECT -54.545 -180.380 -54.300 -179.880 ;
        RECT -54.055 -180.380 -53.825 -179.880 ;
        RECT -53.565 -180.380 -53.335 -179.880 ;
        RECT -53.075 -180.380 -52.845 -179.880 ;
        RECT -52.585 -180.380 -52.355 -179.880 ;
        RECT -52.095 -180.380 -51.865 -179.880 ;
        RECT -51.605 -180.380 -51.375 -179.880 ;
        RECT -51.115 -180.380 -50.885 -179.880 ;
        RECT -50.020 -180.630 -49.790 -180.130 ;
        RECT -49.530 -180.630 -49.300 -180.130 ;
        RECT -49.040 -180.630 -48.810 -180.130 ;
        RECT -48.550 -180.630 -48.320 -180.130 ;
        RECT -48.060 -180.630 -47.830 -180.130 ;
        RECT -47.570 -180.630 -47.340 -180.130 ;
        RECT -46.340 -180.475 -46.050 -179.335 ;
        RECT -44.805 -179.530 -44.330 -179.285 ;
        RECT -44.980 -179.830 -44.295 -179.530 ;
        RECT -51.745 -180.980 -50.900 -180.945 ;
        RECT -65.245 -181.315 -64.400 -181.265 ;
        RECT -72.235 -182.530 -72.005 -181.530 ;
        RECT -71.255 -182.530 -71.025 -181.530 ;
        RECT -70.275 -182.530 -70.045 -181.530 ;
        RECT -68.045 -182.295 -67.815 -181.955 ;
        RECT -68.045 -182.455 -67.790 -182.295 ;
        RECT -67.555 -182.455 -67.325 -181.955 ;
        RECT -67.065 -182.170 -66.835 -181.955 ;
        RECT -68.040 -182.870 -67.790 -182.455 ;
        RECT -67.085 -182.870 -66.830 -182.170 ;
        RECT -66.575 -182.455 -66.345 -181.955 ;
        RECT -66.085 -182.265 -65.855 -181.955 ;
        RECT -66.085 -182.870 -65.830 -182.265 ;
        RECT -65.595 -182.455 -65.365 -181.955 ;
        RECT -65.105 -182.265 -64.875 -181.955 ;
        RECT -65.115 -182.870 -64.860 -182.265 ;
        RECT -64.615 -182.455 -64.385 -181.955 ;
        RECT -63.520 -182.530 -63.290 -181.530 ;
        RECT -62.540 -182.530 -62.310 -181.530 ;
        RECT -61.560 -182.530 -61.330 -181.530 ;
        RECT -60.540 -182.440 -60.255 -181.265 ;
        RECT -51.745 -181.265 -46.755 -180.980 ;
        RECT -46.350 -181.135 -46.050 -180.475 ;
        RECT -45.610 -180.630 -45.380 -180.130 ;
        RECT -45.120 -180.630 -44.890 -180.130 ;
        RECT -44.630 -180.630 -44.400 -180.130 ;
        RECT -44.140 -180.630 -43.910 -180.130 ;
        RECT -43.650 -180.630 -43.420 -180.130 ;
        RECT -43.160 -180.630 -42.930 -180.130 ;
        RECT -51.745 -181.315 -50.900 -181.265 ;
        RECT -58.735 -182.530 -58.505 -181.530 ;
        RECT -57.755 -182.530 -57.525 -181.530 ;
        RECT -56.775 -182.530 -56.545 -181.530 ;
        RECT -54.545 -182.455 -54.315 -181.955 ;
        RECT -54.055 -182.455 -53.825 -181.955 ;
        RECT -53.565 -182.455 -53.335 -181.955 ;
        RECT -53.075 -182.455 -52.845 -181.955 ;
        RECT -52.585 -182.455 -52.355 -181.955 ;
        RECT -52.095 -182.455 -51.865 -181.955 ;
        RECT -51.605 -182.455 -51.375 -181.955 ;
        RECT -51.115 -182.455 -50.885 -181.955 ;
        RECT -50.020 -182.530 -49.790 -181.530 ;
        RECT -49.040 -182.530 -48.810 -181.530 ;
        RECT -48.060 -182.530 -47.830 -181.530 ;
        RECT -47.040 -182.870 -46.755 -181.265 ;
        RECT -45.610 -182.530 -45.380 -181.530 ;
        RECT -44.630 -182.530 -44.400 -181.530 ;
        RECT -43.650 -182.530 -43.420 -181.530 ;
        RECT -68.040 -183.155 -46.755 -182.870 ;
        RECT -42.130 -183.955 -41.655 -179.285 ;
        RECT -40.500 -181.050 -40.270 -179.550 ;
        RECT -40.010 -181.050 -39.780 -179.550 ;
        RECT -38.800 -181.050 -38.570 -179.550 ;
        RECT -38.310 -181.050 -38.080 -179.550 ;
        RECT -37.820 -181.050 -37.590 -179.550 ;
        RECT -56.490 -184.520 -41.650 -183.955 ;
        RECT -67.115 -186.310 -64.920 -186.075 ;
        RECT -67.115 -186.495 -66.880 -186.310 ;
        RECT -67.110 -187.990 -66.880 -186.495 ;
        RECT -66.620 -187.990 -66.390 -186.490 ;
        RECT -66.130 -187.990 -65.900 -186.310 ;
        RECT -69.805 -188.645 -68.875 -188.435 ;
        RECT -74.115 -188.965 -68.875 -188.645 ;
        RECT -69.805 -189.205 -68.875 -188.965 ;
        RECT -81.590 -191.185 -78.050 -190.620 ;
        RECT -66.620 -190.675 -66.390 -189.175 ;
        RECT -65.640 -190.675 -65.410 -186.490 ;
        RECT -65.150 -187.990 -64.920 -186.310 ;
        RECT -59.385 -186.560 -59.155 -185.060 ;
        RECT -58.895 -186.560 -58.665 -185.060 ;
        RECT -58.405 -186.560 -58.175 -185.060 ;
        RECT -57.195 -186.560 -56.965 -185.060 ;
        RECT -56.705 -186.560 -56.475 -185.060 ;
        RECT -59.880 -187.050 -54.780 -186.725 ;
        RECT -55.105 -187.465 -54.780 -187.050 ;
        RECT -55.135 -187.825 -54.610 -187.465 ;
        RECT -63.575 -189.525 -63.345 -189.025 ;
        RECT -63.085 -189.670 -62.855 -189.025 ;
        RECT -62.595 -189.525 -62.365 -189.025 ;
        RECT -62.105 -189.670 -61.875 -189.025 ;
        RECT -63.575 -189.900 -60.390 -189.670 ;
        RECT -63.575 -190.680 -63.345 -189.900 ;
        RECT -63.085 -189.910 -61.875 -189.900 ;
        RECT -62.595 -190.680 -62.365 -189.910 ;
        RECT -61.615 -190.680 -61.385 -189.900 ;
        RECT -59.385 -191.120 -59.155 -188.120 ;
        RECT -58.330 -191.120 -58.100 -188.120 ;
        RECT -57.840 -191.120 -57.610 -188.120 ;
        RECT -57.350 -191.120 -57.120 -188.120 ;
        RECT -56.290 -191.120 -56.060 -188.120 ;
        RECT -85.100 -193.160 -84.870 -191.480 ;
        RECT -87.065 -193.395 -84.870 -193.160 ;
        RECT -82.005 -194.940 -80.665 -193.615 ;
        RECT -81.760 -197.715 -80.820 -194.940 ;
        RECT -81.980 -199.040 -80.640 -197.715 ;
        RECT -78.615 -204.075 -78.050 -191.185 ;
        RECT -66.490 -195.600 -66.260 -194.320 ;
        RECT -65.510 -195.590 -65.280 -194.320 ;
        RECT -66.000 -195.600 -64.790 -195.590 ;
        RECT -64.530 -195.600 -64.300 -194.320 ;
        RECT -61.625 -195.175 -61.395 -193.675 ;
        RECT -81.435 -204.640 -78.050 -204.075 ;
        RECT -109.130 -208.000 -108.900 -205.000 ;
        RECT -108.070 -208.000 -107.840 -205.000 ;
        RECT -107.580 -208.000 -107.350 -205.000 ;
        RECT -107.090 -208.000 -106.860 -205.000 ;
        RECT -106.525 -208.000 -106.295 -205.000 ;
        RECT -106.035 -208.000 -105.805 -205.000 ;
        RECT -105.545 -208.000 -105.315 -205.000 ;
        RECT -103.100 -206.645 -102.870 -204.645 ;
        RECT -102.045 -206.645 -101.815 -204.645 ;
        RECT -101.555 -206.645 -101.325 -204.645 ;
        RECT -101.065 -206.645 -100.835 -204.645 ;
        RECT -98.575 -206.650 -98.345 -204.650 ;
        RECT -97.520 -206.650 -97.290 -204.650 ;
        RECT -97.030 -206.650 -96.800 -204.650 ;
        RECT -96.540 -206.650 -96.310 -204.650 ;
        RECT -92.060 -206.430 -89.865 -206.195 ;
        RECT -92.060 -206.615 -91.825 -206.430 ;
        RECT -99.880 -207.460 -99.590 -206.775 ;
        RECT -104.085 -207.645 -103.795 -207.625 ;
        RECT -104.090 -208.310 -103.795 -207.645 ;
        RECT -101.005 -207.885 -100.320 -207.595 ;
        RECT -105.440 -209.630 -104.755 -209.340 ;
        RECT -109.130 -210.820 -108.900 -209.820 ;
        RECT -108.640 -210.820 -108.410 -209.820 ;
        RECT -108.150 -210.820 -107.920 -209.820 ;
        RECT -107.660 -210.820 -107.430 -209.820 ;
        RECT -109.800 -212.050 -105.780 -211.300 ;
        RECT -109.740 -214.110 -109.305 -212.050 ;
        RECT -108.840 -214.110 -108.405 -212.050 ;
        RECT -107.975 -214.110 -107.540 -212.050 ;
        RECT -107.055 -214.110 -106.620 -212.050 ;
        RECT -106.430 -214.110 -105.995 -212.050 ;
        RECT -110.865 -214.320 -105.950 -214.110 ;
        RECT -112.075 -214.620 -105.950 -214.320 ;
        RECT -112.915 -229.560 -112.300 -228.945 ;
        RECT -112.075 -230.780 -111.775 -214.620 ;
        RECT -110.865 -214.685 -105.950 -214.620 ;
        RECT -105.380 -214.620 -104.930 -209.630 ;
        RECT -104.090 -212.395 -103.875 -208.310 ;
        RECT -103.100 -209.105 -102.870 -208.105 ;
        RECT -102.610 -209.105 -102.380 -208.105 ;
        RECT -102.120 -209.105 -101.890 -208.105 ;
        RECT -104.095 -213.080 -103.805 -212.395 ;
        RECT -105.380 -215.070 -103.795 -214.620 ;
        RECT -110.815 -216.550 -110.585 -215.550 ;
        RECT -110.325 -216.550 -110.095 -215.550 ;
        RECT -108.750 -217.050 -108.520 -215.550 ;
        RECT -108.260 -217.050 -108.030 -215.550 ;
        RECT -107.770 -217.050 -107.540 -215.550 ;
        RECT -107.205 -217.050 -106.975 -215.550 ;
        RECT -106.715 -217.050 -106.485 -215.550 ;
        RECT -106.225 -217.050 -105.995 -215.550 ;
        RECT -105.655 -217.055 -105.425 -215.555 ;
        RECT -105.165 -217.055 -104.935 -215.555 ;
        RECT -104.675 -217.055 -104.445 -215.555 ;
        RECT -104.245 -218.010 -103.795 -215.070 ;
        RECT -100.550 -217.735 -100.375 -207.885 ;
        RECT -99.880 -212.790 -99.705 -207.460 ;
        RECT -99.495 -208.320 -99.205 -207.635 ;
        RECT -96.350 -207.890 -95.665 -207.600 ;
        RECT -99.990 -213.475 -99.700 -212.790 ;
        RECT -99.495 -213.175 -99.320 -208.320 ;
        RECT -98.575 -209.110 -98.345 -208.110 ;
        RECT -98.085 -209.110 -97.855 -208.110 ;
        RECT -97.595 -209.110 -97.365 -208.110 ;
        RECT -99.525 -213.860 -99.235 -213.175 ;
        RECT -100.590 -218.420 -100.300 -217.735 ;
        RECT -95.925 -218.165 -95.750 -207.890 ;
        RECT -92.055 -208.110 -91.825 -206.615 ;
        RECT -91.565 -208.110 -91.335 -206.610 ;
        RECT -91.075 -208.110 -90.845 -206.430 ;
        RECT -93.330 -208.590 -92.345 -208.320 ;
        RECT -95.045 -209.380 -94.460 -208.765 ;
        RECT -95.540 -216.405 -95.250 -215.720 ;
        RECT -95.965 -218.850 -95.675 -218.165 ;
        RECT -110.815 -220.090 -110.585 -219.090 ;
        RECT -107.125 -220.090 -106.895 -219.090 ;
        RECT -106.145 -220.090 -105.915 -219.090 ;
        RECT -105.165 -220.090 -104.935 -219.090 ;
        RECT -110.810 -221.445 -110.595 -220.090 ;
        RECT -111.060 -222.025 -110.270 -221.445 ;
        RECT -95.535 -221.585 -95.340 -216.405 ;
        RECT -95.030 -220.700 -94.570 -209.380 ;
        RECT -92.615 -215.610 -92.345 -208.590 ;
        RECT -91.565 -210.795 -91.335 -209.295 ;
        RECT -90.585 -210.795 -90.355 -206.610 ;
        RECT -90.095 -208.110 -89.865 -206.430 ;
        RECT -84.330 -206.680 -84.100 -205.180 ;
        RECT -83.840 -206.680 -83.610 -205.180 ;
        RECT -83.350 -206.680 -83.120 -205.180 ;
        RECT -82.140 -206.680 -81.910 -205.180 ;
        RECT -81.650 -206.680 -81.420 -205.180 ;
        RECT -84.825 -207.170 -79.725 -206.845 ;
        RECT -80.050 -207.585 -79.725 -207.170 ;
        RECT -80.080 -207.945 -79.555 -207.585 ;
        RECT -88.520 -209.645 -88.290 -209.145 ;
        RECT -88.030 -209.790 -87.800 -209.145 ;
        RECT -87.540 -209.645 -87.310 -209.145 ;
        RECT -87.050 -209.790 -86.820 -209.145 ;
        RECT -88.520 -210.020 -85.335 -209.790 ;
        RECT -88.520 -210.800 -88.290 -210.020 ;
        RECT -88.030 -210.030 -86.820 -210.020 ;
        RECT -87.540 -210.800 -87.310 -210.030 ;
        RECT -86.560 -210.800 -86.330 -210.020 ;
        RECT -84.330 -211.240 -84.100 -208.240 ;
        RECT -83.275 -211.240 -83.045 -208.240 ;
        RECT -82.785 -211.240 -82.555 -208.240 ;
        RECT -82.295 -211.240 -82.065 -208.240 ;
        RECT -81.235 -211.240 -81.005 -208.240 ;
        RECT -92.865 -216.360 -92.215 -215.610 ;
        RECT -91.435 -215.720 -91.205 -214.440 ;
        RECT -90.455 -215.710 -90.225 -214.440 ;
        RECT -90.945 -215.720 -89.735 -215.710 ;
        RECT -89.475 -215.720 -89.245 -214.440 ;
        RECT -86.570 -215.295 -86.340 -213.795 ;
        RECT -91.435 -215.950 -88.250 -215.720 ;
        RECT -87.540 -215.815 -86.745 -215.525 ;
        RECT -91.435 -217.090 -91.205 -216.090 ;
        RECT -90.945 -217.090 -90.715 -215.950 ;
        RECT -90.455 -217.090 -90.225 -216.090 ;
        RECT -89.965 -217.090 -89.735 -215.950 ;
        RECT -87.410 -216.090 -87.140 -215.815 ;
        RECT -88.780 -216.360 -87.140 -216.090 ;
        RECT -88.780 -217.810 -88.510 -216.360 ;
        RECT -93.995 -218.080 -88.510 -217.810 ;
        RECT -87.060 -217.975 -86.830 -216.480 ;
        RECT -93.995 -219.430 -93.725 -218.080 ;
        RECT -87.065 -218.160 -86.830 -217.975 ;
        RECT -86.570 -217.980 -86.340 -216.480 ;
        RECT -86.080 -218.160 -85.850 -216.480 ;
        RECT -85.590 -217.980 -85.360 -213.795 ;
        RECT -83.525 -214.570 -83.295 -213.790 ;
        RECT -82.545 -214.560 -82.315 -213.790 ;
        RECT -83.035 -214.570 -81.825 -214.560 ;
        RECT -81.565 -214.570 -81.335 -213.790 ;
        RECT -83.525 -214.800 -80.340 -214.570 ;
        RECT -83.525 -215.445 -83.295 -214.945 ;
        RECT -83.035 -215.445 -82.805 -214.800 ;
        RECT -82.545 -215.445 -82.315 -214.945 ;
        RECT -82.055 -215.445 -81.825 -214.800 ;
        RECT -78.615 -215.620 -78.050 -204.640 ;
        RECT -77.285 -207.600 -76.245 -195.620 ;
        RECT -66.490 -195.830 -63.305 -195.600 ;
        RECT -62.595 -195.695 -61.800 -195.405 ;
        RECT -66.490 -196.970 -66.260 -195.970 ;
        RECT -66.000 -196.970 -65.770 -195.830 ;
        RECT -65.510 -196.970 -65.280 -195.970 ;
        RECT -65.020 -196.970 -64.790 -195.830 ;
        RECT -62.465 -195.970 -62.195 -195.695 ;
        RECT -63.835 -196.240 -62.195 -195.970 ;
        RECT -63.835 -197.690 -63.565 -196.240 ;
        RECT -74.405 -197.960 -63.565 -197.690 ;
        RECT -62.115 -197.855 -61.885 -196.360 ;
        RECT -74.405 -203.380 -74.135 -197.960 ;
        RECT -62.120 -198.040 -61.885 -197.855 ;
        RECT -61.625 -197.860 -61.395 -196.360 ;
        RECT -61.135 -198.040 -60.905 -196.360 ;
        RECT -60.645 -197.860 -60.415 -193.675 ;
        RECT -58.580 -194.450 -58.350 -193.670 ;
        RECT -57.600 -194.440 -57.370 -193.670 ;
        RECT -58.090 -194.450 -56.880 -194.440 ;
        RECT -56.620 -194.450 -56.390 -193.670 ;
        RECT -58.580 -194.680 -55.395 -194.450 ;
        RECT -58.580 -195.325 -58.350 -194.825 ;
        RECT -58.090 -195.325 -57.860 -194.680 ;
        RECT -57.600 -195.325 -57.370 -194.825 ;
        RECT -57.110 -195.325 -56.880 -194.680 ;
        RECT -53.670 -195.500 -53.105 -184.520 ;
        RECT -56.645 -196.065 -53.105 -195.500 ;
        RECT -60.155 -198.040 -59.925 -196.360 ;
        RECT -62.120 -198.275 -59.925 -198.040 ;
        RECT -71.745 -200.575 -71.515 -199.575 ;
        RECT -70.765 -200.575 -70.535 -199.575 ;
        RECT -69.785 -200.575 -69.555 -199.575 ;
        RECT -68.635 -200.840 -68.350 -199.665 ;
        RECT -67.560 -200.575 -67.330 -199.575 ;
        RECT -66.580 -200.575 -66.350 -199.575 ;
        RECT -65.600 -200.575 -65.370 -199.575 ;
        RECT -64.505 -200.150 -64.275 -199.650 ;
        RECT -64.015 -200.150 -63.785 -199.650 ;
        RECT -63.525 -200.150 -63.295 -199.650 ;
        RECT -63.035 -200.150 -62.805 -199.650 ;
        RECT -62.545 -200.150 -62.315 -199.650 ;
        RECT -62.055 -200.150 -61.825 -199.650 ;
        RECT -61.565 -200.150 -61.335 -199.650 ;
        RECT -61.075 -200.150 -60.845 -199.650 ;
        RECT -58.245 -200.575 -58.015 -199.575 ;
        RECT -57.265 -200.575 -57.035 -199.575 ;
        RECT -56.285 -200.575 -56.055 -199.575 ;
        RECT -64.490 -200.840 -63.645 -200.790 ;
        RECT -68.635 -201.125 -63.645 -200.840 ;
        RECT -55.135 -200.840 -54.850 -199.665 ;
        RECT -54.060 -200.575 -53.830 -199.575 ;
        RECT -53.080 -200.575 -52.850 -199.575 ;
        RECT -52.100 -200.575 -51.870 -199.575 ;
        RECT -51.005 -200.150 -50.775 -199.650 ;
        RECT -50.515 -200.150 -50.285 -199.650 ;
        RECT -50.025 -200.150 -49.795 -199.650 ;
        RECT -49.535 -200.150 -49.305 -199.650 ;
        RECT -49.045 -200.150 -48.815 -199.650 ;
        RECT -48.555 -200.150 -48.325 -199.650 ;
        RECT -48.065 -200.150 -47.835 -199.650 ;
        RECT -47.575 -200.150 -47.345 -199.650 ;
        RECT -50.990 -200.840 -50.145 -200.790 ;
        RECT -59.430 -200.950 -59.130 -200.920 ;
        RECT -60.605 -201.055 -60.400 -201.050 ;
        RECT -64.490 -201.160 -63.645 -201.125 ;
        RECT -72.235 -201.975 -72.005 -201.475 ;
        RECT -71.745 -201.975 -71.515 -201.475 ;
        RECT -71.255 -201.975 -71.025 -201.475 ;
        RECT -70.765 -201.975 -70.535 -201.475 ;
        RECT -70.275 -201.975 -70.045 -201.475 ;
        RECT -69.785 -201.975 -69.555 -201.475 ;
        RECT -71.065 -203.090 -70.380 -202.790 ;
        RECT -72.805 -203.380 -72.505 -203.145 ;
        RECT -74.405 -203.700 -72.505 -203.380 ;
        RECT -72.805 -203.830 -72.505 -203.700 ;
        RECT -70.990 -204.180 -70.515 -203.090 ;
        RECT -68.940 -203.680 -68.640 -201.345 ;
        RECT -61.080 -201.355 -60.395 -201.055 ;
        RECT -59.430 -201.250 -58.715 -200.950 ;
        RECT -55.135 -201.125 -50.145 -200.840 ;
        RECT -50.990 -201.160 -50.145 -201.125 ;
        RECT -68.050 -201.975 -67.820 -201.475 ;
        RECT -67.560 -201.975 -67.330 -201.475 ;
        RECT -67.070 -201.975 -66.840 -201.475 ;
        RECT -66.580 -201.975 -66.350 -201.475 ;
        RECT -66.090 -201.975 -65.860 -201.475 ;
        RECT -65.600 -201.975 -65.370 -201.475 ;
        RECT -64.505 -202.225 -64.275 -201.725 ;
        RECT -64.015 -202.225 -63.785 -201.725 ;
        RECT -63.525 -202.225 -63.295 -201.725 ;
        RECT -63.035 -202.225 -62.805 -201.725 ;
        RECT -62.545 -202.225 -62.315 -201.725 ;
        RECT -62.055 -202.225 -61.825 -201.725 ;
        RECT -61.565 -202.225 -61.335 -201.725 ;
        RECT -61.075 -202.225 -60.845 -201.725 ;
        RECT -69.120 -203.980 -68.460 -203.680 ;
        RECT -60.605 -203.780 -60.400 -201.355 ;
        RECT -60.255 -203.535 -59.570 -203.235 ;
        RECT -68.055 -204.020 -60.400 -203.780 ;
        RECT -71.110 -204.480 -70.450 -204.180 ;
        RECT -72.235 -205.265 -72.005 -204.765 ;
        RECT -71.745 -205.265 -71.515 -204.765 ;
        RECT -71.255 -205.265 -71.025 -204.765 ;
        RECT -70.765 -205.265 -70.535 -204.765 ;
        RECT -70.275 -205.265 -70.045 -204.765 ;
        RECT -69.785 -205.265 -69.555 -204.765 ;
        RECT -68.055 -204.790 -67.815 -204.020 ;
        RECT -68.045 -205.015 -67.815 -204.790 ;
        RECT -67.555 -205.015 -67.325 -204.515 ;
        RECT -67.095 -204.610 -66.790 -204.020 ;
        RECT -67.065 -205.015 -66.835 -204.610 ;
        RECT -66.575 -205.015 -66.345 -204.515 ;
        RECT -66.115 -204.620 -65.810 -204.020 ;
        RECT -66.085 -205.015 -65.855 -204.620 ;
        RECT -65.595 -205.015 -65.365 -204.515 ;
        RECT -65.160 -204.610 -64.855 -204.020 ;
        RECT -65.105 -205.015 -64.875 -204.610 ;
        RECT -64.615 -205.015 -64.385 -204.515 ;
        RECT -63.520 -205.265 -63.290 -204.765 ;
        RECT -63.030 -205.265 -62.800 -204.765 ;
        RECT -62.540 -205.265 -62.310 -204.765 ;
        RECT -62.050 -205.265 -61.820 -204.765 ;
        RECT -61.560 -205.265 -61.330 -204.765 ;
        RECT -61.070 -205.265 -60.840 -204.765 ;
        RECT -65.245 -205.615 -64.400 -205.580 ;
        RECT -65.245 -205.900 -60.255 -205.615 ;
        RECT -60.010 -205.775 -59.710 -203.535 ;
        RECT -59.430 -204.990 -59.130 -201.250 ;
        RECT -47.635 -201.365 -46.865 -201.065 ;
        RECT -58.735 -201.975 -58.505 -201.475 ;
        RECT -58.245 -201.975 -58.015 -201.475 ;
        RECT -57.755 -201.975 -57.525 -201.475 ;
        RECT -57.265 -201.975 -57.035 -201.475 ;
        RECT -56.775 -201.975 -56.545 -201.475 ;
        RECT -56.285 -201.975 -56.055 -201.475 ;
        RECT -58.080 -203.120 -57.395 -202.820 ;
        RECT -58.025 -204.160 -57.550 -203.120 ;
        RECT -55.380 -203.240 -55.080 -201.420 ;
        RECT -54.550 -201.975 -54.320 -201.475 ;
        RECT -54.060 -201.975 -53.830 -201.475 ;
        RECT -53.570 -201.975 -53.340 -201.475 ;
        RECT -53.080 -201.975 -52.850 -201.475 ;
        RECT -52.590 -201.975 -52.360 -201.475 ;
        RECT -52.100 -201.975 -51.870 -201.475 ;
        RECT -51.005 -202.225 -50.775 -201.725 ;
        RECT -50.515 -202.225 -50.285 -201.725 ;
        RECT -50.025 -202.225 -49.795 -201.725 ;
        RECT -49.535 -202.225 -49.305 -201.725 ;
        RECT -49.045 -202.225 -48.815 -201.725 ;
        RECT -48.555 -202.225 -48.325 -201.725 ;
        RECT -48.065 -202.225 -47.835 -201.725 ;
        RECT -47.575 -202.225 -47.345 -201.725 ;
        RECT -47.095 -202.740 -46.865 -201.365 ;
        RECT -50.960 -202.965 -46.865 -202.740 ;
        RECT -44.805 -202.820 -44.330 -184.520 ;
        RECT -50.960 -202.970 -46.905 -202.965 ;
        RECT -55.525 -203.540 -54.865 -203.240 ;
        RECT -50.960 -203.800 -50.730 -202.970 ;
        RECT -44.890 -203.120 -44.230 -202.820 ;
        RECT -54.530 -204.030 -50.730 -203.800 ;
        RECT -46.505 -203.970 -45.845 -203.670 ;
        RECT -58.115 -204.460 -57.430 -204.160 ;
        RECT -54.530 -204.515 -54.300 -204.030 ;
        RECT -53.555 -204.515 -53.345 -204.030 ;
        RECT -52.580 -204.515 -52.370 -204.030 ;
        RECT -51.600 -204.515 -51.390 -204.030 ;
        RECT -59.435 -205.215 -59.130 -204.990 ;
        RECT -59.435 -205.650 -59.135 -205.215 ;
        RECT -58.735 -205.265 -58.505 -204.765 ;
        RECT -58.245 -205.265 -58.015 -204.765 ;
        RECT -57.755 -205.265 -57.525 -204.765 ;
        RECT -57.265 -205.265 -57.035 -204.765 ;
        RECT -56.775 -205.265 -56.545 -204.765 ;
        RECT -56.285 -205.265 -56.055 -204.765 ;
        RECT -54.545 -205.015 -54.300 -204.515 ;
        RECT -54.055 -205.015 -53.825 -204.515 ;
        RECT -53.565 -205.015 -53.335 -204.515 ;
        RECT -53.075 -205.015 -52.845 -204.515 ;
        RECT -52.585 -205.015 -52.355 -204.515 ;
        RECT -52.095 -205.015 -51.865 -204.515 ;
        RECT -51.605 -205.015 -51.375 -204.515 ;
        RECT -51.115 -205.015 -50.885 -204.515 ;
        RECT -50.020 -205.265 -49.790 -204.765 ;
        RECT -49.530 -205.265 -49.300 -204.765 ;
        RECT -49.040 -205.265 -48.810 -204.765 ;
        RECT -48.550 -205.265 -48.320 -204.765 ;
        RECT -48.060 -205.265 -47.830 -204.765 ;
        RECT -47.570 -205.265 -47.340 -204.765 ;
        RECT -46.340 -205.110 -46.050 -203.970 ;
        RECT -44.805 -204.165 -44.330 -203.120 ;
        RECT -44.980 -204.465 -44.295 -204.165 ;
        RECT -51.745 -205.615 -50.900 -205.580 ;
        RECT -65.245 -205.950 -64.400 -205.900 ;
        RECT -72.235 -207.165 -72.005 -206.165 ;
        RECT -71.255 -207.165 -71.025 -206.165 ;
        RECT -70.275 -207.165 -70.045 -206.165 ;
        RECT -68.045 -206.930 -67.815 -206.590 ;
        RECT -68.045 -207.090 -67.790 -206.930 ;
        RECT -67.555 -207.090 -67.325 -206.590 ;
        RECT -67.065 -206.805 -66.835 -206.590 ;
        RECT -68.040 -207.505 -67.790 -207.090 ;
        RECT -67.085 -207.505 -66.830 -206.805 ;
        RECT -66.575 -207.090 -66.345 -206.590 ;
        RECT -66.085 -206.900 -65.855 -206.590 ;
        RECT -66.085 -207.505 -65.830 -206.900 ;
        RECT -65.595 -207.090 -65.365 -206.590 ;
        RECT -65.105 -206.900 -64.875 -206.590 ;
        RECT -65.115 -207.505 -64.860 -206.900 ;
        RECT -64.615 -207.090 -64.385 -206.590 ;
        RECT -63.520 -207.165 -63.290 -206.165 ;
        RECT -62.540 -207.165 -62.310 -206.165 ;
        RECT -61.560 -207.165 -61.330 -206.165 ;
        RECT -60.540 -207.075 -60.255 -205.900 ;
        RECT -51.745 -205.900 -46.755 -205.615 ;
        RECT -46.350 -205.770 -46.050 -205.110 ;
        RECT -45.610 -205.265 -45.380 -204.765 ;
        RECT -45.120 -205.265 -44.890 -204.765 ;
        RECT -44.630 -205.265 -44.400 -204.765 ;
        RECT -44.140 -205.265 -43.910 -204.765 ;
        RECT -43.650 -205.265 -43.420 -204.765 ;
        RECT -43.160 -205.265 -42.930 -204.765 ;
        RECT -51.745 -205.950 -50.900 -205.900 ;
        RECT -58.735 -207.165 -58.505 -206.165 ;
        RECT -57.755 -207.165 -57.525 -206.165 ;
        RECT -56.775 -207.165 -56.545 -206.165 ;
        RECT -54.545 -207.090 -54.315 -206.590 ;
        RECT -54.055 -207.090 -53.825 -206.590 ;
        RECT -53.565 -207.090 -53.335 -206.590 ;
        RECT -53.075 -207.090 -52.845 -206.590 ;
        RECT -52.585 -207.090 -52.355 -206.590 ;
        RECT -52.095 -207.090 -51.865 -206.590 ;
        RECT -51.605 -207.090 -51.375 -206.590 ;
        RECT -51.115 -207.090 -50.885 -206.590 ;
        RECT -50.020 -207.165 -49.790 -206.165 ;
        RECT -49.040 -207.165 -48.810 -206.165 ;
        RECT -48.060 -207.165 -47.830 -206.165 ;
        RECT -47.040 -207.505 -46.755 -205.900 ;
        RECT -45.610 -207.165 -45.380 -206.165 ;
        RECT -44.630 -207.165 -44.400 -206.165 ;
        RECT -43.650 -207.165 -43.420 -206.165 ;
        RECT -68.040 -207.790 -46.755 -207.505 ;
        RECT -81.590 -216.185 -78.050 -215.620 ;
        RECT -85.100 -218.160 -84.870 -216.480 ;
        RECT -87.065 -218.395 -84.870 -218.160 ;
        RECT -42.175 -219.310 -41.295 -186.735 ;
        RECT -40.780 -202.660 -40.550 -199.660 ;
        RECT -39.720 -202.660 -39.490 -199.660 ;
        RECT -39.230 -202.660 -39.000 -199.660 ;
        RECT -38.740 -202.660 -38.510 -199.660 ;
        RECT -37.685 -202.660 -37.455 -199.660 ;
        RECT -40.365 -205.720 -40.135 -204.220 ;
        RECT -39.875 -205.720 -39.645 -204.220 ;
        RECT -38.665 -205.720 -38.435 -204.220 ;
        RECT -38.175 -205.720 -37.945 -204.220 ;
        RECT -37.685 -205.720 -37.455 -204.220 ;
        RECT -94.145 -220.110 -93.425 -219.430 ;
        RECT -42.240 -220.165 -41.240 -219.310 ;
        RECT -36.500 -220.600 -35.840 -178.240 ;
        RECT -32.110 -178.670 -31.970 -177.945 ;
        RECT -29.995 -177.935 -29.300 -177.890 ;
        RECT -25.810 -177.935 -25.130 -177.890 ;
        RECT -29.995 -178.075 -25.130 -177.935 ;
        RECT -29.995 -178.160 -29.300 -178.075 ;
        RECT -25.810 -178.120 -25.130 -178.075 ;
        RECT -31.830 -178.305 -31.135 -178.260 ;
        RECT -26.440 -178.295 -25.745 -178.290 ;
        RECT -26.440 -178.305 -23.785 -178.295 ;
        RECT -31.830 -178.435 -23.785 -178.305 ;
        RECT -31.830 -178.445 -25.745 -178.435 ;
        RECT -31.830 -178.530 -31.135 -178.445 ;
        RECT -26.440 -178.560 -25.745 -178.445 ;
        RECT -27.340 -178.670 -26.685 -178.610 ;
        RECT -32.110 -178.810 -26.685 -178.670 ;
        RECT -27.340 -178.840 -26.685 -178.810 ;
        RECT -33.765 -180.000 -33.535 -179.000 ;
        RECT -33.275 -180.000 -33.045 -179.000 ;
        RECT -31.695 -180.000 -31.465 -179.000 ;
        RECT -31.205 -180.000 -30.975 -179.000 ;
        RECT -29.885 -180.000 -29.655 -179.000 ;
        RECT -29.395 -180.000 -29.165 -179.000 ;
        RECT -28.415 -180.000 -28.185 -179.000 ;
        RECT -27.925 -180.000 -27.695 -179.000 ;
        RECT -26.865 -180.000 -26.635 -179.000 ;
        RECT -26.375 -180.000 -26.145 -179.000 ;
        RECT -25.320 -180.000 -25.090 -179.000 ;
        RECT -24.830 -180.000 -24.600 -179.000 ;
        RECT -31.580 -181.715 -31.350 -181.215 ;
        RECT -31.090 -181.715 -30.860 -181.215 ;
        RECT -30.600 -181.715 -30.370 -181.215 ;
        RECT -30.110 -181.715 -29.880 -181.215 ;
        RECT -29.620 -181.715 -29.390 -181.215 ;
        RECT -29.130 -181.715 -28.900 -181.215 ;
        RECT -23.925 -181.630 -23.785 -178.435 ;
        RECT -24.015 -182.310 -23.785 -181.630 ;
        RECT -31.090 -183.615 -30.860 -182.615 ;
        RECT -30.110 -183.615 -29.880 -182.615 ;
        RECT -29.130 -183.615 -28.900 -182.615 ;
        RECT -23.565 -183.790 -23.425 -177.750 ;
        RECT -21.240 -177.805 -20.545 -177.740 ;
        RECT -15.450 -177.750 -10.570 -177.610 ;
        RECT -15.450 -177.790 -14.755 -177.750 ;
        RECT -21.240 -177.945 -19.470 -177.805 ;
        RECT -12.375 -177.820 -11.680 -177.750 ;
        RECT -21.240 -178.010 -20.545 -177.945 ;
        RECT -19.610 -178.670 -19.470 -177.945 ;
        RECT -17.495 -177.935 -16.800 -177.890 ;
        RECT -13.310 -177.935 -12.630 -177.890 ;
        RECT -17.495 -178.075 -12.630 -177.935 ;
        RECT -17.495 -178.160 -16.800 -178.075 ;
        RECT -13.310 -178.120 -12.630 -178.075 ;
        RECT -19.330 -178.305 -18.635 -178.260 ;
        RECT -13.940 -178.295 -13.245 -178.290 ;
        RECT -13.940 -178.305 -11.000 -178.295 ;
        RECT -19.330 -178.435 -11.000 -178.305 ;
        RECT -19.330 -178.445 -13.245 -178.435 ;
        RECT -19.330 -178.530 -18.635 -178.445 ;
        RECT -13.940 -178.560 -13.245 -178.445 ;
        RECT -14.840 -178.670 -14.185 -178.610 ;
        RECT -19.610 -178.810 -14.185 -178.670 ;
        RECT -14.840 -178.840 -14.185 -178.810 ;
        RECT -22.105 -179.835 -21.875 -179.155 ;
        RECT -22.100 -182.685 -21.880 -179.835 ;
        RECT -21.265 -180.000 -21.035 -179.000 ;
        RECT -20.775 -180.000 -20.545 -179.000 ;
        RECT -19.195 -180.000 -18.965 -179.000 ;
        RECT -18.705 -180.000 -18.475 -179.000 ;
        RECT -17.385 -180.000 -17.155 -179.000 ;
        RECT -16.895 -180.000 -16.665 -179.000 ;
        RECT -15.915 -180.000 -15.685 -179.000 ;
        RECT -15.425 -180.000 -15.195 -179.000 ;
        RECT -14.365 -180.000 -14.135 -179.000 ;
        RECT -13.875 -180.000 -13.645 -179.000 ;
        RECT -12.820 -180.000 -12.590 -179.000 ;
        RECT -12.330 -180.000 -12.100 -179.000 ;
        RECT -22.105 -183.365 -21.875 -182.685 ;
        RECT -11.140 -183.455 -11.000 -178.435 ;
        RECT -10.710 -183.040 -10.570 -177.750 ;
        RECT -8.740 -177.805 -8.045 -177.740 ;
        RECT -2.950 -177.750 1.790 -177.610 ;
        RECT -2.950 -177.790 -2.255 -177.750 ;
        RECT -8.740 -177.945 -6.970 -177.805 ;
        RECT 0.125 -177.820 0.820 -177.750 ;
        RECT -8.740 -178.010 -8.045 -177.945 ;
        RECT -7.110 -178.670 -6.970 -177.945 ;
        RECT -4.995 -177.935 -4.300 -177.890 ;
        RECT -0.810 -177.935 -0.130 -177.890 ;
        RECT -4.995 -178.075 -0.130 -177.935 ;
        RECT -4.995 -178.160 -4.300 -178.075 ;
        RECT -0.810 -178.120 -0.130 -178.075 ;
        RECT -6.830 -178.305 -6.135 -178.260 ;
        RECT -1.440 -178.295 -0.745 -178.290 ;
        RECT -1.440 -178.305 1.420 -178.295 ;
        RECT -6.830 -178.435 1.420 -178.305 ;
        RECT -6.830 -178.445 -0.745 -178.435 ;
        RECT -6.830 -178.530 -6.135 -178.445 ;
        RECT -1.440 -178.560 -0.745 -178.445 ;
        RECT -2.340 -178.670 -1.685 -178.610 ;
        RECT -7.110 -178.810 -1.685 -178.670 ;
        RECT -2.340 -178.840 -1.685 -178.810 ;
        RECT -9.365 -179.855 -9.135 -179.175 ;
        RECT -9.360 -181.040 -9.140 -179.855 ;
        RECT -8.765 -180.000 -8.535 -179.000 ;
        RECT -8.275 -180.000 -8.045 -179.000 ;
        RECT -6.695 -180.000 -6.465 -179.000 ;
        RECT -6.205 -180.000 -5.975 -179.000 ;
        RECT -4.885 -180.000 -4.655 -179.000 ;
        RECT -4.395 -180.000 -4.165 -179.000 ;
        RECT -3.415 -180.000 -3.185 -179.000 ;
        RECT -2.925 -180.000 -2.695 -179.000 ;
        RECT -1.865 -180.000 -1.635 -179.000 ;
        RECT -1.375 -180.000 -1.145 -179.000 ;
        RECT -0.320 -180.000 -0.090 -179.000 ;
        RECT 0.170 -180.000 0.400 -179.000 ;
        RECT -8.540 -181.040 -7.860 -181.035 ;
        RECT -9.365 -181.260 -7.860 -181.040 ;
        RECT -8.540 -181.265 -7.860 -181.260 ;
        RECT 1.280 -182.760 1.420 -178.435 ;
        RECT 1.650 -182.475 1.790 -177.750 ;
        RECT 3.760 -177.805 4.455 -177.740 ;
        RECT 9.550 -177.750 14.165 -177.610 ;
        RECT 9.550 -177.790 10.245 -177.750 ;
        RECT 3.760 -177.945 5.530 -177.805 ;
        RECT 12.625 -177.820 13.320 -177.750 ;
        RECT 3.760 -178.010 4.455 -177.945 ;
        RECT 5.390 -178.670 5.530 -177.945 ;
        RECT 7.505 -177.935 8.200 -177.890 ;
        RECT 11.690 -177.935 12.370 -177.890 ;
        RECT 7.505 -178.075 12.370 -177.935 ;
        RECT 7.505 -178.160 8.200 -178.075 ;
        RECT 11.690 -178.120 12.370 -178.075 ;
        RECT 5.670 -178.305 6.365 -178.260 ;
        RECT 11.060 -178.295 11.755 -178.290 ;
        RECT 11.060 -178.305 13.750 -178.295 ;
        RECT 5.670 -178.435 13.750 -178.305 ;
        RECT 5.670 -178.445 11.755 -178.435 ;
        RECT 5.670 -178.530 6.365 -178.445 ;
        RECT 11.060 -178.560 11.755 -178.445 ;
        RECT 10.160 -178.670 10.815 -178.610 ;
        RECT 5.390 -178.810 10.815 -178.670 ;
        RECT 10.160 -178.840 10.815 -178.810 ;
        RECT 3.035 -179.855 3.265 -179.175 ;
        RECT 3.040 -181.105 3.260 -179.855 ;
        RECT 3.735 -180.000 3.965 -179.000 ;
        RECT 4.225 -180.000 4.455 -179.000 ;
        RECT 5.805 -180.000 6.035 -179.000 ;
        RECT 6.295 -180.000 6.525 -179.000 ;
        RECT 7.615 -180.000 7.845 -179.000 ;
        RECT 8.105 -180.000 8.335 -179.000 ;
        RECT 9.085 -180.000 9.315 -179.000 ;
        RECT 9.575 -180.000 9.805 -179.000 ;
        RECT 10.635 -180.000 10.865 -179.000 ;
        RECT 11.125 -180.000 11.355 -179.000 ;
        RECT 12.180 -180.000 12.410 -179.000 ;
        RECT 12.670 -180.000 12.900 -179.000 ;
        RECT 3.945 -181.105 4.625 -181.100 ;
        RECT 3.040 -181.325 4.625 -181.105 ;
        RECT 3.945 -181.330 4.625 -181.325 ;
        RECT 13.610 -182.160 13.750 -178.435 ;
        RECT 14.025 -181.790 14.165 -177.750 ;
        RECT 16.260 -177.805 16.955 -177.740 ;
        RECT 22.050 -177.750 30.690 -177.610 ;
        RECT 22.050 -177.790 22.745 -177.750 ;
        RECT 16.260 -177.945 18.030 -177.805 ;
        RECT 25.125 -177.820 25.820 -177.750 ;
        RECT 16.260 -178.010 16.955 -177.945 ;
        RECT 17.890 -178.670 18.030 -177.945 ;
        RECT 20.005 -177.935 20.700 -177.890 ;
        RECT 24.190 -177.935 24.870 -177.890 ;
        RECT 20.005 -178.075 24.870 -177.935 ;
        RECT 20.005 -178.160 20.700 -178.075 ;
        RECT 24.190 -178.120 24.870 -178.075 ;
        RECT 22.660 -178.670 23.315 -178.610 ;
        RECT 17.890 -178.810 23.315 -178.670 ;
        RECT 22.660 -178.840 23.315 -178.810 ;
        RECT 15.120 -179.855 15.350 -179.175 ;
        RECT 15.125 -181.415 15.345 -179.855 ;
        RECT 16.235 -180.000 16.465 -179.000 ;
        RECT 16.725 -180.000 16.955 -179.000 ;
        RECT 18.305 -180.000 18.535 -179.000 ;
        RECT 18.795 -180.000 19.025 -179.000 ;
        RECT 20.115 -180.000 20.345 -179.000 ;
        RECT 20.605 -180.000 20.835 -179.000 ;
        RECT 21.585 -180.000 21.815 -179.000 ;
        RECT 22.075 -180.000 22.305 -179.000 ;
        RECT 23.135 -180.000 23.365 -179.000 ;
        RECT 23.625 -180.000 23.855 -179.000 ;
        RECT 24.680 -180.000 24.910 -179.000 ;
        RECT 25.170 -180.000 25.400 -179.000 ;
        RECT 29.645 -179.855 29.875 -179.175 ;
        RECT 29.650 -181.335 29.870 -179.855 ;
        RECT 30.550 -181.125 30.690 -177.750 ;
        RECT 31.260 -177.805 31.955 -177.740 ;
        RECT 37.050 -177.750 51.475 -177.610 ;
        RECT 37.050 -177.790 37.745 -177.750 ;
        RECT 31.260 -177.945 33.030 -177.805 ;
        RECT 40.125 -177.820 40.820 -177.750 ;
        RECT 31.260 -178.010 31.955 -177.945 ;
        RECT 32.890 -178.670 33.030 -177.945 ;
        RECT 35.005 -177.935 35.700 -177.890 ;
        RECT 39.190 -177.935 39.870 -177.890 ;
        RECT 35.005 -178.075 39.870 -177.935 ;
        RECT 35.005 -178.160 35.700 -178.075 ;
        RECT 39.190 -178.120 39.870 -178.075 ;
        RECT 37.660 -178.670 38.315 -178.610 ;
        RECT 32.890 -178.810 38.315 -178.670 ;
        RECT 37.660 -178.840 38.315 -178.810 ;
        RECT 31.235 -180.000 31.465 -179.000 ;
        RECT 31.725 -180.000 31.955 -179.000 ;
        RECT 33.305 -180.000 33.535 -179.000 ;
        RECT 33.795 -180.000 34.025 -179.000 ;
        RECT 35.115 -180.000 35.345 -179.000 ;
        RECT 35.605 -180.000 35.835 -179.000 ;
        RECT 36.585 -180.000 36.815 -179.000 ;
        RECT 37.075 -180.000 37.305 -179.000 ;
        RECT 38.135 -180.000 38.365 -179.000 ;
        RECT 38.625 -180.000 38.855 -179.000 ;
        RECT 39.680 -180.000 39.910 -179.000 ;
        RECT 40.170 -180.000 40.400 -179.000 ;
        RECT 44.690 -181.125 50.650 -180.540 ;
        RECT 30.550 -181.265 50.695 -181.125 ;
        RECT 14.860 -181.645 15.540 -181.415 ;
        RECT 29.385 -181.565 30.065 -181.335 ;
        RECT 14.025 -181.980 49.930 -181.790 ;
        RECT 13.610 -182.300 49.555 -182.160 ;
        RECT 1.650 -182.615 49.170 -182.475 ;
        RECT 1.280 -182.900 48.745 -182.760 ;
        RECT -10.710 -183.295 48.375 -183.040 ;
        RECT -11.140 -183.635 47.950 -183.455 ;
        RECT -23.565 -184.045 47.595 -183.790 ;
        RECT -22.090 -184.640 -21.410 -184.630 ;
        RECT 13.155 -184.640 13.835 -184.620 ;
        RECT -22.090 -184.850 13.835 -184.640 ;
        RECT -22.090 -184.860 -21.410 -184.850 ;
        RECT -34.490 -185.050 -33.810 -185.040 ;
        RECT 12.635 -185.050 13.410 -185.040 ;
        RECT -34.490 -185.260 13.410 -185.050 ;
        RECT -34.490 -185.270 -33.810 -185.260 ;
        RECT 12.635 -185.270 13.410 -185.260 ;
        RECT -32.865 -188.130 -32.635 -187.130 ;
        RECT -31.885 -188.130 -31.655 -187.130 ;
        RECT -30.905 -188.130 -30.675 -187.130 ;
        RECT -28.675 -187.705 -28.445 -187.205 ;
        RECT -28.185 -187.705 -27.955 -187.205 ;
        RECT -27.695 -187.705 -27.465 -187.205 ;
        RECT -27.205 -187.705 -26.975 -187.205 ;
        RECT -26.715 -187.705 -26.485 -187.205 ;
        RECT -26.225 -187.705 -25.995 -187.205 ;
        RECT -25.735 -187.705 -25.505 -187.205 ;
        RECT -25.245 -187.705 -25.015 -187.205 ;
        RECT -24.150 -188.130 -23.920 -187.130 ;
        RECT -23.170 -188.130 -22.940 -187.130 ;
        RECT -22.190 -188.130 -21.960 -187.130 ;
        RECT -25.875 -188.395 -25.030 -188.345 ;
        RECT -21.170 -188.395 -20.885 -187.220 ;
        RECT -19.365 -188.130 -19.135 -187.130 ;
        RECT -18.385 -188.130 -18.155 -187.130 ;
        RECT -17.405 -188.130 -17.175 -187.130 ;
        RECT -15.175 -187.705 -14.945 -187.205 ;
        RECT -14.685 -187.705 -14.455 -187.205 ;
        RECT -14.195 -187.705 -13.965 -187.205 ;
        RECT -13.705 -187.705 -13.475 -187.205 ;
        RECT -13.215 -187.705 -12.985 -187.205 ;
        RECT -12.725 -187.705 -12.495 -187.205 ;
        RECT -12.235 -187.705 -12.005 -187.205 ;
        RECT -11.745 -187.705 -11.515 -187.205 ;
        RECT -10.650 -188.130 -10.420 -187.130 ;
        RECT -9.670 -188.130 -9.440 -187.130 ;
        RECT -8.690 -188.130 -8.460 -187.130 ;
        RECT -25.875 -188.680 -20.885 -188.395 ;
        RECT -12.375 -188.395 -11.530 -188.345 ;
        RECT -7.670 -188.395 -7.385 -187.220 ;
        RECT -6.240 -188.130 -6.010 -187.130 ;
        RECT -5.260 -188.130 -5.030 -187.130 ;
        RECT -4.280 -188.130 -4.050 -187.130 ;
        RECT -1.590 -188.215 -1.360 -187.215 ;
        RECT 2.100 -188.215 2.330 -187.215 ;
        RECT 3.080 -188.215 3.310 -187.215 ;
        RECT 4.060 -188.215 4.290 -187.215 ;
        RECT 5.190 -188.020 5.420 -188.010 ;
        RECT -25.875 -188.715 -25.030 -188.680 ;
        RECT -32.865 -189.530 -32.635 -189.030 ;
        RECT -32.375 -189.530 -32.145 -189.030 ;
        RECT -31.885 -189.530 -31.655 -189.030 ;
        RECT -31.395 -189.530 -31.165 -189.030 ;
        RECT -30.905 -189.530 -30.675 -189.030 ;
        RECT -30.415 -189.530 -30.185 -189.030 ;
        RECT -28.675 -189.505 -28.445 -189.280 ;
        RECT -31.740 -190.115 -31.080 -189.815 ;
        RECT -33.435 -190.595 -33.135 -190.465 ;
        RECT -35.210 -190.910 -33.135 -190.595 ;
        RECT -35.125 -190.915 -33.135 -190.910 ;
        RECT -33.435 -191.150 -33.135 -190.915 ;
        RECT -31.620 -191.205 -31.145 -190.115 ;
        RECT -28.685 -190.275 -28.445 -189.505 ;
        RECT -28.185 -189.780 -27.955 -189.280 ;
        RECT -27.695 -189.685 -27.465 -189.280 ;
        RECT -27.725 -190.275 -27.420 -189.685 ;
        RECT -27.205 -189.780 -26.975 -189.280 ;
        RECT -26.715 -189.675 -26.485 -189.280 ;
        RECT -26.745 -190.275 -26.440 -189.675 ;
        RECT -26.225 -189.780 -25.995 -189.280 ;
        RECT -25.735 -189.685 -25.505 -189.280 ;
        RECT -25.790 -190.275 -25.485 -189.685 ;
        RECT -25.245 -189.780 -25.015 -189.280 ;
        RECT -24.150 -189.530 -23.920 -189.030 ;
        RECT -23.660 -189.530 -23.430 -189.030 ;
        RECT -23.170 -189.530 -22.940 -189.030 ;
        RECT -22.680 -189.530 -22.450 -189.030 ;
        RECT -22.190 -189.530 -21.960 -189.030 ;
        RECT -21.700 -189.530 -21.470 -189.030 ;
        RECT -28.685 -190.515 -21.030 -190.275 ;
        RECT -31.695 -191.505 -31.010 -191.205 ;
        RECT -32.865 -192.820 -32.635 -192.320 ;
        RECT -32.375 -192.820 -32.145 -192.320 ;
        RECT -31.885 -192.820 -31.655 -192.320 ;
        RECT -31.395 -192.820 -31.165 -192.320 ;
        RECT -30.905 -192.820 -30.675 -192.320 ;
        RECT -30.415 -192.820 -30.185 -192.320 ;
        RECT -28.680 -192.820 -28.450 -192.320 ;
        RECT -28.190 -192.820 -27.960 -192.320 ;
        RECT -27.700 -192.820 -27.470 -192.320 ;
        RECT -27.210 -192.820 -26.980 -192.320 ;
        RECT -26.720 -192.820 -26.490 -192.320 ;
        RECT -26.230 -192.820 -26.000 -192.320 ;
        RECT -25.135 -192.570 -24.905 -192.070 ;
        RECT -24.645 -192.570 -24.415 -192.070 ;
        RECT -24.155 -192.570 -23.925 -192.070 ;
        RECT -23.665 -192.570 -23.435 -192.070 ;
        RECT -23.175 -192.570 -22.945 -192.070 ;
        RECT -22.685 -192.570 -22.455 -192.070 ;
        RECT -22.195 -192.570 -21.965 -192.070 ;
        RECT -21.705 -192.570 -21.475 -192.070 ;
        RECT -21.235 -192.940 -21.030 -190.515 ;
        RECT -20.640 -190.760 -20.340 -188.520 ;
        RECT -20.065 -189.080 -19.765 -188.645 ;
        RECT -12.375 -188.680 -7.385 -188.395 ;
        RECT -12.375 -188.715 -11.530 -188.680 ;
        RECT -20.065 -189.305 -19.760 -189.080 ;
        RECT -20.885 -191.060 -20.200 -190.760 ;
        RECT -25.120 -193.170 -24.275 -193.135 ;
        RECT -29.265 -193.455 -24.275 -193.170 ;
        RECT -21.710 -193.240 -21.025 -192.940 ;
        RECT -20.060 -193.045 -19.760 -189.305 ;
        RECT -19.365 -189.530 -19.135 -189.030 ;
        RECT -18.875 -189.530 -18.645 -189.030 ;
        RECT -18.385 -189.530 -18.155 -189.030 ;
        RECT -17.895 -189.530 -17.665 -189.030 ;
        RECT -17.405 -189.530 -17.175 -189.030 ;
        RECT -16.915 -189.530 -16.685 -189.030 ;
        RECT -15.175 -189.780 -14.930 -189.280 ;
        RECT -14.685 -189.780 -14.455 -189.280 ;
        RECT -14.195 -189.780 -13.965 -189.280 ;
        RECT -13.705 -189.780 -13.475 -189.280 ;
        RECT -13.215 -189.780 -12.985 -189.280 ;
        RECT -12.725 -189.780 -12.495 -189.280 ;
        RECT -12.235 -189.780 -12.005 -189.280 ;
        RECT -11.745 -189.780 -11.515 -189.280 ;
        RECT -10.650 -189.530 -10.420 -189.030 ;
        RECT -10.160 -189.530 -9.930 -189.030 ;
        RECT -9.670 -189.530 -9.440 -189.030 ;
        RECT -9.180 -189.530 -8.950 -189.030 ;
        RECT -8.690 -189.530 -8.460 -189.030 ;
        RECT -8.200 -189.530 -7.970 -189.030 ;
        RECT -18.745 -190.135 -18.060 -189.835 ;
        RECT -18.655 -191.175 -18.180 -190.135 ;
        RECT -15.160 -190.265 -14.930 -189.780 ;
        RECT -14.185 -190.265 -13.975 -189.780 ;
        RECT -13.210 -190.265 -13.000 -189.780 ;
        RECT -12.230 -190.265 -12.020 -189.780 ;
        RECT -15.160 -190.495 -11.360 -190.265 ;
        RECT -16.155 -191.055 -15.495 -190.755 ;
        RECT -18.710 -191.475 -18.025 -191.175 ;
        RECT -19.365 -192.820 -19.135 -192.320 ;
        RECT -18.875 -192.820 -18.645 -192.320 ;
        RECT -18.385 -192.820 -18.155 -192.320 ;
        RECT -17.895 -192.820 -17.665 -192.320 ;
        RECT -17.405 -192.820 -17.175 -192.320 ;
        RECT -16.915 -192.820 -16.685 -192.320 ;
        RECT -16.010 -192.875 -15.710 -191.055 ;
        RECT -11.590 -191.325 -11.360 -190.495 ;
        RECT -7.670 -190.865 -7.385 -188.680 ;
        RECT -6.980 -189.185 -6.680 -188.525 ;
        RECT 5.150 -188.690 5.420 -188.020 ;
        RECT 7.075 -188.060 7.305 -187.280 ;
        RECT 8.055 -188.050 8.285 -187.280 ;
        RECT 7.565 -188.060 8.775 -188.050 ;
        RECT 9.035 -188.060 9.265 -187.280 ;
        RECT 6.950 -188.290 9.265 -188.060 ;
        RECT -6.970 -190.325 -6.680 -189.185 ;
        RECT -6.240 -189.530 -6.010 -189.030 ;
        RECT -5.750 -189.530 -5.520 -189.030 ;
        RECT -5.260 -189.530 -5.030 -189.030 ;
        RECT -4.770 -189.530 -4.540 -189.030 ;
        RECT -4.280 -189.530 -4.050 -189.030 ;
        RECT -3.790 -189.530 -3.560 -189.030 ;
        RECT -2.315 -189.510 -1.610 -189.245 ;
        RECT -4.960 -190.130 -4.275 -189.830 ;
        RECT -6.970 -190.615 -5.775 -190.325 ;
        RECT -6.065 -190.760 -5.775 -190.615 ;
        RECT -7.670 -191.150 -6.340 -190.865 ;
        RECT -6.085 -191.060 -5.425 -190.760 ;
        RECT -11.590 -191.330 -7.535 -191.325 ;
        RECT -11.590 -191.555 -7.495 -191.330 ;
        RECT -15.180 -192.820 -14.950 -192.320 ;
        RECT -14.690 -192.820 -14.460 -192.320 ;
        RECT -14.200 -192.820 -13.970 -192.320 ;
        RECT -13.710 -192.820 -13.480 -192.320 ;
        RECT -13.220 -192.820 -12.990 -192.320 ;
        RECT -12.730 -192.820 -12.500 -192.320 ;
        RECT -11.635 -192.570 -11.405 -192.070 ;
        RECT -11.145 -192.570 -10.915 -192.070 ;
        RECT -10.655 -192.570 -10.425 -192.070 ;
        RECT -10.165 -192.570 -9.935 -192.070 ;
        RECT -9.675 -192.570 -9.445 -192.070 ;
        RECT -9.185 -192.570 -8.955 -192.070 ;
        RECT -8.695 -192.570 -8.465 -192.070 ;
        RECT -8.205 -192.570 -7.975 -192.070 ;
        RECT -7.725 -192.930 -7.495 -191.555 ;
        RECT -6.625 -191.755 -6.340 -191.150 ;
        RECT -4.785 -191.175 -4.310 -190.130 ;
        RECT -4.870 -191.475 -4.210 -191.175 ;
        RECT -2.315 -191.755 -2.030 -189.510 ;
        RECT -1.590 -191.755 -1.360 -190.755 ;
        RECT -1.100 -191.755 -0.870 -190.755 ;
        RECT 0.475 -191.755 0.705 -190.255 ;
        RECT 0.965 -191.755 1.195 -190.255 ;
        RECT 1.455 -191.755 1.685 -190.255 ;
        RECT 2.020 -191.755 2.250 -190.255 ;
        RECT 2.510 -191.755 2.740 -190.255 ;
        RECT 3.000 -191.755 3.230 -190.255 ;
        RECT 3.570 -191.750 3.800 -190.250 ;
        RECT 4.060 -191.750 4.290 -190.250 ;
        RECT 4.550 -191.750 4.780 -190.250 ;
        RECT -6.625 -192.040 -2.030 -191.755 ;
        RECT -21.235 -193.245 -21.030 -193.240 ;
        RECT -20.060 -193.345 -19.345 -193.045 ;
        RECT -11.620 -193.170 -10.775 -193.135 ;
        RECT -20.060 -193.375 -19.760 -193.345 ;
        RECT -32.375 -194.720 -32.145 -193.720 ;
        RECT -31.395 -194.720 -31.165 -193.720 ;
        RECT -30.415 -194.720 -30.185 -193.720 ;
        RECT -29.265 -194.630 -28.980 -193.455 ;
        RECT -25.120 -193.505 -24.275 -193.455 ;
        RECT -15.765 -193.455 -10.775 -193.170 ;
        RECT -8.265 -193.230 -7.495 -192.930 ;
        RECT 5.150 -192.715 5.380 -188.690 ;
        RECT 5.595 -189.110 6.275 -188.880 ;
        RECT 7.565 -188.935 7.795 -188.290 ;
        RECT 8.055 -188.935 8.285 -188.435 ;
        RECT 8.545 -188.935 8.775 -188.290 ;
        RECT 9.035 -188.935 9.265 -188.435 ;
        RECT 5.915 -192.155 6.145 -189.110 ;
        RECT 10.610 -191.650 10.840 -189.970 ;
        RECT 11.100 -191.470 11.330 -187.285 ;
        RECT 12.080 -188.785 12.310 -187.285 ;
        RECT 15.100 -188.070 15.330 -187.290 ;
        RECT 16.080 -188.060 16.310 -187.290 ;
        RECT 15.590 -188.070 16.800 -188.060 ;
        RECT 17.060 -188.070 17.290 -187.290 ;
        RECT 14.975 -188.300 17.290 -188.070 ;
        RECT 15.590 -188.945 15.820 -188.300 ;
        RECT 16.080 -188.945 16.310 -188.445 ;
        RECT 16.570 -188.945 16.800 -188.300 ;
        RECT 17.060 -188.945 17.290 -188.445 ;
        RECT 11.590 -191.650 11.820 -189.970 ;
        RECT 12.080 -191.470 12.310 -189.970 ;
        RECT 12.570 -191.465 12.800 -189.970 ;
        RECT 12.570 -191.650 12.805 -191.465 ;
        RECT 10.610 -191.885 12.805 -191.650 ;
        RECT 18.635 -191.660 18.865 -189.980 ;
        RECT 19.125 -191.480 19.355 -187.295 ;
        RECT 20.105 -188.795 20.335 -187.295 ;
        RECT 23.220 -188.170 23.450 -187.170 ;
        RECT 26.910 -188.170 27.140 -187.170 ;
        RECT 27.890 -188.170 28.120 -187.170 ;
        RECT 28.870 -188.170 29.100 -187.170 ;
        RECT 31.285 -188.225 31.515 -187.225 ;
        RECT 31.775 -188.380 32.005 -187.225 ;
        RECT 32.265 -188.225 32.495 -187.225 ;
        RECT 32.865 -188.225 33.095 -187.225 ;
        RECT 33.355 -188.225 33.585 -187.225 ;
        RECT 33.845 -188.225 34.075 -187.225 ;
        RECT 35.655 -188.225 35.885 -187.225 ;
        RECT 36.635 -188.225 36.865 -187.225 ;
        RECT 38.185 -188.225 38.415 -187.225 ;
        RECT 39.730 -188.225 39.960 -187.225 ;
        RECT 29.245 -188.610 32.005 -188.380 ;
        RECT 29.265 -188.655 29.945 -188.610 ;
        RECT 37.100 -188.865 37.795 -188.775 ;
        RECT 40.175 -188.830 40.870 -188.805 ;
        RECT 44.830 -188.830 45.920 -188.535 ;
        RECT 40.175 -188.865 45.920 -188.830 ;
        RECT 37.100 -188.970 45.920 -188.865 ;
        RECT 31.310 -189.060 32.005 -188.995 ;
        RECT 37.100 -189.005 41.375 -188.970 ;
        RECT 44.830 -188.980 45.920 -188.970 ;
        RECT 37.100 -189.045 37.795 -189.005 ;
        RECT 31.310 -189.200 33.080 -189.060 ;
        RECT 40.175 -189.075 40.870 -189.005 ;
        RECT 31.310 -189.265 32.005 -189.200 ;
        RECT 32.940 -189.925 33.080 -189.200 ;
        RECT 35.055 -189.190 35.750 -189.145 ;
        RECT 39.240 -189.190 39.920 -189.145 ;
        RECT 35.055 -189.330 39.920 -189.190 ;
        RECT 35.055 -189.415 35.750 -189.330 ;
        RECT 39.240 -189.375 39.920 -189.330 ;
        RECT 37.710 -189.925 38.365 -189.865 ;
        RECT 19.615 -191.660 19.845 -189.980 ;
        RECT 20.105 -191.480 20.335 -189.980 ;
        RECT 20.595 -191.475 20.825 -189.980 ;
        RECT 32.940 -190.065 38.365 -189.925 ;
        RECT 37.710 -190.095 38.365 -190.065 ;
        RECT 20.595 -191.660 20.830 -191.475 ;
        RECT 18.635 -191.895 20.830 -191.660 ;
        RECT 23.220 -191.710 23.450 -190.710 ;
        RECT 23.710 -191.710 23.940 -190.710 ;
        RECT 25.285 -191.710 25.515 -190.210 ;
        RECT 25.775 -191.710 26.005 -190.210 ;
        RECT 26.265 -191.710 26.495 -190.210 ;
        RECT 26.830 -191.710 27.060 -190.210 ;
        RECT 27.320 -191.710 27.550 -190.210 ;
        RECT 27.810 -191.710 28.040 -190.210 ;
        RECT 28.380 -191.705 28.610 -190.205 ;
        RECT 28.870 -191.705 29.100 -190.205 ;
        RECT 29.360 -191.705 29.590 -190.205 ;
        RECT 31.285 -191.255 31.515 -190.255 ;
        RECT 31.775 -191.255 32.005 -190.255 ;
        RECT 33.355 -191.255 33.585 -190.255 ;
        RECT 33.845 -191.255 34.075 -190.255 ;
        RECT 35.165 -191.255 35.395 -190.255 ;
        RECT 35.655 -191.255 35.885 -190.255 ;
        RECT 36.635 -191.255 36.865 -190.255 ;
        RECT 37.125 -191.255 37.355 -190.255 ;
        RECT 38.185 -191.255 38.415 -190.255 ;
        RECT 38.675 -191.255 38.905 -190.255 ;
        RECT 39.730 -191.255 39.960 -190.255 ;
        RECT 40.220 -191.255 40.450 -190.255 ;
        RECT 5.915 -192.385 14.660 -192.155 ;
        RECT 5.150 -192.945 22.500 -192.715 ;
        RECT -28.190 -194.720 -27.960 -193.720 ;
        RECT -27.210 -194.720 -26.980 -193.720 ;
        RECT -26.230 -194.720 -26.000 -193.720 ;
        RECT -25.135 -194.645 -24.905 -194.145 ;
        RECT -24.645 -194.645 -24.415 -194.145 ;
        RECT -24.155 -194.645 -23.925 -194.145 ;
        RECT -23.665 -194.645 -23.435 -194.145 ;
        RECT -23.175 -194.645 -22.945 -194.145 ;
        RECT -22.685 -194.645 -22.455 -194.145 ;
        RECT -22.195 -194.645 -21.965 -194.145 ;
        RECT -21.705 -194.645 -21.475 -194.145 ;
        RECT -18.875 -194.720 -18.645 -193.720 ;
        RECT -17.895 -194.720 -17.665 -193.720 ;
        RECT -16.915 -194.720 -16.685 -193.720 ;
        RECT -15.765 -194.630 -15.480 -193.455 ;
        RECT -11.620 -193.505 -10.775 -193.455 ;
        RECT -14.690 -194.720 -14.460 -193.720 ;
        RECT -13.710 -194.720 -13.480 -193.720 ;
        RECT -12.730 -194.720 -12.500 -193.720 ;
        RECT -11.635 -194.645 -11.405 -194.145 ;
        RECT -11.145 -194.645 -10.915 -194.145 ;
        RECT -10.655 -194.645 -10.425 -194.145 ;
        RECT -10.165 -194.645 -9.935 -194.145 ;
        RECT -9.675 -194.645 -9.445 -194.145 ;
        RECT -9.185 -194.645 -8.955 -194.145 ;
        RECT -8.695 -194.645 -8.465 -194.145 ;
        RECT -8.205 -194.645 -7.975 -194.145 ;
        RECT -32.375 -201.910 -32.145 -200.910 ;
        RECT -31.395 -201.910 -31.165 -200.910 ;
        RECT -30.415 -201.910 -30.185 -200.910 ;
        RECT -29.265 -202.175 -28.980 -201.000 ;
        RECT -28.190 -201.910 -27.960 -200.910 ;
        RECT -27.210 -201.910 -26.980 -200.910 ;
        RECT -26.230 -201.910 -26.000 -200.910 ;
        RECT -25.135 -201.485 -24.905 -200.985 ;
        RECT -24.645 -201.485 -24.415 -200.985 ;
        RECT -24.155 -201.485 -23.925 -200.985 ;
        RECT -23.665 -201.485 -23.435 -200.985 ;
        RECT -23.175 -201.485 -22.945 -200.985 ;
        RECT -22.685 -201.485 -22.455 -200.985 ;
        RECT -22.195 -201.485 -21.965 -200.985 ;
        RECT -21.705 -201.485 -21.475 -200.985 ;
        RECT -18.875 -201.910 -18.645 -200.910 ;
        RECT -17.895 -201.910 -17.665 -200.910 ;
        RECT -16.915 -201.910 -16.685 -200.910 ;
        RECT -25.120 -202.175 -24.275 -202.125 ;
        RECT -29.265 -202.460 -24.275 -202.175 ;
        RECT -15.765 -202.175 -15.480 -201.000 ;
        RECT -14.690 -201.910 -14.460 -200.910 ;
        RECT -13.710 -201.910 -13.480 -200.910 ;
        RECT -12.730 -201.910 -12.500 -200.910 ;
        RECT -11.635 -201.485 -11.405 -200.985 ;
        RECT -11.145 -201.485 -10.915 -200.985 ;
        RECT -10.655 -201.485 -10.425 -200.985 ;
        RECT -10.165 -201.485 -9.935 -200.985 ;
        RECT -9.675 -201.485 -9.445 -200.985 ;
        RECT -9.185 -201.485 -8.955 -200.985 ;
        RECT -8.695 -201.485 -8.465 -200.985 ;
        RECT -8.205 -201.485 -7.975 -200.985 ;
        RECT -11.620 -202.175 -10.775 -202.125 ;
        RECT -20.060 -202.285 -19.760 -202.255 ;
        RECT -21.235 -202.390 -21.030 -202.385 ;
        RECT -25.120 -202.495 -24.275 -202.460 ;
        RECT -32.865 -203.310 -32.635 -202.810 ;
        RECT -32.375 -203.310 -32.145 -202.810 ;
        RECT -31.885 -203.310 -31.655 -202.810 ;
        RECT -31.395 -203.310 -31.165 -202.810 ;
        RECT -30.905 -203.310 -30.675 -202.810 ;
        RECT -30.415 -203.310 -30.185 -202.810 ;
        RECT -35.165 -204.715 -34.290 -203.620 ;
        RECT -31.695 -204.425 -31.010 -204.125 ;
        RECT -33.435 -204.715 -33.135 -204.480 ;
        RECT -35.165 -205.035 -33.135 -204.715 ;
        RECT -35.165 -205.190 -34.290 -205.035 ;
        RECT -33.435 -205.165 -33.135 -205.035 ;
        RECT -31.620 -205.365 -31.145 -204.425 ;
        RECT -29.570 -205.015 -29.270 -202.680 ;
        RECT -21.710 -202.690 -21.025 -202.390 ;
        RECT -20.060 -202.585 -19.345 -202.285 ;
        RECT -15.765 -202.460 -10.775 -202.175 ;
        RECT -11.620 -202.495 -10.775 -202.460 ;
        RECT -28.680 -203.310 -28.450 -202.810 ;
        RECT -28.190 -203.310 -27.960 -202.810 ;
        RECT -27.700 -203.310 -27.470 -202.810 ;
        RECT -27.210 -203.310 -26.980 -202.810 ;
        RECT -26.720 -203.310 -26.490 -202.810 ;
        RECT -26.230 -203.310 -26.000 -202.810 ;
        RECT -25.135 -203.560 -24.905 -203.060 ;
        RECT -24.645 -203.560 -24.415 -203.060 ;
        RECT -24.155 -203.560 -23.925 -203.060 ;
        RECT -23.665 -203.560 -23.435 -203.060 ;
        RECT -23.175 -203.560 -22.945 -203.060 ;
        RECT -22.685 -203.560 -22.455 -203.060 ;
        RECT -22.195 -203.560 -21.965 -203.060 ;
        RECT -21.705 -203.560 -21.475 -203.060 ;
        RECT -29.750 -205.315 -29.090 -205.015 ;
        RECT -21.235 -205.115 -21.030 -202.690 ;
        RECT -34.055 -205.515 -31.145 -205.365 ;
        RECT -28.685 -205.355 -21.030 -205.115 ;
        RECT -34.055 -205.815 -31.080 -205.515 ;
        RECT -34.055 -205.840 -31.145 -205.815 ;
        RECT -34.055 -206.235 -33.580 -205.840 ;
        RECT -35.130 -206.710 -33.580 -206.235 ;
        RECT -32.865 -206.600 -32.635 -206.100 ;
        RECT -32.375 -206.600 -32.145 -206.100 ;
        RECT -31.885 -206.600 -31.655 -206.100 ;
        RECT -31.395 -206.600 -31.165 -206.100 ;
        RECT -30.905 -206.600 -30.675 -206.100 ;
        RECT -30.415 -206.600 -30.185 -206.100 ;
        RECT -28.685 -206.125 -28.445 -205.355 ;
        RECT -28.675 -206.350 -28.445 -206.125 ;
        RECT -28.185 -206.350 -27.955 -205.850 ;
        RECT -27.725 -205.945 -27.420 -205.355 ;
        RECT -27.695 -206.350 -27.465 -205.945 ;
        RECT -27.205 -206.350 -26.975 -205.850 ;
        RECT -26.745 -205.955 -26.440 -205.355 ;
        RECT -26.715 -206.350 -26.485 -205.955 ;
        RECT -26.225 -206.350 -25.995 -205.850 ;
        RECT -25.790 -205.945 -25.485 -205.355 ;
        RECT -25.735 -206.350 -25.505 -205.945 ;
        RECT -25.245 -206.350 -25.015 -205.850 ;
        RECT -24.150 -206.600 -23.920 -206.100 ;
        RECT -23.660 -206.600 -23.430 -206.100 ;
        RECT -23.170 -206.600 -22.940 -206.100 ;
        RECT -22.680 -206.600 -22.450 -206.100 ;
        RECT -22.190 -206.600 -21.960 -206.100 ;
        RECT -21.700 -206.600 -21.470 -206.100 ;
        RECT -20.060 -206.325 -19.760 -202.585 ;
        RECT -8.265 -202.700 -7.495 -202.400 ;
        RECT -19.365 -203.310 -19.135 -202.810 ;
        RECT -18.875 -203.310 -18.645 -202.810 ;
        RECT -18.385 -203.310 -18.155 -202.810 ;
        RECT -17.895 -203.310 -17.665 -202.810 ;
        RECT -17.405 -203.310 -17.175 -202.810 ;
        RECT -16.915 -203.310 -16.685 -202.810 ;
        RECT -15.180 -203.310 -14.950 -202.810 ;
        RECT -14.690 -203.310 -14.460 -202.810 ;
        RECT -14.200 -203.310 -13.970 -202.810 ;
        RECT -13.710 -203.310 -13.480 -202.810 ;
        RECT -13.220 -203.310 -12.990 -202.810 ;
        RECT -12.730 -203.310 -12.500 -202.810 ;
        RECT -11.635 -203.560 -11.405 -203.060 ;
        RECT -11.145 -203.560 -10.915 -203.060 ;
        RECT -10.655 -203.560 -10.425 -203.060 ;
        RECT -10.165 -203.560 -9.935 -203.060 ;
        RECT -9.675 -203.560 -9.445 -203.060 ;
        RECT -9.185 -203.560 -8.955 -203.060 ;
        RECT -8.695 -203.560 -8.465 -203.060 ;
        RECT -8.205 -203.560 -7.975 -203.060 ;
        RECT -7.725 -204.075 -7.495 -202.700 ;
        RECT 5.150 -202.915 22.500 -202.685 ;
        RECT -18.710 -204.455 -18.025 -204.155 ;
        RECT -11.590 -204.300 -7.495 -204.075 ;
        RECT -6.625 -203.875 -2.030 -203.590 ;
        RECT -11.590 -204.305 -7.535 -204.300 ;
        RECT -18.655 -205.495 -18.180 -204.455 ;
        RECT -11.590 -205.135 -11.360 -204.305 ;
        RECT -6.625 -204.480 -6.340 -203.875 ;
        RECT -5.520 -204.455 -4.860 -204.155 ;
        RECT -15.160 -205.365 -11.360 -205.135 ;
        RECT -7.670 -204.765 -6.340 -204.480 ;
        RECT -18.745 -205.795 -18.060 -205.495 ;
        RECT -15.160 -205.850 -14.930 -205.365 ;
        RECT -14.185 -205.850 -13.975 -205.365 ;
        RECT -13.210 -205.850 -13.000 -205.365 ;
        RECT -12.230 -205.850 -12.020 -205.365 ;
        RECT -20.065 -206.550 -19.760 -206.325 ;
        RECT -25.875 -206.950 -25.030 -206.915 ;
        RECT -25.875 -207.235 -20.885 -206.950 ;
        RECT -20.065 -206.985 -19.765 -206.550 ;
        RECT -19.365 -206.600 -19.135 -206.100 ;
        RECT -18.875 -206.600 -18.645 -206.100 ;
        RECT -18.385 -206.600 -18.155 -206.100 ;
        RECT -17.895 -206.600 -17.665 -206.100 ;
        RECT -17.405 -206.600 -17.175 -206.100 ;
        RECT -16.915 -206.600 -16.685 -206.100 ;
        RECT -15.175 -206.350 -14.930 -205.850 ;
        RECT -14.685 -206.350 -14.455 -205.850 ;
        RECT -14.195 -206.350 -13.965 -205.850 ;
        RECT -13.705 -206.350 -13.475 -205.850 ;
        RECT -13.215 -206.350 -12.985 -205.850 ;
        RECT -12.725 -206.350 -12.495 -205.850 ;
        RECT -12.235 -206.350 -12.005 -205.850 ;
        RECT -11.745 -206.350 -11.515 -205.850 ;
        RECT -10.650 -206.600 -10.420 -206.100 ;
        RECT -10.160 -206.600 -9.930 -206.100 ;
        RECT -9.670 -206.600 -9.440 -206.100 ;
        RECT -9.180 -206.600 -8.950 -206.100 ;
        RECT -8.690 -206.600 -8.460 -206.100 ;
        RECT -8.200 -206.600 -7.970 -206.100 ;
        RECT -12.375 -206.950 -11.530 -206.915 ;
        RECT -7.670 -206.950 -7.385 -204.765 ;
        RECT -7.135 -205.305 -6.475 -205.005 ;
        RECT -6.970 -206.445 -6.680 -205.305 ;
        RECT -5.435 -205.500 -4.960 -204.455 ;
        RECT -5.610 -205.800 -4.925 -205.500 ;
        RECT -25.875 -207.285 -25.030 -207.235 ;
        RECT -32.865 -208.500 -32.635 -207.500 ;
        RECT -31.885 -208.500 -31.655 -207.500 ;
        RECT -30.905 -208.500 -30.675 -207.500 ;
        RECT -28.675 -208.425 -28.445 -207.925 ;
        RECT -28.185 -208.425 -27.955 -207.925 ;
        RECT -27.695 -208.425 -27.465 -207.925 ;
        RECT -27.205 -208.425 -26.975 -207.925 ;
        RECT -26.715 -208.425 -26.485 -207.925 ;
        RECT -26.225 -208.425 -25.995 -207.925 ;
        RECT -25.735 -208.425 -25.505 -207.925 ;
        RECT -25.245 -208.425 -25.015 -207.925 ;
        RECT -24.150 -208.500 -23.920 -207.500 ;
        RECT -23.170 -208.500 -22.940 -207.500 ;
        RECT -22.190 -208.500 -21.960 -207.500 ;
        RECT -21.170 -208.410 -20.885 -207.235 ;
        RECT -12.375 -207.235 -7.385 -206.950 ;
        RECT -6.980 -207.105 -6.680 -206.445 ;
        RECT -6.240 -206.600 -6.010 -206.100 ;
        RECT -5.750 -206.600 -5.520 -206.100 ;
        RECT -5.260 -206.600 -5.030 -206.100 ;
        RECT -4.770 -206.600 -4.540 -206.100 ;
        RECT -4.280 -206.600 -4.050 -206.100 ;
        RECT -3.790 -206.600 -3.560 -206.100 ;
        RECT -2.315 -206.120 -2.030 -203.875 ;
        RECT -1.590 -204.875 -1.360 -203.875 ;
        RECT -1.100 -204.875 -0.870 -203.875 ;
        RECT 0.475 -205.375 0.705 -203.875 ;
        RECT 0.965 -205.375 1.195 -203.875 ;
        RECT 1.455 -205.375 1.685 -203.875 ;
        RECT 2.020 -205.375 2.250 -203.875 ;
        RECT 2.510 -205.375 2.740 -203.875 ;
        RECT 3.000 -205.375 3.230 -203.875 ;
        RECT 3.570 -205.380 3.800 -203.880 ;
        RECT 4.060 -205.380 4.290 -203.880 ;
        RECT 4.550 -205.380 4.780 -203.880 ;
        RECT -2.315 -206.385 -1.610 -206.120 ;
        RECT 5.150 -206.940 5.380 -202.915 ;
        RECT 5.915 -203.475 14.660 -203.245 ;
        RECT 5.915 -206.520 6.145 -203.475 ;
        RECT 10.610 -203.980 12.805 -203.745 ;
        RECT 10.610 -205.660 10.840 -203.980 ;
        RECT 5.595 -206.750 6.275 -206.520 ;
        RECT -12.375 -207.285 -11.530 -207.235 ;
        RECT -19.365 -208.500 -19.135 -207.500 ;
        RECT -18.385 -208.500 -18.155 -207.500 ;
        RECT -17.405 -208.500 -17.175 -207.500 ;
        RECT -15.175 -208.425 -14.945 -207.925 ;
        RECT -14.685 -208.425 -14.455 -207.925 ;
        RECT -14.195 -208.425 -13.965 -207.925 ;
        RECT -13.705 -208.425 -13.475 -207.925 ;
        RECT -13.215 -208.425 -12.985 -207.925 ;
        RECT -12.725 -208.425 -12.495 -207.925 ;
        RECT -12.235 -208.425 -12.005 -207.925 ;
        RECT -11.745 -208.425 -11.515 -207.925 ;
        RECT -10.650 -208.500 -10.420 -207.500 ;
        RECT -9.670 -208.500 -9.440 -207.500 ;
        RECT -8.690 -208.500 -8.460 -207.500 ;
        RECT -7.670 -208.410 -7.385 -207.235 ;
        RECT -6.240 -208.500 -6.010 -207.500 ;
        RECT -5.260 -208.500 -5.030 -207.500 ;
        RECT -4.280 -208.500 -4.050 -207.500 ;
        RECT -1.590 -208.415 -1.360 -207.415 ;
        RECT 2.100 -208.415 2.330 -207.415 ;
        RECT 3.080 -208.415 3.310 -207.415 ;
        RECT 4.060 -208.415 4.290 -207.415 ;
        RECT 5.150 -207.610 5.420 -206.940 ;
        RECT 7.565 -207.340 7.795 -206.695 ;
        RECT 8.055 -207.195 8.285 -206.695 ;
        RECT 8.545 -207.340 8.775 -206.695 ;
        RECT 9.035 -207.195 9.265 -206.695 ;
        RECT 6.950 -207.570 9.265 -207.340 ;
        RECT 5.190 -207.620 5.420 -207.610 ;
        RECT 7.075 -208.350 7.305 -207.570 ;
        RECT 7.565 -207.580 8.775 -207.570 ;
        RECT 8.055 -208.350 8.285 -207.580 ;
        RECT 9.035 -208.350 9.265 -207.570 ;
        RECT 11.100 -208.345 11.330 -204.160 ;
        RECT 11.590 -205.660 11.820 -203.980 ;
        RECT 12.080 -205.660 12.310 -204.160 ;
        RECT 12.570 -204.165 12.805 -203.980 ;
        RECT 18.635 -203.970 20.830 -203.735 ;
        RECT 12.570 -205.660 12.800 -204.165 ;
        RECT 18.635 -205.650 18.865 -203.970 ;
        RECT 12.080 -208.345 12.310 -206.845 ;
        RECT 15.590 -207.330 15.820 -206.685 ;
        RECT 16.080 -207.185 16.310 -206.685 ;
        RECT 16.570 -207.330 16.800 -206.685 ;
        RECT 17.060 -207.185 17.290 -206.685 ;
        RECT 14.975 -207.560 17.290 -207.330 ;
        RECT 15.100 -208.340 15.330 -207.560 ;
        RECT 15.590 -207.570 16.800 -207.560 ;
        RECT 16.080 -208.340 16.310 -207.570 ;
        RECT 17.060 -208.340 17.290 -207.560 ;
        RECT 19.125 -208.335 19.355 -204.150 ;
        RECT 19.615 -205.650 19.845 -203.970 ;
        RECT 20.105 -205.650 20.335 -204.150 ;
        RECT 20.595 -204.155 20.830 -203.970 ;
        RECT 20.595 -205.650 20.825 -204.155 ;
        RECT 23.220 -204.920 23.450 -203.920 ;
        RECT 23.710 -204.920 23.940 -203.920 ;
        RECT 25.285 -205.420 25.515 -203.920 ;
        RECT 25.775 -205.420 26.005 -203.920 ;
        RECT 26.265 -205.420 26.495 -203.920 ;
        RECT 26.830 -205.420 27.060 -203.920 ;
        RECT 27.320 -205.420 27.550 -203.920 ;
        RECT 27.810 -205.420 28.040 -203.920 ;
        RECT 28.380 -205.425 28.610 -203.925 ;
        RECT 28.870 -205.425 29.100 -203.925 ;
        RECT 29.360 -205.425 29.590 -203.925 ;
        RECT 31.285 -205.375 31.515 -204.375 ;
        RECT 31.775 -205.375 32.005 -204.375 ;
        RECT 33.355 -205.375 33.585 -204.375 ;
        RECT 33.845 -205.375 34.075 -204.375 ;
        RECT 35.165 -205.375 35.395 -204.375 ;
        RECT 35.655 -205.375 35.885 -204.375 ;
        RECT 36.635 -205.375 36.865 -204.375 ;
        RECT 37.125 -205.375 37.355 -204.375 ;
        RECT 38.185 -205.375 38.415 -204.375 ;
        RECT 38.675 -205.375 38.905 -204.375 ;
        RECT 39.730 -205.375 39.960 -204.375 ;
        RECT 40.220 -205.375 40.450 -204.375 ;
        RECT 37.710 -205.565 38.365 -205.535 ;
        RECT 32.940 -205.705 38.365 -205.565 ;
        RECT 31.310 -206.430 32.005 -206.365 ;
        RECT 32.940 -206.430 33.080 -205.705 ;
        RECT 37.710 -205.765 38.365 -205.705 ;
        RECT 31.310 -206.570 33.080 -206.430 ;
        RECT 35.055 -206.300 35.750 -206.215 ;
        RECT 39.240 -206.300 39.920 -206.255 ;
        RECT 35.055 -206.440 39.920 -206.300 ;
        RECT 35.055 -206.485 35.750 -206.440 ;
        RECT 39.240 -206.485 39.920 -206.440 ;
        RECT 31.310 -206.635 32.005 -206.570 ;
        RECT 37.100 -206.625 37.795 -206.585 ;
        RECT 40.175 -206.625 40.870 -206.555 ;
        RECT 37.100 -206.660 41.375 -206.625 ;
        RECT 45.665 -206.660 45.805 -188.980 ;
        RECT 47.340 -202.435 47.595 -184.045 ;
        RECT 47.325 -202.910 47.620 -202.435 ;
        RECT 37.100 -206.765 45.805 -206.660 ;
        RECT 20.105 -208.335 20.335 -206.835 ;
        RECT 37.100 -206.855 37.795 -206.765 ;
        RECT 40.175 -206.800 45.805 -206.765 ;
        RECT 40.175 -206.825 40.870 -206.800 ;
        RECT 29.265 -207.020 29.945 -206.975 ;
        RECT 29.245 -207.250 32.005 -207.020 ;
        RECT 23.220 -208.460 23.450 -207.460 ;
        RECT 26.910 -208.460 27.140 -207.460 ;
        RECT 27.890 -208.460 28.120 -207.460 ;
        RECT 28.870 -208.460 29.100 -207.460 ;
        RECT 31.285 -208.405 31.515 -207.405 ;
        RECT 31.775 -208.405 32.005 -207.250 ;
        RECT 32.265 -208.405 32.495 -207.405 ;
        RECT 32.865 -208.405 33.095 -207.405 ;
        RECT 33.355 -208.405 33.585 -207.405 ;
        RECT 33.845 -208.405 34.075 -207.405 ;
        RECT 35.655 -208.405 35.885 -207.405 ;
        RECT 36.635 -208.405 36.865 -207.405 ;
        RECT 38.185 -208.405 38.415 -207.405 ;
        RECT 39.730 -208.405 39.960 -207.405 ;
        RECT 12.635 -210.370 13.410 -210.360 ;
        RECT -33.870 -210.405 13.410 -210.370 ;
        RECT -34.490 -210.580 13.410 -210.405 ;
        RECT -34.490 -210.635 -33.810 -210.580 ;
        RECT 12.635 -210.590 13.410 -210.580 ;
        RECT -22.090 -210.780 -21.410 -210.770 ;
        RECT -22.090 -210.990 13.835 -210.780 ;
        RECT -22.090 -211.000 -21.410 -210.990 ;
        RECT 13.155 -211.010 13.835 -210.990 ;
        RECT 47.340 -211.585 47.595 -202.910 ;
        RECT -23.565 -211.815 47.595 -211.585 ;
        RECT -23.565 -211.840 45.475 -211.815 ;
        RECT -33.765 -216.630 -33.535 -215.630 ;
        RECT -33.275 -216.630 -33.045 -215.630 ;
        RECT -31.695 -216.630 -31.465 -215.630 ;
        RECT -31.205 -216.630 -30.975 -215.630 ;
        RECT -29.885 -216.630 -29.655 -215.630 ;
        RECT -29.395 -216.630 -29.165 -215.630 ;
        RECT -28.415 -216.630 -28.185 -215.630 ;
        RECT -27.925 -216.630 -27.695 -215.630 ;
        RECT -26.865 -216.630 -26.635 -215.630 ;
        RECT -26.375 -216.630 -26.145 -215.630 ;
        RECT -25.320 -216.630 -25.090 -215.630 ;
        RECT -24.830 -216.630 -24.600 -215.630 ;
        RECT -27.340 -216.820 -26.685 -216.790 ;
        RECT -32.110 -216.960 -26.685 -216.820 ;
        RECT -33.740 -217.685 -33.045 -217.620 ;
        RECT -32.110 -217.685 -31.970 -216.960 ;
        RECT -27.340 -217.020 -26.685 -216.960 ;
        RECT -33.740 -217.825 -31.970 -217.685 ;
        RECT -29.995 -217.555 -29.300 -217.470 ;
        RECT -25.810 -217.555 -25.130 -217.510 ;
        RECT -29.995 -217.695 -25.130 -217.555 ;
        RECT -29.995 -217.740 -29.300 -217.695 ;
        RECT -25.810 -217.740 -25.130 -217.695 ;
        RECT -33.740 -217.890 -33.045 -217.825 ;
        RECT -27.950 -217.880 -27.255 -217.840 ;
        RECT -24.875 -217.880 -24.180 -217.810 ;
        RECT -23.565 -217.880 -23.425 -211.840 ;
        RECT 46.415 -211.995 47.155 -211.955 ;
        RECT 47.770 -211.995 47.950 -183.635 ;
        RECT 48.120 -206.395 48.375 -183.295 ;
        RECT 48.090 -207.090 48.435 -206.395 ;
        RECT -11.140 -212.175 47.950 -211.995 ;
        RECT -22.105 -212.945 -21.875 -212.265 ;
        RECT -22.100 -215.795 -21.880 -212.945 ;
        RECT -22.105 -216.475 -21.875 -215.795 ;
        RECT -21.265 -216.630 -21.035 -215.630 ;
        RECT -20.775 -216.630 -20.545 -215.630 ;
        RECT -19.195 -216.630 -18.965 -215.630 ;
        RECT -18.705 -216.630 -18.475 -215.630 ;
        RECT -17.385 -216.630 -17.155 -215.630 ;
        RECT -16.895 -216.630 -16.665 -215.630 ;
        RECT -15.915 -216.630 -15.685 -215.630 ;
        RECT -15.425 -216.630 -15.195 -215.630 ;
        RECT -14.365 -216.630 -14.135 -215.630 ;
        RECT -13.875 -216.630 -13.645 -215.630 ;
        RECT -12.820 -216.630 -12.590 -215.630 ;
        RECT -12.330 -216.630 -12.100 -215.630 ;
        RECT -14.840 -216.820 -14.185 -216.790 ;
        RECT -19.610 -216.960 -14.185 -216.820 ;
        RECT -27.950 -218.020 -23.425 -217.880 ;
        RECT -21.240 -217.685 -20.545 -217.620 ;
        RECT -19.610 -217.685 -19.470 -216.960 ;
        RECT -14.840 -217.020 -14.185 -216.960 ;
        RECT -19.330 -217.185 -18.635 -217.100 ;
        RECT -13.940 -217.185 -13.245 -217.070 ;
        RECT -19.330 -217.195 -13.245 -217.185 ;
        RECT -11.140 -217.195 -11.000 -212.175 ;
        RECT 46.415 -212.195 47.155 -212.175 ;
        RECT 48.120 -212.335 48.375 -207.090 ;
        RECT -19.330 -217.325 -11.000 -217.195 ;
        RECT -19.330 -217.370 -18.635 -217.325 ;
        RECT -13.940 -217.335 -11.000 -217.325 ;
        RECT -10.710 -212.490 48.375 -212.335 ;
        RECT -10.710 -212.590 45.475 -212.490 ;
        RECT 46.440 -212.525 48.375 -212.490 ;
        RECT -13.940 -217.340 -13.245 -217.335 ;
        RECT -21.240 -217.825 -19.470 -217.685 ;
        RECT -17.495 -217.555 -16.800 -217.470 ;
        RECT -13.310 -217.555 -12.630 -217.510 ;
        RECT -17.495 -217.695 -12.630 -217.555 ;
        RECT -17.495 -217.740 -16.800 -217.695 ;
        RECT -13.310 -217.740 -12.630 -217.695 ;
        RECT -21.240 -217.890 -20.545 -217.825 ;
        RECT -15.450 -217.880 -14.755 -217.840 ;
        RECT -12.375 -217.880 -11.680 -217.810 ;
        RECT -10.710 -217.880 -10.570 -212.590 ;
        RECT 45.615 -212.730 46.330 -212.640 ;
        RECT 48.605 -212.730 48.745 -182.900 ;
        RECT 49.030 -200.835 49.170 -182.615 ;
        RECT 48.930 -201.425 49.250 -200.835 ;
        RECT 1.280 -212.870 48.745 -212.730 ;
        RECT -8.540 -214.370 -7.860 -214.365 ;
        RECT -9.365 -214.590 -7.860 -214.370 ;
        RECT -9.360 -215.775 -9.140 -214.590 ;
        RECT -8.540 -214.595 -7.860 -214.590 ;
        RECT -9.365 -216.455 -9.135 -215.775 ;
        RECT -8.765 -216.630 -8.535 -215.630 ;
        RECT -8.275 -216.630 -8.045 -215.630 ;
        RECT -6.695 -216.630 -6.465 -215.630 ;
        RECT -6.205 -216.630 -5.975 -215.630 ;
        RECT -4.885 -216.630 -4.655 -215.630 ;
        RECT -4.395 -216.630 -4.165 -215.630 ;
        RECT -3.415 -216.630 -3.185 -215.630 ;
        RECT -2.925 -216.630 -2.695 -215.630 ;
        RECT -1.865 -216.630 -1.635 -215.630 ;
        RECT -1.375 -216.630 -1.145 -215.630 ;
        RECT -0.320 -216.630 -0.090 -215.630 ;
        RECT 0.170 -216.630 0.400 -215.630 ;
        RECT -2.340 -216.820 -1.685 -216.790 ;
        RECT -7.110 -216.960 -1.685 -216.820 ;
        RECT -15.450 -218.020 -10.570 -217.880 ;
        RECT -8.740 -217.685 -8.045 -217.620 ;
        RECT -7.110 -217.685 -6.970 -216.960 ;
        RECT -2.340 -217.020 -1.685 -216.960 ;
        RECT -6.830 -217.185 -6.135 -217.100 ;
        RECT -1.440 -217.185 -0.745 -217.070 ;
        RECT -6.830 -217.195 -0.745 -217.185 ;
        RECT 1.280 -217.195 1.420 -212.870 ;
        RECT 45.615 -212.875 46.330 -212.870 ;
        RECT 49.030 -213.015 49.170 -201.425 ;
        RECT -6.830 -217.325 1.420 -217.195 ;
        RECT -6.830 -217.370 -6.135 -217.325 ;
        RECT -1.440 -217.335 1.420 -217.325 ;
        RECT 1.650 -213.155 49.170 -213.015 ;
        RECT -1.440 -217.340 -0.745 -217.335 ;
        RECT -8.740 -217.825 -6.970 -217.685 ;
        RECT -4.995 -217.555 -4.300 -217.470 ;
        RECT -0.810 -217.555 -0.130 -217.510 ;
        RECT -4.995 -217.695 -0.130 -217.555 ;
        RECT -4.995 -217.740 -4.300 -217.695 ;
        RECT -0.810 -217.740 -0.130 -217.695 ;
        RECT -8.740 -217.890 -8.045 -217.825 ;
        RECT -2.950 -217.880 -2.255 -217.840 ;
        RECT 0.125 -217.880 0.820 -217.810 ;
        RECT 1.650 -217.880 1.790 -213.155 ;
        RECT 44.985 -213.330 45.705 -213.295 ;
        RECT 49.415 -213.330 49.555 -182.300 ;
        RECT 13.610 -213.470 49.555 -213.330 ;
        RECT 49.740 -189.650 49.930 -181.980 ;
        RECT 49.740 -190.315 49.990 -189.650 ;
        RECT 3.945 -214.305 4.625 -214.300 ;
        RECT 3.040 -214.525 4.625 -214.305 ;
        RECT 3.040 -215.775 3.260 -214.525 ;
        RECT 3.945 -214.530 4.625 -214.525 ;
        RECT 3.035 -216.455 3.265 -215.775 ;
        RECT 3.735 -216.630 3.965 -215.630 ;
        RECT 4.225 -216.630 4.455 -215.630 ;
        RECT 5.805 -216.630 6.035 -215.630 ;
        RECT 6.295 -216.630 6.525 -215.630 ;
        RECT 7.615 -216.630 7.845 -215.630 ;
        RECT 8.105 -216.630 8.335 -215.630 ;
        RECT 9.085 -216.630 9.315 -215.630 ;
        RECT 9.575 -216.630 9.805 -215.630 ;
        RECT 10.635 -216.630 10.865 -215.630 ;
        RECT 11.125 -216.630 11.355 -215.630 ;
        RECT 12.180 -216.630 12.410 -215.630 ;
        RECT 12.670 -216.630 12.900 -215.630 ;
        RECT 10.160 -216.820 10.815 -216.790 ;
        RECT 5.390 -216.960 10.815 -216.820 ;
        RECT -2.950 -218.020 1.790 -217.880 ;
        RECT 3.760 -217.685 4.455 -217.620 ;
        RECT 5.390 -217.685 5.530 -216.960 ;
        RECT 10.160 -217.020 10.815 -216.960 ;
        RECT 5.670 -217.185 6.365 -217.100 ;
        RECT 11.060 -217.185 11.755 -217.070 ;
        RECT 5.670 -217.195 11.755 -217.185 ;
        RECT 13.610 -217.195 13.750 -213.470 ;
        RECT 44.985 -213.530 45.705 -213.470 ;
        RECT 49.740 -213.650 49.930 -190.315 ;
        RECT 5.670 -217.325 13.750 -217.195 ;
        RECT 5.670 -217.370 6.365 -217.325 ;
        RECT 11.060 -217.335 13.750 -217.325 ;
        RECT 14.025 -213.700 42.515 -213.650 ;
        RECT 45.915 -213.700 49.930 -213.650 ;
        RECT 14.025 -213.840 49.930 -213.700 ;
        RECT 11.060 -217.340 11.755 -217.335 ;
        RECT 3.760 -217.825 5.530 -217.685 ;
        RECT 7.505 -217.555 8.200 -217.470 ;
        RECT 11.690 -217.555 12.370 -217.510 ;
        RECT 7.505 -217.695 12.370 -217.555 ;
        RECT 7.505 -217.740 8.200 -217.695 ;
        RECT 11.690 -217.740 12.370 -217.695 ;
        RECT 3.760 -217.890 4.455 -217.825 ;
        RECT 9.550 -217.880 10.245 -217.840 ;
        RECT 12.625 -217.880 13.320 -217.810 ;
        RECT 14.025 -217.880 14.165 -213.840 ;
        RECT 14.860 -214.215 15.540 -213.985 ;
        RECT 15.125 -215.775 15.345 -214.215 ;
        RECT 29.385 -214.295 30.065 -214.065 ;
        RECT 15.120 -216.455 15.350 -215.775 ;
        RECT 16.235 -216.630 16.465 -215.630 ;
        RECT 16.725 -216.630 16.955 -215.630 ;
        RECT 18.305 -216.630 18.535 -215.630 ;
        RECT 18.795 -216.630 19.025 -215.630 ;
        RECT 20.115 -216.630 20.345 -215.630 ;
        RECT 20.605 -216.630 20.835 -215.630 ;
        RECT 21.585 -216.630 21.815 -215.630 ;
        RECT 22.075 -216.630 22.305 -215.630 ;
        RECT 23.135 -216.630 23.365 -215.630 ;
        RECT 23.625 -216.630 23.855 -215.630 ;
        RECT 24.680 -216.630 24.910 -215.630 ;
        RECT 25.170 -216.630 25.400 -215.630 ;
        RECT 29.650 -215.775 29.870 -214.295 ;
        RECT 50.555 -214.365 50.695 -181.265 ;
        RECT 30.550 -214.505 50.695 -214.365 ;
        RECT 29.645 -216.455 29.875 -215.775 ;
        RECT 22.660 -216.820 23.315 -216.790 ;
        RECT 17.890 -216.960 23.315 -216.820 ;
        RECT 9.550 -218.020 14.165 -217.880 ;
        RECT 16.260 -217.685 16.955 -217.620 ;
        RECT 17.890 -217.685 18.030 -216.960 ;
        RECT 22.660 -217.020 23.315 -216.960 ;
        RECT 16.260 -217.825 18.030 -217.685 ;
        RECT 20.005 -217.555 20.700 -217.470 ;
        RECT 24.190 -217.555 24.870 -217.510 ;
        RECT 20.005 -217.695 24.870 -217.555 ;
        RECT 20.005 -217.740 20.700 -217.695 ;
        RECT 24.190 -217.740 24.870 -217.695 ;
        RECT 16.260 -217.890 16.955 -217.825 ;
        RECT 22.050 -217.880 22.745 -217.840 ;
        RECT 25.125 -217.880 25.820 -217.810 ;
        RECT 30.550 -217.880 30.690 -214.505 ;
        RECT 31.235 -216.630 31.465 -215.630 ;
        RECT 31.725 -216.630 31.955 -215.630 ;
        RECT 33.305 -216.630 33.535 -215.630 ;
        RECT 33.795 -216.630 34.025 -215.630 ;
        RECT 35.115 -216.630 35.345 -215.630 ;
        RECT 35.605 -216.630 35.835 -215.630 ;
        RECT 36.585 -216.630 36.815 -215.630 ;
        RECT 37.075 -216.630 37.305 -215.630 ;
        RECT 38.135 -216.630 38.365 -215.630 ;
        RECT 38.625 -216.630 38.855 -215.630 ;
        RECT 39.680 -216.630 39.910 -215.630 ;
        RECT 40.170 -216.630 40.400 -215.630 ;
        RECT 37.660 -216.820 38.315 -216.790 ;
        RECT 32.890 -216.960 38.315 -216.820 ;
        RECT 22.050 -218.020 30.690 -217.880 ;
        RECT 31.260 -217.685 31.955 -217.620 ;
        RECT 32.890 -217.685 33.030 -216.960 ;
        RECT 37.660 -217.020 38.315 -216.960 ;
        RECT 31.260 -217.825 33.030 -217.685 ;
        RECT 35.005 -217.555 35.700 -217.470 ;
        RECT 39.190 -217.555 39.870 -217.510 ;
        RECT 35.005 -217.695 39.870 -217.555 ;
        RECT 35.005 -217.740 35.700 -217.695 ;
        RECT 39.190 -217.740 39.870 -217.695 ;
        RECT 31.260 -217.890 31.955 -217.825 ;
        RECT 37.050 -217.880 37.745 -217.840 ;
        RECT 40.125 -217.880 40.820 -217.810 ;
        RECT 51.335 -217.880 51.475 -177.750 ;
        RECT 37.050 -218.020 51.475 -217.880 ;
        RECT 54.545 -215.880 55.545 -185.600 ;
        RECT 63.865 -203.310 65.210 -160.180 ;
        RECT 68.825 -164.845 394.450 -163.290 ;
        RECT 63.560 -205.015 65.490 -203.310 ;
        RECT 68.825 -204.760 70.080 -164.845 ;
        RECT 71.760 -167.095 348.110 -166.210 ;
        RECT 71.760 -198.510 73.415 -167.095 ;
        RECT 77.320 -169.890 304.565 -168.785 ;
        RECT 77.320 -189.610 77.770 -169.890 ;
        RECT 84.225 -172.675 258.620 -171.545 ;
        RECT 82.265 -175.075 214.495 -173.750 ;
        RECT 80.855 -177.105 172.090 -175.860 ;
        RECT 80.985 -180.505 83.810 -180.500 ;
        RECT 79.560 -181.205 83.810 -180.505 ;
        RECT 132.985 -182.665 165.310 -181.820 ;
        RECT 79.395 -185.815 80.730 -185.425 ;
        RECT 79.395 -186.590 128.965 -185.815 ;
        RECT 79.395 -186.915 80.730 -186.590 ;
        RECT 80.710 -189.135 84.845 -188.380 ;
        RECT 101.375 -189.050 101.605 -188.550 ;
        RECT 101.865 -189.050 102.095 -188.550 ;
        RECT 102.355 -189.050 102.585 -188.550 ;
        RECT 102.845 -189.050 103.075 -188.550 ;
        RECT 103.335 -189.050 103.565 -188.550 ;
        RECT 103.825 -189.050 104.055 -188.550 ;
        RECT 104.315 -189.050 104.545 -188.550 ;
        RECT 104.805 -189.050 105.035 -188.550 ;
        RECT 105.900 -189.475 106.130 -188.475 ;
        RECT 106.880 -189.475 107.110 -188.475 ;
        RECT 107.860 -189.475 108.090 -188.475 ;
        RECT 77.300 -190.430 77.790 -189.610 ;
        RECT 71.240 -200.635 73.810 -198.510 ;
        RECT 77.320 -201.255 77.770 -190.430 ;
        RECT 90.845 -190.645 91.075 -189.645 ;
        RECT 91.335 -190.645 91.565 -189.645 ;
        RECT 91.825 -190.645 92.055 -189.645 ;
        RECT 92.315 -190.645 92.545 -189.645 ;
        RECT 104.175 -189.740 105.020 -189.690 ;
        RECT 108.880 -189.740 109.165 -188.565 ;
        RECT 110.085 -189.475 110.315 -188.475 ;
        RECT 111.065 -189.475 111.295 -188.475 ;
        RECT 112.045 -189.475 112.275 -188.475 ;
        RECT 114.875 -189.050 115.105 -188.550 ;
        RECT 115.365 -189.050 115.595 -188.550 ;
        RECT 115.855 -189.050 116.085 -188.550 ;
        RECT 116.345 -189.050 116.575 -188.550 ;
        RECT 116.835 -189.050 117.065 -188.550 ;
        RECT 117.325 -189.050 117.555 -188.550 ;
        RECT 117.815 -189.050 118.045 -188.550 ;
        RECT 118.305 -189.050 118.535 -188.550 ;
        RECT 119.400 -189.475 119.630 -188.475 ;
        RECT 120.380 -189.475 120.610 -188.475 ;
        RECT 121.360 -189.475 121.590 -188.475 ;
        RECT 100.895 -190.265 101.665 -189.965 ;
        RECT 104.175 -190.025 109.165 -189.740 ;
        RECT 117.675 -189.740 118.520 -189.690 ;
        RECT 122.380 -189.740 122.665 -188.565 ;
        RECT 123.585 -189.475 123.815 -188.475 ;
        RECT 124.565 -189.475 124.795 -188.475 ;
        RECT 125.545 -189.475 125.775 -188.475 ;
        RECT 113.160 -189.850 113.460 -189.820 ;
        RECT 104.175 -190.060 105.020 -190.025 ;
        RECT 112.745 -190.150 113.460 -189.850 ;
        RECT 114.430 -189.955 114.635 -189.950 ;
        RECT 95.025 -190.835 95.235 -190.815 ;
        RECT 94.615 -191.135 95.275 -190.835 ;
        RECT 90.845 -195.465 91.075 -192.465 ;
        RECT 91.905 -195.465 92.135 -192.465 ;
        RECT 92.395 -195.465 92.625 -192.465 ;
        RECT 92.885 -195.465 93.115 -192.465 ;
        RECT 93.450 -195.465 93.680 -192.465 ;
        RECT 93.940 -195.465 94.170 -192.465 ;
        RECT 94.430 -195.465 94.660 -192.465 ;
        RECT 80.020 -200.150 90.570 -199.170 ;
        RECT 89.590 -200.180 90.570 -200.150 ;
        RECT 89.590 -200.950 90.580 -200.180 ;
        RECT 89.555 -201.160 94.740 -200.950 ;
        RECT 77.320 -201.320 87.235 -201.255 ;
        RECT 77.320 -201.530 94.290 -201.320 ;
        RECT 77.320 -201.705 87.235 -201.530 ;
        RECT 90.820 -203.735 91.050 -202.735 ;
        RECT 91.310 -203.735 91.540 -202.735 ;
        RECT 91.800 -203.735 92.030 -202.735 ;
        RECT 92.870 -204.260 93.530 -203.960 ;
        RECT 68.745 -205.910 70.185 -204.760 ;
        RECT 93.305 -204.825 93.515 -204.260 ;
        RECT 94.080 -204.385 94.290 -201.530 ;
        RECT 94.530 -203.965 94.740 -201.160 ;
        RECT 95.025 -201.305 95.235 -191.135 ;
        RECT 95.475 -191.440 100.025 -191.155 ;
        RECT 95.475 -198.195 95.760 -191.440 ;
        RECT 98.260 -192.020 98.920 -191.720 ;
        RECT 98.360 -193.065 98.835 -192.020 ;
        RECT 99.740 -192.045 100.025 -191.440 ;
        RECT 100.895 -191.640 101.125 -190.265 ;
        RECT 101.375 -191.125 101.605 -190.625 ;
        RECT 101.865 -191.125 102.095 -190.625 ;
        RECT 102.355 -191.125 102.585 -190.625 ;
        RECT 102.845 -191.125 103.075 -190.625 ;
        RECT 103.335 -191.125 103.565 -190.625 ;
        RECT 103.825 -191.125 104.055 -190.625 ;
        RECT 104.315 -191.125 104.545 -190.625 ;
        RECT 104.805 -191.125 105.035 -190.625 ;
        RECT 105.900 -190.875 106.130 -190.375 ;
        RECT 106.390 -190.875 106.620 -190.375 ;
        RECT 106.880 -190.875 107.110 -190.375 ;
        RECT 107.370 -190.875 107.600 -190.375 ;
        RECT 107.860 -190.875 108.090 -190.375 ;
        RECT 108.350 -190.875 108.580 -190.375 ;
        RECT 110.085 -190.875 110.315 -190.375 ;
        RECT 110.575 -190.875 110.805 -190.375 ;
        RECT 111.065 -190.875 111.295 -190.375 ;
        RECT 111.555 -190.875 111.785 -190.375 ;
        RECT 112.045 -190.875 112.275 -190.375 ;
        RECT 112.535 -190.875 112.765 -190.375 ;
        RECT 100.895 -191.865 104.990 -191.640 ;
        RECT 100.935 -191.870 104.990 -191.865 ;
        RECT 99.740 -192.330 101.070 -192.045 ;
        RECT 99.875 -192.870 100.535 -192.570 ;
        RECT 98.325 -193.365 99.010 -193.065 ;
        RECT 96.960 -194.165 97.190 -193.665 ;
        RECT 97.450 -194.165 97.680 -193.665 ;
        RECT 97.940 -194.165 98.170 -193.665 ;
        RECT 98.430 -194.165 98.660 -193.665 ;
        RECT 98.920 -194.165 99.150 -193.665 ;
        RECT 99.410 -194.165 99.640 -193.665 ;
        RECT 100.080 -194.010 100.370 -192.870 ;
        RECT 100.080 -194.670 100.380 -194.010 ;
        RECT 100.785 -194.515 101.070 -192.330 ;
        RECT 104.760 -192.700 104.990 -191.870 ;
        RECT 111.425 -192.020 112.110 -191.720 ;
        RECT 104.760 -192.930 108.560 -192.700 ;
        RECT 105.420 -193.415 105.630 -192.930 ;
        RECT 106.400 -193.415 106.610 -192.930 ;
        RECT 107.375 -193.415 107.585 -192.930 ;
        RECT 108.330 -193.415 108.560 -192.930 ;
        RECT 111.580 -193.060 112.055 -192.020 ;
        RECT 111.460 -193.360 112.145 -193.060 ;
        RECT 101.370 -194.165 101.600 -193.665 ;
        RECT 101.860 -194.165 102.090 -193.665 ;
        RECT 102.350 -194.165 102.580 -193.665 ;
        RECT 102.840 -194.165 103.070 -193.665 ;
        RECT 103.330 -194.165 103.560 -193.665 ;
        RECT 103.820 -194.165 104.050 -193.665 ;
        RECT 104.915 -193.915 105.145 -193.415 ;
        RECT 105.405 -193.915 105.635 -193.415 ;
        RECT 105.895 -193.915 106.125 -193.415 ;
        RECT 106.385 -193.915 106.615 -193.415 ;
        RECT 106.875 -193.915 107.105 -193.415 ;
        RECT 107.365 -193.915 107.595 -193.415 ;
        RECT 107.855 -193.915 108.085 -193.415 ;
        RECT 108.330 -193.915 108.575 -193.415 ;
        RECT 110.085 -194.165 110.315 -193.665 ;
        RECT 110.575 -194.165 110.805 -193.665 ;
        RECT 111.065 -194.165 111.295 -193.665 ;
        RECT 111.555 -194.165 111.785 -193.665 ;
        RECT 112.045 -194.165 112.275 -193.665 ;
        RECT 112.535 -194.165 112.765 -193.665 ;
        RECT 113.160 -193.890 113.460 -190.150 ;
        RECT 114.425 -190.255 115.110 -189.955 ;
        RECT 117.675 -190.025 122.665 -189.740 ;
        RECT 117.675 -190.060 118.520 -190.025 ;
        RECT 114.430 -192.680 114.635 -190.255 ;
        RECT 114.875 -191.125 115.105 -190.625 ;
        RECT 115.365 -191.125 115.595 -190.625 ;
        RECT 115.855 -191.125 116.085 -190.625 ;
        RECT 116.345 -191.125 116.575 -190.625 ;
        RECT 116.835 -191.125 117.065 -190.625 ;
        RECT 117.325 -191.125 117.555 -190.625 ;
        RECT 117.815 -191.125 118.045 -190.625 ;
        RECT 118.305 -191.125 118.535 -190.625 ;
        RECT 119.400 -190.875 119.630 -190.375 ;
        RECT 119.890 -190.875 120.120 -190.375 ;
        RECT 120.380 -190.875 120.610 -190.375 ;
        RECT 120.870 -190.875 121.100 -190.375 ;
        RECT 121.360 -190.875 121.590 -190.375 ;
        RECT 121.850 -190.875 122.080 -190.375 ;
        RECT 122.670 -192.580 122.970 -190.245 ;
        RECT 123.585 -190.875 123.815 -190.375 ;
        RECT 124.075 -190.875 124.305 -190.375 ;
        RECT 124.565 -190.875 124.795 -190.375 ;
        RECT 125.055 -190.875 125.285 -190.375 ;
        RECT 125.545 -190.875 125.775 -190.375 ;
        RECT 126.035 -190.875 126.265 -190.375 ;
        RECT 124.410 -191.990 125.095 -191.690 ;
        RECT 114.430 -192.920 122.085 -192.680 ;
        RECT 122.490 -192.880 123.150 -192.580 ;
        RECT 113.160 -194.115 113.465 -193.890 ;
        RECT 104.930 -194.515 105.775 -194.480 ;
        RECT 100.785 -194.800 105.775 -194.515 ;
        RECT 113.165 -194.550 113.465 -194.115 ;
        RECT 114.870 -194.165 115.100 -193.665 ;
        RECT 115.360 -194.165 115.590 -193.665 ;
        RECT 115.850 -194.165 116.080 -193.665 ;
        RECT 116.340 -194.165 116.570 -193.665 ;
        RECT 116.830 -194.165 117.060 -193.665 ;
        RECT 117.320 -194.165 117.550 -193.665 ;
        RECT 118.415 -193.915 118.645 -193.415 ;
        RECT 118.885 -193.510 119.190 -192.920 ;
        RECT 118.905 -193.915 119.135 -193.510 ;
        RECT 119.395 -193.915 119.625 -193.415 ;
        RECT 119.840 -193.520 120.145 -192.920 ;
        RECT 119.885 -193.915 120.115 -193.520 ;
        RECT 120.375 -193.915 120.605 -193.415 ;
        RECT 120.820 -193.510 121.125 -192.920 ;
        RECT 120.865 -193.915 121.095 -193.510 ;
        RECT 121.355 -193.915 121.585 -193.415 ;
        RECT 121.845 -193.690 122.085 -192.920 ;
        RECT 124.545 -193.080 125.020 -191.990 ;
        RECT 126.535 -192.280 126.835 -192.045 ;
        RECT 126.535 -192.600 127.880 -192.280 ;
        RECT 126.535 -192.730 127.265 -192.600 ;
        RECT 124.480 -193.380 125.140 -193.080 ;
        RECT 121.845 -193.915 122.075 -193.690 ;
        RECT 123.585 -194.165 123.815 -193.665 ;
        RECT 124.075 -194.165 124.305 -193.665 ;
        RECT 124.565 -194.165 124.795 -193.665 ;
        RECT 125.055 -194.165 125.285 -193.665 ;
        RECT 125.545 -194.165 125.775 -193.665 ;
        RECT 126.035 -194.165 126.265 -193.665 ;
        RECT 118.430 -194.515 119.275 -194.480 ;
        RECT 97.450 -196.065 97.680 -195.065 ;
        RECT 98.430 -196.065 98.660 -195.065 ;
        RECT 99.410 -196.065 99.640 -195.065 ;
        RECT 100.785 -195.975 101.070 -194.800 ;
        RECT 104.930 -194.850 105.775 -194.800 ;
        RECT 114.285 -194.800 119.275 -194.515 ;
        RECT 101.860 -196.065 102.090 -195.065 ;
        RECT 102.840 -196.065 103.070 -195.065 ;
        RECT 103.820 -196.065 104.050 -195.065 ;
        RECT 104.915 -195.990 105.145 -195.490 ;
        RECT 105.405 -195.990 105.635 -195.490 ;
        RECT 105.895 -195.990 106.125 -195.490 ;
        RECT 106.385 -195.990 106.615 -195.490 ;
        RECT 106.875 -195.990 107.105 -195.490 ;
        RECT 107.365 -195.990 107.595 -195.490 ;
        RECT 107.855 -195.990 108.085 -195.490 ;
        RECT 108.345 -195.990 108.575 -195.490 ;
        RECT 110.575 -196.065 110.805 -195.065 ;
        RECT 111.555 -196.065 111.785 -195.065 ;
        RECT 112.535 -196.065 112.765 -195.065 ;
        RECT 114.285 -195.975 114.570 -194.800 ;
        RECT 118.430 -194.850 119.275 -194.800 ;
        RECT 115.360 -196.065 115.590 -195.065 ;
        RECT 116.340 -196.065 116.570 -195.065 ;
        RECT 117.320 -196.065 117.550 -195.065 ;
        RECT 118.415 -195.990 118.645 -195.490 ;
        RECT 118.905 -195.990 119.135 -195.490 ;
        RECT 119.395 -195.990 119.625 -195.490 ;
        RECT 119.885 -195.990 120.115 -195.490 ;
        RECT 120.375 -195.990 120.605 -195.490 ;
        RECT 120.865 -195.990 121.095 -195.490 ;
        RECT 121.355 -195.990 121.585 -195.490 ;
        RECT 121.845 -195.990 122.075 -195.490 ;
        RECT 124.075 -196.065 124.305 -195.065 ;
        RECT 125.055 -196.065 125.285 -195.065 ;
        RECT 126.035 -196.065 126.265 -195.065 ;
        RECT 126.815 -196.950 127.265 -192.730 ;
        RECT 107.105 -197.400 127.265 -196.950 ;
        RECT 107.105 -197.855 107.905 -197.400 ;
        RECT 95.475 -198.480 111.835 -198.195 ;
        RECT 107.090 -199.430 107.890 -198.770 ;
        RECT 95.025 -201.515 98.875 -201.305 ;
        RECT 106.575 -201.345 107.235 -201.045 ;
        RECT 95.550 -203.735 95.780 -202.735 ;
        RECT 96.040 -203.735 96.270 -202.735 ;
        RECT 96.530 -203.735 96.760 -202.735 ;
        RECT 95.110 -203.965 95.770 -203.930 ;
        RECT 94.530 -204.175 95.770 -203.965 ;
        RECT 95.110 -204.230 95.770 -204.175 ;
        RECT 96.225 -204.385 96.885 -204.330 ;
        RECT 94.080 -204.595 96.885 -204.385 ;
        RECT 96.225 -204.630 96.885 -204.595 ;
        RECT 98.050 -204.825 98.350 -204.675 ;
        RECT 93.305 -205.035 98.350 -204.825 ;
        RECT 90.820 -207.195 91.050 -205.195 ;
        RECT 91.875 -207.195 92.105 -205.195 ;
        RECT 92.365 -207.195 92.595 -205.195 ;
        RECT 92.855 -207.195 93.085 -205.195 ;
        RECT 95.550 -207.195 95.780 -205.195 ;
        RECT 96.605 -207.195 96.835 -205.195 ;
        RECT 97.095 -207.195 97.325 -205.195 ;
        RECT 97.585 -207.195 97.815 -205.195 ;
        RECT 98.050 -205.335 98.350 -205.035 ;
        RECT 98.665 -205.925 98.875 -201.515 ;
        RECT 99.640 -204.330 99.870 -202.830 ;
        RECT 100.130 -204.330 100.360 -202.830 ;
        RECT 100.620 -204.330 100.850 -202.830 ;
        RECT 101.190 -204.325 101.420 -202.825 ;
        RECT 101.680 -204.325 101.910 -202.825 ;
        RECT 102.170 -204.325 102.400 -202.825 ;
        RECT 102.735 -204.325 102.965 -202.825 ;
        RECT 103.225 -204.325 103.455 -202.825 ;
        RECT 103.715 -204.325 103.945 -202.825 ;
        RECT 105.290 -203.825 105.520 -202.825 ;
        RECT 105.780 -203.825 106.010 -202.825 ;
        RECT 106.735 -204.770 107.035 -201.345 ;
        RECT 107.430 -201.550 107.730 -199.430 ;
        RECT 109.675 -200.825 109.905 -198.825 ;
        RECT 110.655 -200.825 110.885 -198.825 ;
        RECT 111.550 -201.090 111.835 -198.480 ;
        RECT 128.190 -198.535 128.965 -186.590 ;
        RECT 112.530 -198.885 128.965 -198.535 ;
        RECT 112.530 -199.780 112.880 -198.885 ;
        RECT 107.430 -201.555 109.135 -201.550 ;
        RECT 107.430 -201.845 109.140 -201.555 ;
        RECT 111.405 -201.760 111.835 -201.090 ;
        RECT 107.430 -201.850 109.135 -201.845 ;
        RECT 106.540 -205.070 107.195 -204.770 ;
        RECT 107.430 -205.620 107.730 -201.850 ;
        RECT 109.185 -203.095 109.415 -202.095 ;
        RECT 109.675 -203.095 109.905 -202.095 ;
        RECT 110.235 -203.095 110.465 -202.095 ;
        RECT 110.725 -203.095 110.955 -202.095 ;
        RECT 113.335 -202.550 113.565 -199.050 ;
        RECT 113.825 -202.550 114.055 -199.050 ;
        RECT 115.335 -202.550 115.565 -199.050 ;
        RECT 115.825 -202.550 116.055 -199.050 ;
        RECT 117.750 -202.535 118.100 -198.885 ;
        RECT 118.335 -202.550 118.565 -199.050 ;
        RECT 118.825 -202.550 119.055 -199.050 ;
        RECT 120.335 -202.550 120.565 -199.050 ;
        RECT 120.825 -202.550 121.055 -199.050 ;
        RECT 122.705 -202.540 123.055 -198.885 ;
        RECT 123.335 -202.550 123.565 -199.050 ;
        RECT 123.825 -202.550 124.055 -199.050 ;
        RECT 125.335 -202.550 125.565 -199.050 ;
        RECT 125.825 -202.550 126.055 -199.050 ;
        RECT 132.985 -200.905 133.830 -182.665 ;
        RECT 143.110 -183.990 145.305 -183.755 ;
        RECT 143.110 -184.175 143.345 -183.990 ;
        RECT 137.310 -186.540 137.960 -185.790 ;
        RECT 138.740 -186.060 138.970 -185.060 ;
        RECT 139.230 -186.200 139.460 -185.060 ;
        RECT 139.720 -186.060 139.950 -185.060 ;
        RECT 140.210 -186.200 140.440 -185.060 ;
        RECT 143.115 -185.670 143.345 -184.175 ;
        RECT 143.605 -185.670 143.835 -184.170 ;
        RECT 144.095 -185.670 144.325 -183.990 ;
        RECT 138.740 -186.430 141.925 -186.200 ;
        RECT 137.560 -193.560 137.830 -186.540 ;
        RECT 138.740 -187.710 138.970 -186.430 ;
        RECT 139.230 -186.440 140.440 -186.430 ;
        RECT 139.720 -187.710 139.950 -186.440 ;
        RECT 140.700 -187.710 140.930 -186.430 ;
        RECT 143.605 -188.355 143.835 -186.855 ;
        RECT 144.585 -188.355 144.815 -184.170 ;
        RECT 145.075 -185.670 145.305 -183.990 ;
        RECT 148.585 -186.530 152.125 -185.965 ;
        RECT 146.650 -187.205 146.880 -186.705 ;
        RECT 147.140 -187.350 147.370 -186.705 ;
        RECT 147.630 -187.205 147.860 -186.705 ;
        RECT 148.120 -187.350 148.350 -186.705 ;
        RECT 146.650 -187.580 149.835 -187.350 ;
        RECT 146.650 -188.360 146.880 -187.580 ;
        RECT 147.140 -187.590 148.350 -187.580 ;
        RECT 147.630 -188.360 147.860 -187.590 ;
        RECT 148.610 -188.360 148.840 -187.580 ;
        RECT 138.610 -192.855 138.840 -191.355 ;
        RECT 136.845 -193.830 137.830 -193.560 ;
        RECT 138.120 -195.535 138.350 -194.040 ;
        RECT 138.115 -195.720 138.350 -195.535 ;
        RECT 138.610 -195.540 138.840 -194.040 ;
        RECT 139.100 -195.720 139.330 -194.040 ;
        RECT 139.590 -195.540 139.820 -191.355 ;
        RECT 141.655 -192.130 141.885 -191.350 ;
        RECT 142.635 -192.120 142.865 -191.350 ;
        RECT 142.145 -192.130 143.355 -192.120 ;
        RECT 143.615 -192.130 143.845 -191.350 ;
        RECT 141.655 -192.360 144.840 -192.130 ;
        RECT 141.655 -193.005 141.885 -192.505 ;
        RECT 142.145 -193.005 142.375 -192.360 ;
        RECT 142.635 -193.005 142.865 -192.505 ;
        RECT 143.125 -193.005 143.355 -192.360 ;
        RECT 145.845 -193.910 146.075 -190.910 ;
        RECT 146.900 -193.910 147.130 -190.910 ;
        RECT 147.390 -193.910 147.620 -190.910 ;
        RECT 147.880 -193.910 148.110 -190.910 ;
        RECT 148.940 -193.910 149.170 -190.910 ;
        RECT 140.080 -195.720 140.310 -194.040 ;
        RECT 150.095 -194.565 150.620 -194.205 ;
        RECT 150.125 -194.980 150.450 -194.565 ;
        RECT 145.350 -195.305 150.450 -194.980 ;
        RECT 138.115 -195.955 140.310 -195.720 ;
        RECT 145.845 -196.970 146.075 -195.470 ;
        RECT 146.335 -196.970 146.565 -195.470 ;
        RECT 146.825 -196.970 147.055 -195.470 ;
        RECT 148.035 -196.970 148.265 -195.470 ;
        RECT 148.525 -196.970 148.755 -195.470 ;
        RECT 149.690 -197.510 150.255 -197.505 ;
        RECT 151.560 -197.510 152.125 -186.530 ;
        RECT 155.805 -192.700 156.035 -190.200 ;
        RECT 157.150 -192.700 157.380 -190.200 ;
        RECT 157.640 -192.700 157.870 -190.200 ;
        RECT 158.130 -192.700 158.360 -190.200 ;
        RECT 158.780 -192.700 159.010 -190.200 ;
        RECT 160.410 -192.700 160.640 -190.200 ;
        RECT 161.550 -191.700 161.780 -190.200 ;
        RECT 154.650 -193.500 155.340 -193.480 ;
        RECT 158.680 -193.500 159.370 -193.480 ;
        RECT 160.605 -193.500 160.875 -193.135 ;
        RECT 154.650 -193.720 160.875 -193.500 ;
        RECT 154.650 -193.750 155.340 -193.720 ;
        RECT 158.680 -193.750 159.370 -193.720 ;
        RECT 160.605 -193.825 160.875 -193.720 ;
        RECT 161.465 -193.900 161.795 -193.840 ;
        RECT 164.465 -193.900 165.310 -182.665 ;
        RECT 170.845 -183.275 172.090 -177.105 ;
        RECT 172.900 -182.405 208.310 -181.450 ;
        RECT 170.390 -183.955 172.175 -183.275 ;
        RECT 170.390 -184.225 172.205 -183.955 ;
        RECT 170.390 -184.610 172.175 -184.225 ;
        RECT 153.845 -195.435 154.360 -194.980 ;
        RECT 148.740 -198.075 152.125 -197.510 ;
        RECT 132.985 -201.335 134.735 -200.905 ;
        RECT 143.070 -201.255 145.265 -201.020 ;
        RECT 132.985 -201.605 141.625 -201.335 ;
        RECT 143.070 -201.440 143.305 -201.255 ;
        RECT 132.985 -201.750 134.735 -201.605 ;
        RECT 116.395 -202.800 116.985 -202.740 ;
        RECT 116.395 -202.970 117.430 -202.800 ;
        RECT 126.260 -202.835 126.850 -202.815 ;
        RECT 129.015 -202.835 129.620 -202.720 ;
        RECT 116.395 -203.030 116.985 -202.970 ;
        RECT 108.935 -205.430 109.165 -204.930 ;
        RECT 109.425 -205.430 109.655 -204.930 ;
        RECT 109.915 -205.430 110.145 -204.930 ;
        RECT 110.405 -205.430 110.635 -204.930 ;
        RECT 110.895 -205.430 111.125 -204.930 ;
        RECT 111.385 -205.430 111.615 -204.930 ;
        RECT 107.430 -205.920 109.065 -205.620 ;
        RECT 98.625 -206.585 98.925 -205.925 ;
        RECT 100.130 -207.365 100.360 -206.365 ;
        RECT 101.110 -207.365 101.340 -206.365 ;
        RECT 102.090 -207.365 102.320 -206.365 ;
        RECT 105.780 -207.365 106.010 -206.365 ;
        RECT 109.425 -207.330 109.655 -206.330 ;
        RECT 110.405 -207.330 110.635 -206.330 ;
        RECT 111.385 -207.330 111.615 -206.330 ;
        RECT 113.825 -206.975 114.055 -203.475 ;
        RECT 115.825 -206.975 116.055 -203.475 ;
        RECT 117.260 -207.475 117.430 -202.970 ;
        RECT 121.780 -203.165 122.370 -202.875 ;
        RECT 126.260 -203.060 129.620 -202.835 ;
        RECT 126.260 -203.105 126.850 -203.060 ;
        RECT 118.825 -206.975 119.055 -203.475 ;
        RECT 120.825 -206.975 121.055 -203.475 ;
        RECT 121.810 -207.150 121.980 -203.165 ;
        RECT 123.825 -206.975 124.055 -203.475 ;
        RECT 125.825 -206.975 126.055 -203.475 ;
        RECT 121.810 -207.320 128.350 -207.150 ;
        RECT 117.260 -207.645 127.910 -207.475 ;
        RECT 56.810 -212.255 57.040 -211.255 ;
        RECT 57.790 -212.255 58.020 -211.255 ;
        RECT 58.770 -212.255 59.000 -211.255 ;
        RECT 60.145 -212.520 60.430 -211.345 ;
        RECT 61.220 -212.255 61.450 -211.255 ;
        RECT 62.200 -212.255 62.430 -211.255 ;
        RECT 63.180 -212.255 63.410 -211.255 ;
        RECT 64.275 -211.830 64.505 -211.330 ;
        RECT 64.765 -211.830 64.995 -211.330 ;
        RECT 65.255 -211.830 65.485 -211.330 ;
        RECT 65.745 -211.830 65.975 -211.330 ;
        RECT 66.235 -211.830 66.465 -211.330 ;
        RECT 66.725 -211.830 66.955 -211.330 ;
        RECT 67.215 -211.830 67.445 -211.330 ;
        RECT 67.705 -211.830 67.935 -211.330 ;
        RECT 69.935 -212.255 70.165 -211.255 ;
        RECT 70.915 -212.255 71.145 -211.255 ;
        RECT 71.895 -212.255 72.125 -211.255 ;
        RECT 64.290 -212.520 65.135 -212.470 ;
        RECT 56.320 -213.655 56.550 -213.155 ;
        RECT 56.810 -213.655 57.040 -213.155 ;
        RECT 57.300 -213.655 57.530 -213.155 ;
        RECT 57.790 -213.655 58.020 -213.155 ;
        RECT 58.280 -213.655 58.510 -213.155 ;
        RECT 58.770 -213.655 59.000 -213.155 ;
        RECT 59.440 -213.310 59.740 -212.650 ;
        RECT 60.145 -212.805 65.135 -212.520 ;
        RECT 73.645 -212.520 73.930 -211.345 ;
        RECT 74.720 -212.255 74.950 -211.255 ;
        RECT 75.700 -212.255 75.930 -211.255 ;
        RECT 76.680 -212.255 76.910 -211.255 ;
        RECT 77.775 -211.830 78.005 -211.330 ;
        RECT 78.265 -211.830 78.495 -211.330 ;
        RECT 78.755 -211.830 78.985 -211.330 ;
        RECT 79.245 -211.830 79.475 -211.330 ;
        RECT 79.735 -211.830 79.965 -211.330 ;
        RECT 80.225 -211.830 80.455 -211.330 ;
        RECT 80.715 -211.830 80.945 -211.330 ;
        RECT 81.205 -211.830 81.435 -211.330 ;
        RECT 83.435 -212.255 83.665 -211.255 ;
        RECT 84.415 -212.255 84.645 -211.255 ;
        RECT 85.395 -212.255 85.625 -211.255 ;
        RECT 77.790 -212.520 78.635 -212.470 ;
        RECT 57.685 -214.255 58.370 -213.955 ;
        RECT 57.720 -215.300 58.195 -214.255 ;
        RECT 59.440 -214.450 59.730 -213.310 ;
        RECT 59.235 -214.750 59.895 -214.450 ;
        RECT 60.145 -214.990 60.430 -212.805 ;
        RECT 64.290 -212.840 65.135 -212.805 ;
        RECT 60.730 -213.655 60.960 -213.155 ;
        RECT 61.220 -213.655 61.450 -213.155 ;
        RECT 61.710 -213.655 61.940 -213.155 ;
        RECT 62.200 -213.655 62.430 -213.155 ;
        RECT 62.690 -213.655 62.920 -213.155 ;
        RECT 63.180 -213.655 63.410 -213.155 ;
        RECT 64.275 -213.905 64.505 -213.405 ;
        RECT 64.765 -213.905 64.995 -213.405 ;
        RECT 65.255 -213.905 65.485 -213.405 ;
        RECT 65.745 -213.905 65.975 -213.405 ;
        RECT 66.235 -213.905 66.465 -213.405 ;
        RECT 66.725 -213.905 66.955 -213.405 ;
        RECT 67.215 -213.905 67.445 -213.405 ;
        RECT 67.690 -213.905 67.935 -213.405 ;
        RECT 69.445 -213.655 69.675 -213.155 ;
        RECT 69.935 -213.655 70.165 -213.155 ;
        RECT 70.425 -213.655 70.655 -213.155 ;
        RECT 70.915 -213.655 71.145 -213.155 ;
        RECT 71.405 -213.655 71.635 -213.155 ;
        RECT 71.895 -213.655 72.125 -213.155 ;
        RECT 72.525 -213.205 72.825 -212.770 ;
        RECT 73.645 -212.805 78.635 -212.520 ;
        RECT 77.790 -212.840 78.635 -212.805 ;
        RECT 72.520 -213.430 72.825 -213.205 ;
        RECT 64.780 -214.390 64.990 -213.905 ;
        RECT 65.760 -214.390 65.970 -213.905 ;
        RECT 66.735 -214.390 66.945 -213.905 ;
        RECT 67.690 -214.390 67.920 -213.905 ;
        RECT 70.820 -214.260 71.505 -213.960 ;
        RECT 59.100 -215.275 60.430 -214.990 ;
        RECT 64.120 -214.620 67.920 -214.390 ;
        RECT 57.620 -215.600 58.280 -215.300 ;
        RECT 59.100 -215.880 59.385 -215.275 ;
        RECT 64.120 -215.450 64.350 -214.620 ;
        RECT 70.940 -215.300 71.415 -214.260 ;
        RECT 60.295 -215.455 64.350 -215.450 ;
        RECT 54.545 -216.165 59.385 -215.880 ;
        RECT 60.255 -215.680 64.350 -215.455 ;
        RECT 70.785 -215.600 71.470 -215.300 ;
        RECT -27.950 -218.110 -27.255 -218.020 ;
        RECT -24.875 -218.080 -24.180 -218.020 ;
        RECT -15.450 -218.110 -14.755 -218.020 ;
        RECT -12.375 -218.080 -11.680 -218.020 ;
        RECT -2.950 -218.110 -2.255 -218.020 ;
        RECT 0.125 -218.080 0.820 -218.020 ;
        RECT 9.550 -218.110 10.245 -218.020 ;
        RECT 12.625 -218.080 13.320 -218.020 ;
        RECT 22.050 -218.110 22.745 -218.020 ;
        RECT 25.125 -218.080 25.820 -218.020 ;
        RECT 37.050 -218.110 37.745 -218.020 ;
        RECT 40.125 -218.080 40.820 -218.020 ;
        RECT -33.765 -219.660 -33.535 -218.660 ;
        RECT -33.275 -219.660 -33.045 -218.660 ;
        RECT -32.785 -219.660 -32.555 -218.660 ;
        RECT -32.185 -219.660 -31.955 -218.660 ;
        RECT -31.695 -219.660 -31.465 -218.660 ;
        RECT -31.205 -219.660 -30.975 -218.660 ;
        RECT -29.395 -219.660 -29.165 -218.660 ;
        RECT -28.415 -219.660 -28.185 -218.660 ;
        RECT -26.865 -219.660 -26.635 -218.660 ;
        RECT -25.320 -219.660 -25.090 -218.660 ;
        RECT -21.265 -219.660 -21.035 -218.660 ;
        RECT -20.775 -219.660 -20.545 -218.660 ;
        RECT -20.285 -219.660 -20.055 -218.660 ;
        RECT -19.685 -219.660 -19.455 -218.660 ;
        RECT -19.195 -219.660 -18.965 -218.660 ;
        RECT -18.705 -219.660 -18.475 -218.660 ;
        RECT -16.895 -219.660 -16.665 -218.660 ;
        RECT -15.915 -219.660 -15.685 -218.660 ;
        RECT -14.365 -219.660 -14.135 -218.660 ;
        RECT -12.820 -219.660 -12.590 -218.660 ;
        RECT -8.765 -219.660 -8.535 -218.660 ;
        RECT -8.275 -219.660 -8.045 -218.660 ;
        RECT -7.785 -219.660 -7.555 -218.660 ;
        RECT -7.185 -219.660 -6.955 -218.660 ;
        RECT -6.695 -219.660 -6.465 -218.660 ;
        RECT -6.205 -219.660 -5.975 -218.660 ;
        RECT -4.395 -219.660 -4.165 -218.660 ;
        RECT -3.415 -219.660 -3.185 -218.660 ;
        RECT -1.865 -219.660 -1.635 -218.660 ;
        RECT -0.320 -219.660 -0.090 -218.660 ;
        RECT 3.735 -219.660 3.965 -218.660 ;
        RECT 4.225 -219.660 4.455 -218.660 ;
        RECT 4.715 -219.660 4.945 -218.660 ;
        RECT 5.315 -219.660 5.545 -218.660 ;
        RECT 5.805 -219.660 6.035 -218.660 ;
        RECT 6.295 -219.660 6.525 -218.660 ;
        RECT 8.105 -219.660 8.335 -218.660 ;
        RECT 9.085 -219.660 9.315 -218.660 ;
        RECT 10.635 -219.660 10.865 -218.660 ;
        RECT 12.180 -219.660 12.410 -218.660 ;
        RECT 16.235 -219.660 16.465 -218.660 ;
        RECT 16.725 -219.660 16.955 -218.660 ;
        RECT 17.215 -219.660 17.445 -218.660 ;
        RECT 17.815 -219.660 18.045 -218.660 ;
        RECT 18.305 -219.660 18.535 -218.660 ;
        RECT 18.795 -219.660 19.025 -218.660 ;
        RECT 20.605 -219.660 20.835 -218.660 ;
        RECT 21.585 -219.660 21.815 -218.660 ;
        RECT 23.135 -219.660 23.365 -218.660 ;
        RECT 24.680 -219.660 24.910 -218.660 ;
        RECT 31.235 -219.660 31.465 -218.660 ;
        RECT 31.725 -219.660 31.955 -218.660 ;
        RECT 32.215 -219.660 32.445 -218.660 ;
        RECT 32.815 -219.660 33.045 -218.660 ;
        RECT 33.305 -219.660 33.535 -218.660 ;
        RECT 33.795 -219.660 34.025 -218.660 ;
        RECT 35.605 -219.660 35.835 -218.660 ;
        RECT 36.585 -219.660 36.815 -218.660 ;
        RECT 38.135 -219.660 38.365 -218.660 ;
        RECT 39.680 -219.660 39.910 -218.660 ;
        RECT -95.030 -221.385 -94.340 -220.700 ;
        RECT -36.555 -221.475 -35.740 -220.600 ;
        RECT -95.720 -221.875 -95.035 -221.585 ;
        RECT -112.160 -231.395 -111.545 -230.780 ;
        RECT -36.500 -233.250 -35.840 -221.475 ;
        RECT 44.825 -227.415 45.130 -220.530 ;
        RECT 44.480 -227.420 45.130 -227.415 ;
        RECT 44.480 -227.585 45.135 -227.420 ;
        RECT 44.485 -228.010 45.135 -227.585 ;
        RECT 45.395 -228.055 45.715 -220.510 ;
        RECT 45.385 -228.915 45.715 -228.055 ;
        RECT 45.280 -228.920 45.715 -228.915 ;
        RECT 45.280 -229.535 45.895 -228.920 ;
        RECT 46.120 -230.755 46.420 -220.330 ;
        RECT 46.035 -231.370 46.650 -230.755 ;
        RECT -36.500 -233.930 -35.820 -233.250 ;
        RECT 54.545 -235.115 55.545 -216.165 ;
        RECT 60.255 -217.055 60.485 -215.680 ;
        RECT 60.735 -216.695 60.965 -216.195 ;
        RECT 61.225 -216.695 61.455 -216.195 ;
        RECT 61.715 -216.695 61.945 -216.195 ;
        RECT 62.205 -216.695 62.435 -216.195 ;
        RECT 62.695 -216.695 62.925 -216.195 ;
        RECT 63.185 -216.695 63.415 -216.195 ;
        RECT 63.675 -216.695 63.905 -216.195 ;
        RECT 64.165 -216.695 64.395 -216.195 ;
        RECT 65.260 -216.945 65.490 -216.445 ;
        RECT 65.750 -216.945 65.980 -216.445 ;
        RECT 66.240 -216.945 66.470 -216.445 ;
        RECT 66.730 -216.945 66.960 -216.445 ;
        RECT 67.220 -216.945 67.450 -216.445 ;
        RECT 67.710 -216.945 67.940 -216.445 ;
        RECT 69.445 -216.945 69.675 -216.445 ;
        RECT 69.935 -216.945 70.165 -216.445 ;
        RECT 70.425 -216.945 70.655 -216.445 ;
        RECT 70.915 -216.945 71.145 -216.445 ;
        RECT 71.405 -216.945 71.635 -216.445 ;
        RECT 71.895 -216.945 72.125 -216.445 ;
        RECT 60.255 -217.355 61.025 -217.055 ;
        RECT 72.520 -217.170 72.820 -213.430 ;
        RECT 74.230 -213.655 74.460 -213.155 ;
        RECT 74.720 -213.655 74.950 -213.155 ;
        RECT 75.210 -213.655 75.440 -213.155 ;
        RECT 75.700 -213.655 75.930 -213.155 ;
        RECT 76.190 -213.655 76.420 -213.155 ;
        RECT 76.680 -213.655 76.910 -213.155 ;
        RECT 77.775 -213.905 78.005 -213.405 ;
        RECT 78.265 -213.810 78.495 -213.405 ;
        RECT 78.245 -214.400 78.550 -213.810 ;
        RECT 78.755 -213.905 78.985 -213.405 ;
        RECT 79.245 -213.800 79.475 -213.405 ;
        RECT 79.200 -214.400 79.505 -213.800 ;
        RECT 79.735 -213.905 79.965 -213.405 ;
        RECT 80.225 -213.810 80.455 -213.405 ;
        RECT 80.180 -214.400 80.485 -213.810 ;
        RECT 80.715 -213.905 80.945 -213.405 ;
        RECT 81.205 -213.630 81.435 -213.405 ;
        RECT 81.205 -214.400 81.445 -213.630 ;
        RECT 82.945 -213.655 83.175 -213.155 ;
        RECT 83.435 -213.655 83.665 -213.155 ;
        RECT 83.925 -213.655 84.155 -213.155 ;
        RECT 84.415 -213.655 84.645 -213.155 ;
        RECT 84.905 -213.655 85.135 -213.155 ;
        RECT 85.395 -213.655 85.625 -213.155 ;
        RECT 83.840 -214.240 84.500 -213.940 ;
        RECT 73.790 -214.640 81.445 -214.400 ;
        RECT 73.790 -217.065 73.995 -214.640 ;
        RECT 81.850 -214.740 82.510 -214.440 ;
        RECT 74.235 -216.695 74.465 -216.195 ;
        RECT 74.725 -216.695 74.955 -216.195 ;
        RECT 75.215 -216.695 75.445 -216.195 ;
        RECT 75.705 -216.695 75.935 -216.195 ;
        RECT 76.195 -216.695 76.425 -216.195 ;
        RECT 76.685 -216.695 76.915 -216.195 ;
        RECT 77.175 -216.695 77.405 -216.195 ;
        RECT 77.665 -216.695 77.895 -216.195 ;
        RECT 78.760 -216.945 78.990 -216.445 ;
        RECT 79.250 -216.945 79.480 -216.445 ;
        RECT 79.740 -216.945 79.970 -216.445 ;
        RECT 80.230 -216.945 80.460 -216.445 ;
        RECT 80.720 -216.945 80.950 -216.445 ;
        RECT 81.210 -216.945 81.440 -216.445 ;
        RECT 63.535 -217.295 64.380 -217.260 ;
        RECT 63.535 -217.580 68.525 -217.295 ;
        RECT 72.105 -217.470 72.820 -217.170 ;
        RECT 73.785 -217.365 74.470 -217.065 ;
        RECT 82.030 -217.075 82.330 -214.740 ;
        RECT 83.905 -215.330 84.380 -214.240 ;
        RECT 85.895 -214.720 86.195 -214.590 ;
        RECT 85.895 -215.040 88.175 -214.720 ;
        RECT 85.895 -215.275 86.195 -215.040 ;
        RECT 83.770 -215.630 84.455 -215.330 ;
        RECT 82.945 -216.945 83.175 -216.445 ;
        RECT 83.435 -216.945 83.665 -216.445 ;
        RECT 83.925 -216.945 84.155 -216.445 ;
        RECT 84.415 -216.945 84.645 -216.445 ;
        RECT 84.905 -216.945 85.135 -216.445 ;
        RECT 85.395 -216.945 85.625 -216.445 ;
        RECT 77.035 -217.295 77.880 -217.260 ;
        RECT 73.790 -217.370 73.995 -217.365 ;
        RECT 72.520 -217.500 72.820 -217.470 ;
        RECT 63.535 -217.630 64.380 -217.580 ;
        RECT 60.735 -218.770 60.965 -218.270 ;
        RECT 61.225 -218.770 61.455 -218.270 ;
        RECT 61.715 -218.770 61.945 -218.270 ;
        RECT 62.205 -218.770 62.435 -218.270 ;
        RECT 62.695 -218.770 62.925 -218.270 ;
        RECT 63.185 -218.770 63.415 -218.270 ;
        RECT 63.675 -218.770 63.905 -218.270 ;
        RECT 64.165 -218.770 64.395 -218.270 ;
        RECT 65.260 -218.845 65.490 -217.845 ;
        RECT 66.240 -218.845 66.470 -217.845 ;
        RECT 67.220 -218.845 67.450 -217.845 ;
        RECT 68.240 -218.755 68.525 -217.580 ;
        RECT 77.035 -217.580 82.025 -217.295 ;
        RECT 77.035 -217.630 77.880 -217.580 ;
        RECT 69.445 -218.845 69.675 -217.845 ;
        RECT 70.425 -218.845 70.655 -217.845 ;
        RECT 71.405 -218.845 71.635 -217.845 ;
        RECT 74.235 -218.770 74.465 -218.270 ;
        RECT 74.725 -218.770 74.955 -218.270 ;
        RECT 75.215 -218.770 75.445 -218.270 ;
        RECT 75.705 -218.770 75.935 -218.270 ;
        RECT 76.195 -218.770 76.425 -218.270 ;
        RECT 76.685 -218.770 76.915 -218.270 ;
        RECT 77.175 -218.770 77.405 -218.270 ;
        RECT 77.665 -218.770 77.895 -218.270 ;
        RECT 78.760 -218.845 78.990 -217.845 ;
        RECT 79.740 -218.845 79.970 -217.845 ;
        RECT 80.720 -218.845 80.950 -217.845 ;
        RECT 81.740 -218.755 82.025 -217.580 ;
        RECT 82.945 -218.845 83.175 -217.845 ;
        RECT 83.925 -218.845 84.155 -217.845 ;
        RECT 84.905 -218.845 85.135 -217.845 ;
        RECT 87.535 -233.250 88.175 -215.040 ;
        RECT 125.045 -218.500 125.395 -207.645 ;
        RECT 128.180 -207.960 128.350 -207.320 ;
        RECT 124.450 -219.600 126.305 -218.500 ;
        RECT 127.875 -221.245 128.480 -207.960 ;
        RECT 87.510 -233.930 88.175 -233.250 ;
        RECT 121.475 -221.850 128.480 -221.245 ;
        RECT 121.475 -236.065 122.080 -221.850 ;
        RECT 129.015 -233.055 129.620 -203.060 ;
        RECT 137.270 -203.805 137.920 -203.055 ;
        RECT 138.700 -203.325 138.930 -202.325 ;
        RECT 139.190 -203.465 139.420 -202.325 ;
        RECT 139.680 -203.325 139.910 -202.325 ;
        RECT 140.170 -203.465 140.400 -202.325 ;
        RECT 141.355 -203.055 141.625 -201.605 ;
        RECT 143.075 -202.935 143.305 -201.440 ;
        RECT 143.565 -202.935 143.795 -201.435 ;
        RECT 144.055 -202.935 144.285 -201.255 ;
        RECT 141.355 -203.325 142.995 -203.055 ;
        RECT 138.700 -203.695 141.885 -203.465 ;
        RECT 142.725 -203.600 142.995 -203.325 ;
        RECT 137.520 -210.825 137.790 -203.805 ;
        RECT 138.700 -204.975 138.930 -203.695 ;
        RECT 139.190 -203.705 140.400 -203.695 ;
        RECT 139.680 -204.975 139.910 -203.705 ;
        RECT 140.660 -204.975 140.890 -203.695 ;
        RECT 142.595 -203.890 143.390 -203.600 ;
        RECT 143.565 -205.620 143.795 -204.120 ;
        RECT 144.545 -205.620 144.775 -201.435 ;
        RECT 145.035 -202.935 145.265 -201.255 ;
        RECT 149.690 -203.230 150.255 -198.075 ;
        RECT 153.905 -198.600 154.300 -195.435 ;
        RECT 155.315 -196.680 155.545 -195.180 ;
        RECT 155.805 -196.680 156.035 -195.180 ;
        RECT 157.665 -196.680 157.895 -194.180 ;
        RECT 158.155 -196.680 158.385 -194.180 ;
        RECT 158.780 -196.680 159.010 -194.180 ;
        RECT 159.270 -196.680 159.500 -194.180 ;
        RECT 159.920 -196.680 160.150 -194.180 ;
        RECT 160.410 -196.680 160.640 -194.180 ;
        RECT 160.900 -196.680 161.130 -194.180 ;
        RECT 161.465 -194.210 169.575 -193.900 ;
        RECT 161.465 -194.255 161.795 -194.210 ;
        RECT 161.550 -196.680 161.780 -195.180 ;
        RECT 162.040 -196.680 162.270 -195.180 ;
        RECT 151.405 -198.995 154.300 -198.600 ;
        RECT 151.405 -200.770 151.800 -198.995 ;
        RECT 151.275 -201.255 151.855 -200.770 ;
        RECT 161.410 -201.410 163.605 -201.175 ;
        RECT 154.420 -201.490 154.905 -201.460 ;
        RECT 154.420 -201.760 159.965 -201.490 ;
        RECT 161.410 -201.595 161.645 -201.410 ;
        RECT 154.420 -201.790 154.905 -201.760 ;
        RECT 148.545 -203.795 152.085 -203.230 ;
        RECT 146.610 -204.470 146.840 -203.970 ;
        RECT 147.100 -204.615 147.330 -203.970 ;
        RECT 147.590 -204.470 147.820 -203.970 ;
        RECT 148.080 -204.615 148.310 -203.970 ;
        RECT 146.610 -204.845 149.795 -204.615 ;
        RECT 146.610 -205.625 146.840 -204.845 ;
        RECT 147.100 -204.855 148.310 -204.845 ;
        RECT 147.590 -205.625 147.820 -204.855 ;
        RECT 148.570 -205.625 148.800 -204.845 ;
        RECT 138.570 -210.120 138.800 -208.620 ;
        RECT 136.805 -211.095 137.790 -210.825 ;
        RECT 138.080 -212.800 138.310 -211.305 ;
        RECT 138.075 -212.985 138.310 -212.800 ;
        RECT 138.570 -212.805 138.800 -211.305 ;
        RECT 139.060 -212.985 139.290 -211.305 ;
        RECT 139.550 -212.805 139.780 -208.620 ;
        RECT 141.615 -209.395 141.845 -208.615 ;
        RECT 142.595 -209.385 142.825 -208.615 ;
        RECT 142.105 -209.395 143.315 -209.385 ;
        RECT 143.575 -209.395 143.805 -208.615 ;
        RECT 141.615 -209.625 144.800 -209.395 ;
        RECT 141.615 -210.270 141.845 -209.770 ;
        RECT 142.105 -210.270 142.335 -209.625 ;
        RECT 142.595 -210.270 142.825 -209.770 ;
        RECT 143.085 -210.270 143.315 -209.625 ;
        RECT 145.805 -211.175 146.035 -208.175 ;
        RECT 146.860 -211.175 147.090 -208.175 ;
        RECT 147.350 -211.175 147.580 -208.175 ;
        RECT 147.840 -211.175 148.070 -208.175 ;
        RECT 148.900 -211.175 149.130 -208.175 ;
        RECT 140.040 -212.985 140.270 -211.305 ;
        RECT 150.055 -211.830 150.580 -211.470 ;
        RECT 150.085 -212.245 150.410 -211.830 ;
        RECT 145.310 -212.570 150.410 -212.245 ;
        RECT 138.075 -213.220 140.270 -212.985 ;
        RECT 145.805 -214.235 146.035 -212.735 ;
        RECT 146.295 -214.235 146.525 -212.735 ;
        RECT 146.785 -214.235 147.015 -212.735 ;
        RECT 147.995 -214.235 148.225 -212.735 ;
        RECT 148.485 -214.235 148.715 -212.735 ;
        RECT 151.520 -214.775 152.085 -203.795 ;
        RECT 155.610 -203.960 156.260 -203.210 ;
        RECT 157.040 -203.480 157.270 -202.480 ;
        RECT 157.530 -203.620 157.760 -202.480 ;
        RECT 158.020 -203.480 158.250 -202.480 ;
        RECT 158.510 -203.620 158.740 -202.480 ;
        RECT 159.695 -203.210 159.965 -201.760 ;
        RECT 161.415 -203.090 161.645 -201.595 ;
        RECT 161.905 -203.090 162.135 -201.590 ;
        RECT 162.395 -203.090 162.625 -201.410 ;
        RECT 159.695 -203.480 161.335 -203.210 ;
        RECT 157.040 -203.850 160.225 -203.620 ;
        RECT 161.065 -203.755 161.335 -203.480 ;
        RECT 155.860 -210.980 156.130 -203.960 ;
        RECT 157.040 -205.130 157.270 -203.850 ;
        RECT 157.530 -203.860 158.740 -203.850 ;
        RECT 158.020 -205.130 158.250 -203.860 ;
        RECT 159.000 -205.130 159.230 -203.850 ;
        RECT 160.935 -204.045 161.730 -203.755 ;
        RECT 161.905 -205.775 162.135 -204.275 ;
        RECT 162.885 -205.775 163.115 -201.590 ;
        RECT 163.375 -203.090 163.605 -201.410 ;
        RECT 166.885 -203.950 170.425 -203.385 ;
        RECT 164.950 -204.625 165.180 -204.125 ;
        RECT 165.440 -204.770 165.670 -204.125 ;
        RECT 165.930 -204.625 166.160 -204.125 ;
        RECT 166.420 -204.770 166.650 -204.125 ;
        RECT 164.950 -205.000 168.135 -204.770 ;
        RECT 164.950 -205.780 165.180 -205.000 ;
        RECT 165.440 -205.010 166.650 -205.000 ;
        RECT 165.930 -205.780 166.160 -205.010 ;
        RECT 166.910 -205.780 167.140 -205.000 ;
        RECT 156.910 -210.275 157.140 -208.775 ;
        RECT 155.145 -211.250 156.130 -210.980 ;
        RECT 156.420 -212.955 156.650 -211.460 ;
        RECT 156.415 -213.140 156.650 -212.955 ;
        RECT 156.910 -212.960 157.140 -211.460 ;
        RECT 157.400 -213.140 157.630 -211.460 ;
        RECT 157.890 -212.960 158.120 -208.775 ;
        RECT 159.955 -209.550 160.185 -208.770 ;
        RECT 160.935 -209.540 161.165 -208.770 ;
        RECT 160.445 -209.550 161.655 -209.540 ;
        RECT 161.915 -209.550 162.145 -208.770 ;
        RECT 159.955 -209.780 163.140 -209.550 ;
        RECT 159.955 -210.425 160.185 -209.925 ;
        RECT 160.445 -210.425 160.675 -209.780 ;
        RECT 160.935 -210.425 161.165 -209.925 ;
        RECT 161.425 -210.425 161.655 -209.780 ;
        RECT 164.145 -211.330 164.375 -208.330 ;
        RECT 165.200 -211.330 165.430 -208.330 ;
        RECT 165.690 -211.330 165.920 -208.330 ;
        RECT 166.180 -211.330 166.410 -208.330 ;
        RECT 167.240 -211.330 167.470 -208.330 ;
        RECT 158.380 -213.140 158.610 -211.460 ;
        RECT 168.395 -211.985 168.920 -211.625 ;
        RECT 168.425 -212.400 168.750 -211.985 ;
        RECT 163.650 -212.725 168.750 -212.400 ;
        RECT 156.415 -213.375 158.610 -213.140 ;
        RECT 164.145 -214.390 164.375 -212.890 ;
        RECT 164.635 -214.390 164.865 -212.890 ;
        RECT 165.125 -214.390 165.355 -212.890 ;
        RECT 166.335 -214.390 166.565 -212.890 ;
        RECT 166.825 -214.390 167.055 -212.890 ;
        RECT 148.700 -214.930 152.085 -214.775 ;
        RECT 169.860 -214.930 170.425 -203.950 ;
        RECT 170.845 -212.055 172.090 -184.610 ;
        RECT 172.900 -200.975 173.855 -182.405 ;
        RECT 176.280 -184.125 178.065 -183.445 ;
        RECT 185.310 -184.045 187.505 -183.810 ;
        RECT 176.280 -184.395 183.865 -184.125 ;
        RECT 185.310 -184.230 185.545 -184.045 ;
        RECT 176.280 -184.780 178.065 -184.395 ;
        RECT 179.510 -186.595 180.160 -185.845 ;
        RECT 180.940 -186.115 181.170 -185.115 ;
        RECT 181.430 -186.255 181.660 -185.115 ;
        RECT 181.920 -186.115 182.150 -185.115 ;
        RECT 182.410 -186.255 182.640 -185.115 ;
        RECT 183.595 -185.845 183.865 -184.395 ;
        RECT 185.315 -185.725 185.545 -184.230 ;
        RECT 185.805 -185.725 186.035 -184.225 ;
        RECT 186.295 -185.725 186.525 -184.045 ;
        RECT 183.595 -186.115 185.235 -185.845 ;
        RECT 180.940 -186.485 184.125 -186.255 ;
        RECT 184.965 -186.390 185.235 -186.115 ;
        RECT 179.760 -193.615 180.030 -186.595 ;
        RECT 180.940 -187.765 181.170 -186.485 ;
        RECT 181.430 -186.495 182.640 -186.485 ;
        RECT 181.920 -187.765 182.150 -186.495 ;
        RECT 182.900 -187.765 183.130 -186.485 ;
        RECT 184.835 -186.680 185.630 -186.390 ;
        RECT 185.805 -188.410 186.035 -186.910 ;
        RECT 186.785 -188.410 187.015 -184.225 ;
        RECT 187.275 -185.725 187.505 -184.045 ;
        RECT 190.785 -186.585 194.325 -186.020 ;
        RECT 188.850 -187.260 189.080 -186.760 ;
        RECT 189.340 -187.405 189.570 -186.760 ;
        RECT 189.830 -187.260 190.060 -186.760 ;
        RECT 190.320 -187.405 190.550 -186.760 ;
        RECT 188.850 -187.635 192.035 -187.405 ;
        RECT 188.850 -188.415 189.080 -187.635 ;
        RECT 189.340 -187.645 190.550 -187.635 ;
        RECT 189.830 -188.415 190.060 -187.645 ;
        RECT 190.810 -188.415 191.040 -187.635 ;
        RECT 180.810 -192.910 181.040 -191.410 ;
        RECT 179.045 -193.885 180.030 -193.615 ;
        RECT 180.320 -195.590 180.550 -194.095 ;
        RECT 180.315 -195.775 180.550 -195.590 ;
        RECT 180.810 -195.595 181.040 -194.095 ;
        RECT 181.300 -195.775 181.530 -194.095 ;
        RECT 181.790 -195.595 182.020 -191.410 ;
        RECT 183.855 -192.185 184.085 -191.405 ;
        RECT 184.835 -192.175 185.065 -191.405 ;
        RECT 184.345 -192.185 185.555 -192.175 ;
        RECT 185.815 -192.185 186.045 -191.405 ;
        RECT 183.855 -192.415 187.040 -192.185 ;
        RECT 183.855 -193.060 184.085 -192.560 ;
        RECT 184.345 -193.060 184.575 -192.415 ;
        RECT 184.835 -193.060 185.065 -192.560 ;
        RECT 185.325 -193.060 185.555 -192.415 ;
        RECT 188.045 -193.965 188.275 -190.965 ;
        RECT 189.100 -193.965 189.330 -190.965 ;
        RECT 189.590 -193.965 189.820 -190.965 ;
        RECT 190.080 -193.965 190.310 -190.965 ;
        RECT 191.140 -193.965 191.370 -190.965 ;
        RECT 182.280 -195.775 182.510 -194.095 ;
        RECT 192.295 -194.620 192.820 -194.260 ;
        RECT 192.325 -195.035 192.650 -194.620 ;
        RECT 187.550 -195.360 192.650 -195.035 ;
        RECT 180.315 -196.010 182.510 -195.775 ;
        RECT 188.045 -197.025 188.275 -195.525 ;
        RECT 188.535 -197.025 188.765 -195.525 ;
        RECT 189.025 -197.025 189.255 -195.525 ;
        RECT 190.235 -197.025 190.465 -195.525 ;
        RECT 190.725 -197.025 190.955 -195.525 ;
        RECT 191.890 -197.565 192.455 -197.560 ;
        RECT 193.760 -197.565 194.325 -186.585 ;
        RECT 198.005 -192.755 198.235 -190.255 ;
        RECT 199.350 -192.755 199.580 -190.255 ;
        RECT 199.840 -192.755 200.070 -190.255 ;
        RECT 200.330 -192.755 200.560 -190.255 ;
        RECT 200.980 -192.755 201.210 -190.255 ;
        RECT 202.610 -192.755 202.840 -190.255 ;
        RECT 203.750 -191.755 203.980 -190.255 ;
        RECT 196.850 -193.555 197.540 -193.535 ;
        RECT 200.880 -193.555 201.570 -193.535 ;
        RECT 202.805 -193.555 203.075 -193.190 ;
        RECT 196.850 -193.775 203.075 -193.555 ;
        RECT 196.850 -193.805 197.540 -193.775 ;
        RECT 200.880 -193.805 201.570 -193.775 ;
        RECT 202.805 -193.880 203.075 -193.775 ;
        RECT 203.665 -193.955 203.995 -193.895 ;
        RECT 207.230 -193.955 208.310 -182.405 ;
        RECT 196.045 -195.490 196.560 -195.035 ;
        RECT 190.940 -198.130 194.325 -197.565 ;
        RECT 172.900 -201.390 177.150 -200.975 ;
        RECT 185.270 -201.310 187.465 -201.075 ;
        RECT 172.900 -201.660 183.825 -201.390 ;
        RECT 185.270 -201.495 185.505 -201.310 ;
        RECT 172.900 -201.930 177.150 -201.660 ;
        RECT 179.470 -203.860 180.120 -203.110 ;
        RECT 180.900 -203.380 181.130 -202.380 ;
        RECT 181.390 -203.520 181.620 -202.380 ;
        RECT 181.880 -203.380 182.110 -202.380 ;
        RECT 182.370 -203.520 182.600 -202.380 ;
        RECT 183.555 -203.110 183.825 -201.660 ;
        RECT 185.275 -202.990 185.505 -201.495 ;
        RECT 185.765 -202.990 185.995 -201.490 ;
        RECT 186.255 -202.990 186.485 -201.310 ;
        RECT 183.555 -203.380 185.195 -203.110 ;
        RECT 180.900 -203.750 184.085 -203.520 ;
        RECT 184.925 -203.655 185.195 -203.380 ;
        RECT 179.720 -210.880 179.990 -203.860 ;
        RECT 180.900 -205.030 181.130 -203.750 ;
        RECT 181.390 -203.760 182.600 -203.750 ;
        RECT 181.880 -205.030 182.110 -203.760 ;
        RECT 182.860 -205.030 183.090 -203.750 ;
        RECT 184.795 -203.945 185.590 -203.655 ;
        RECT 185.765 -205.675 185.995 -204.175 ;
        RECT 186.745 -205.675 186.975 -201.490 ;
        RECT 187.235 -202.990 187.465 -201.310 ;
        RECT 191.890 -203.285 192.455 -198.130 ;
        RECT 196.105 -198.655 196.500 -195.490 ;
        RECT 197.515 -196.735 197.745 -195.235 ;
        RECT 198.005 -196.735 198.235 -195.235 ;
        RECT 199.865 -196.735 200.095 -194.235 ;
        RECT 200.355 -196.735 200.585 -194.235 ;
        RECT 200.980 -196.735 201.210 -194.235 ;
        RECT 201.470 -196.735 201.700 -194.235 ;
        RECT 202.120 -196.735 202.350 -194.235 ;
        RECT 202.610 -196.735 202.840 -194.235 ;
        RECT 203.100 -196.735 203.330 -194.235 ;
        RECT 203.665 -194.265 211.775 -193.955 ;
        RECT 203.665 -194.310 203.995 -194.265 ;
        RECT 203.750 -196.735 203.980 -195.235 ;
        RECT 204.240 -196.735 204.470 -195.235 ;
        RECT 193.605 -199.050 196.500 -198.655 ;
        RECT 193.605 -200.825 194.000 -199.050 ;
        RECT 193.475 -201.310 194.055 -200.825 ;
        RECT 203.610 -201.465 205.805 -201.230 ;
        RECT 196.620 -201.545 197.105 -201.515 ;
        RECT 196.620 -201.815 202.165 -201.545 ;
        RECT 203.610 -201.650 203.845 -201.465 ;
        RECT 196.620 -201.845 197.105 -201.815 ;
        RECT 190.745 -203.850 194.285 -203.285 ;
        RECT 188.810 -204.525 189.040 -204.025 ;
        RECT 189.300 -204.670 189.530 -204.025 ;
        RECT 189.790 -204.525 190.020 -204.025 ;
        RECT 190.280 -204.670 190.510 -204.025 ;
        RECT 188.810 -204.900 191.995 -204.670 ;
        RECT 188.810 -205.680 189.040 -204.900 ;
        RECT 189.300 -204.910 190.510 -204.900 ;
        RECT 189.790 -205.680 190.020 -204.910 ;
        RECT 190.770 -205.680 191.000 -204.900 ;
        RECT 180.770 -210.175 181.000 -208.675 ;
        RECT 179.005 -211.150 179.990 -210.880 ;
        RECT 170.925 -212.900 172.040 -212.055 ;
        RECT 180.280 -212.855 180.510 -211.360 ;
        RECT 180.275 -213.040 180.510 -212.855 ;
        RECT 180.770 -212.860 181.000 -211.360 ;
        RECT 181.260 -213.040 181.490 -211.360 ;
        RECT 181.750 -212.860 181.980 -208.675 ;
        RECT 183.815 -209.450 184.045 -208.670 ;
        RECT 184.795 -209.440 185.025 -208.670 ;
        RECT 184.305 -209.450 185.515 -209.440 ;
        RECT 185.775 -209.450 186.005 -208.670 ;
        RECT 183.815 -209.680 187.000 -209.450 ;
        RECT 183.815 -210.325 184.045 -209.825 ;
        RECT 184.305 -210.325 184.535 -209.680 ;
        RECT 184.795 -210.325 185.025 -209.825 ;
        RECT 185.285 -210.325 185.515 -209.680 ;
        RECT 188.005 -211.230 188.235 -208.230 ;
        RECT 189.060 -211.230 189.290 -208.230 ;
        RECT 189.550 -211.230 189.780 -208.230 ;
        RECT 190.040 -211.230 190.270 -208.230 ;
        RECT 191.100 -211.230 191.330 -208.230 ;
        RECT 182.240 -213.040 182.470 -211.360 ;
        RECT 192.255 -211.885 192.780 -211.525 ;
        RECT 192.285 -212.300 192.610 -211.885 ;
        RECT 187.510 -212.625 192.610 -212.300 ;
        RECT 180.275 -213.275 182.470 -213.040 ;
        RECT 188.005 -214.290 188.235 -212.790 ;
        RECT 188.495 -214.290 188.725 -212.790 ;
        RECT 188.985 -214.290 189.215 -212.790 ;
        RECT 190.195 -214.290 190.425 -212.790 ;
        RECT 190.685 -214.290 190.915 -212.790 ;
        RECT 193.720 -214.830 194.285 -203.850 ;
        RECT 197.810 -204.015 198.460 -203.265 ;
        RECT 199.240 -203.535 199.470 -202.535 ;
        RECT 199.730 -203.675 199.960 -202.535 ;
        RECT 200.220 -203.535 200.450 -202.535 ;
        RECT 200.710 -203.675 200.940 -202.535 ;
        RECT 201.895 -203.265 202.165 -201.815 ;
        RECT 203.615 -203.145 203.845 -201.650 ;
        RECT 204.105 -203.145 204.335 -201.645 ;
        RECT 204.595 -203.145 204.825 -201.465 ;
        RECT 201.895 -203.535 203.535 -203.265 ;
        RECT 199.240 -203.905 202.425 -203.675 ;
        RECT 203.265 -203.810 203.535 -203.535 ;
        RECT 198.060 -211.035 198.330 -204.015 ;
        RECT 199.240 -205.185 199.470 -203.905 ;
        RECT 199.730 -203.915 200.940 -203.905 ;
        RECT 200.220 -205.185 200.450 -203.915 ;
        RECT 201.200 -205.185 201.430 -203.905 ;
        RECT 203.135 -204.100 203.930 -203.810 ;
        RECT 204.105 -205.830 204.335 -204.330 ;
        RECT 205.085 -205.830 205.315 -201.645 ;
        RECT 205.575 -203.145 205.805 -201.465 ;
        RECT 209.085 -204.005 212.625 -203.440 ;
        RECT 207.150 -204.680 207.380 -204.180 ;
        RECT 207.640 -204.825 207.870 -204.180 ;
        RECT 208.130 -204.680 208.360 -204.180 ;
        RECT 208.620 -204.825 208.850 -204.180 ;
        RECT 207.150 -205.055 210.335 -204.825 ;
        RECT 207.150 -205.835 207.380 -205.055 ;
        RECT 207.640 -205.065 208.850 -205.055 ;
        RECT 208.130 -205.835 208.360 -205.065 ;
        RECT 209.110 -205.835 209.340 -205.055 ;
        RECT 199.110 -210.330 199.340 -208.830 ;
        RECT 197.345 -211.305 198.330 -211.035 ;
        RECT 198.620 -213.010 198.850 -211.515 ;
        RECT 198.615 -213.195 198.850 -213.010 ;
        RECT 199.110 -213.015 199.340 -211.515 ;
        RECT 199.600 -213.195 199.830 -211.515 ;
        RECT 200.090 -213.015 200.320 -208.830 ;
        RECT 202.155 -209.605 202.385 -208.825 ;
        RECT 203.135 -209.595 203.365 -208.825 ;
        RECT 202.645 -209.605 203.855 -209.595 ;
        RECT 204.115 -209.605 204.345 -208.825 ;
        RECT 202.155 -209.835 205.340 -209.605 ;
        RECT 202.155 -210.480 202.385 -209.980 ;
        RECT 202.645 -210.480 202.875 -209.835 ;
        RECT 203.135 -210.480 203.365 -209.980 ;
        RECT 203.625 -210.480 203.855 -209.835 ;
        RECT 206.345 -211.385 206.575 -208.385 ;
        RECT 207.400 -211.385 207.630 -208.385 ;
        RECT 207.890 -211.385 208.120 -208.385 ;
        RECT 208.380 -211.385 208.610 -208.385 ;
        RECT 209.440 -211.385 209.670 -208.385 ;
        RECT 200.580 -213.195 200.810 -211.515 ;
        RECT 210.595 -212.040 211.120 -211.680 ;
        RECT 210.625 -212.455 210.950 -212.040 ;
        RECT 205.850 -212.780 210.950 -212.455 ;
        RECT 198.615 -213.430 200.810 -213.195 ;
        RECT 206.345 -214.445 206.575 -212.945 ;
        RECT 206.835 -214.445 207.065 -212.945 ;
        RECT 207.325 -214.445 207.555 -212.945 ;
        RECT 208.535 -214.445 208.765 -212.945 ;
        RECT 209.025 -214.445 209.255 -212.945 ;
        RECT 148.700 -215.340 170.425 -214.930 ;
        RECT 148.720 -215.495 170.425 -215.340 ;
        RECT 190.900 -214.985 194.285 -214.830 ;
        RECT 212.060 -214.985 212.625 -204.005 ;
        RECT 213.170 -211.740 214.495 -175.075 ;
        RECT 215.380 -182.370 255.185 -181.360 ;
        RECT 215.380 -201.320 216.390 -182.370 ;
        RECT 220.800 -184.320 222.285 -183.890 ;
        RECT 229.625 -184.240 231.820 -184.005 ;
        RECT 220.800 -184.590 228.180 -184.320 ;
        RECT 229.625 -184.425 229.860 -184.240 ;
        RECT 220.800 -185.000 222.285 -184.590 ;
        RECT 223.825 -186.790 224.475 -186.040 ;
        RECT 225.255 -186.310 225.485 -185.310 ;
        RECT 225.745 -186.450 225.975 -185.310 ;
        RECT 226.235 -186.310 226.465 -185.310 ;
        RECT 226.725 -186.450 226.955 -185.310 ;
        RECT 227.910 -186.040 228.180 -184.590 ;
        RECT 229.630 -185.920 229.860 -184.425 ;
        RECT 230.120 -185.920 230.350 -184.420 ;
        RECT 230.610 -185.920 230.840 -184.240 ;
        RECT 227.910 -186.310 229.550 -186.040 ;
        RECT 225.255 -186.680 228.440 -186.450 ;
        RECT 229.280 -186.585 229.550 -186.310 ;
        RECT 224.075 -193.810 224.345 -186.790 ;
        RECT 225.255 -187.960 225.485 -186.680 ;
        RECT 225.745 -186.690 226.955 -186.680 ;
        RECT 226.235 -187.960 226.465 -186.690 ;
        RECT 227.215 -187.960 227.445 -186.680 ;
        RECT 229.150 -186.875 229.945 -186.585 ;
        RECT 230.120 -188.605 230.350 -187.105 ;
        RECT 231.100 -188.605 231.330 -184.420 ;
        RECT 231.590 -185.920 231.820 -184.240 ;
        RECT 235.100 -186.780 238.640 -186.215 ;
        RECT 233.165 -187.455 233.395 -186.955 ;
        RECT 233.655 -187.600 233.885 -186.955 ;
        RECT 234.145 -187.455 234.375 -186.955 ;
        RECT 234.635 -187.600 234.865 -186.955 ;
        RECT 233.165 -187.830 236.350 -187.600 ;
        RECT 233.165 -188.610 233.395 -187.830 ;
        RECT 233.655 -187.840 234.865 -187.830 ;
        RECT 234.145 -188.610 234.375 -187.840 ;
        RECT 235.125 -188.610 235.355 -187.830 ;
        RECT 225.125 -193.105 225.355 -191.605 ;
        RECT 223.360 -194.080 224.345 -193.810 ;
        RECT 224.635 -195.785 224.865 -194.290 ;
        RECT 224.630 -195.970 224.865 -195.785 ;
        RECT 225.125 -195.790 225.355 -194.290 ;
        RECT 225.615 -195.970 225.845 -194.290 ;
        RECT 226.105 -195.790 226.335 -191.605 ;
        RECT 228.170 -192.380 228.400 -191.600 ;
        RECT 229.150 -192.370 229.380 -191.600 ;
        RECT 228.660 -192.380 229.870 -192.370 ;
        RECT 230.130 -192.380 230.360 -191.600 ;
        RECT 228.170 -192.610 231.355 -192.380 ;
        RECT 228.170 -193.255 228.400 -192.755 ;
        RECT 228.660 -193.255 228.890 -192.610 ;
        RECT 229.150 -193.255 229.380 -192.755 ;
        RECT 229.640 -193.255 229.870 -192.610 ;
        RECT 232.360 -194.160 232.590 -191.160 ;
        RECT 233.415 -194.160 233.645 -191.160 ;
        RECT 233.905 -194.160 234.135 -191.160 ;
        RECT 234.395 -194.160 234.625 -191.160 ;
        RECT 235.455 -194.160 235.685 -191.160 ;
        RECT 226.595 -195.970 226.825 -194.290 ;
        RECT 236.610 -194.815 237.135 -194.455 ;
        RECT 236.640 -195.230 236.965 -194.815 ;
        RECT 231.865 -195.555 236.965 -195.230 ;
        RECT 224.630 -196.205 226.825 -195.970 ;
        RECT 232.360 -197.220 232.590 -195.720 ;
        RECT 232.850 -197.220 233.080 -195.720 ;
        RECT 233.340 -197.220 233.570 -195.720 ;
        RECT 234.550 -197.220 234.780 -195.720 ;
        RECT 235.040 -197.220 235.270 -195.720 ;
        RECT 236.205 -197.760 236.770 -197.755 ;
        RECT 238.075 -197.760 238.640 -186.780 ;
        RECT 242.320 -192.950 242.550 -190.450 ;
        RECT 243.665 -192.950 243.895 -190.450 ;
        RECT 244.155 -192.950 244.385 -190.450 ;
        RECT 244.645 -192.950 244.875 -190.450 ;
        RECT 245.295 -192.950 245.525 -190.450 ;
        RECT 246.925 -192.950 247.155 -190.450 ;
        RECT 248.065 -191.950 248.295 -190.450 ;
        RECT 241.165 -193.750 241.855 -193.730 ;
        RECT 245.195 -193.750 245.885 -193.730 ;
        RECT 247.120 -193.750 247.390 -193.385 ;
        RECT 241.165 -193.970 247.390 -193.750 ;
        RECT 241.165 -194.000 241.855 -193.970 ;
        RECT 245.195 -194.000 245.885 -193.970 ;
        RECT 247.120 -194.075 247.390 -193.970 ;
        RECT 247.980 -194.150 248.310 -194.090 ;
        RECT 254.175 -194.150 255.185 -182.370 ;
        RECT 240.360 -195.685 240.875 -195.230 ;
        RECT 235.255 -198.325 238.640 -197.760 ;
        RECT 215.380 -201.585 222.030 -201.320 ;
        RECT 229.585 -201.505 231.780 -201.270 ;
        RECT 215.380 -201.855 228.140 -201.585 ;
        RECT 229.585 -201.690 229.820 -201.505 ;
        RECT 215.380 -202.330 222.030 -201.855 ;
        RECT 223.785 -204.055 224.435 -203.305 ;
        RECT 225.215 -203.575 225.445 -202.575 ;
        RECT 225.705 -203.715 225.935 -202.575 ;
        RECT 226.195 -203.575 226.425 -202.575 ;
        RECT 226.685 -203.715 226.915 -202.575 ;
        RECT 227.870 -203.305 228.140 -201.855 ;
        RECT 229.590 -203.185 229.820 -201.690 ;
        RECT 230.080 -203.185 230.310 -201.685 ;
        RECT 230.570 -203.185 230.800 -201.505 ;
        RECT 227.870 -203.575 229.510 -203.305 ;
        RECT 225.215 -203.945 228.400 -203.715 ;
        RECT 229.240 -203.850 229.510 -203.575 ;
        RECT 224.035 -211.075 224.305 -204.055 ;
        RECT 225.215 -205.225 225.445 -203.945 ;
        RECT 225.705 -203.955 226.915 -203.945 ;
        RECT 226.195 -205.225 226.425 -203.955 ;
        RECT 227.175 -205.225 227.405 -203.945 ;
        RECT 229.110 -204.140 229.905 -203.850 ;
        RECT 230.080 -205.870 230.310 -204.370 ;
        RECT 231.060 -205.870 231.290 -201.685 ;
        RECT 231.550 -203.185 231.780 -201.505 ;
        RECT 236.205 -203.480 236.770 -198.325 ;
        RECT 240.420 -198.850 240.815 -195.685 ;
        RECT 241.830 -196.930 242.060 -195.430 ;
        RECT 242.320 -196.930 242.550 -195.430 ;
        RECT 244.180 -196.930 244.410 -194.430 ;
        RECT 244.670 -196.930 244.900 -194.430 ;
        RECT 245.295 -196.930 245.525 -194.430 ;
        RECT 245.785 -196.930 246.015 -194.430 ;
        RECT 246.435 -196.930 246.665 -194.430 ;
        RECT 246.925 -196.930 247.155 -194.430 ;
        RECT 247.415 -196.930 247.645 -194.430 ;
        RECT 247.980 -194.460 256.090 -194.150 ;
        RECT 247.980 -194.505 248.310 -194.460 ;
        RECT 248.065 -196.930 248.295 -195.430 ;
        RECT 248.555 -196.930 248.785 -195.430 ;
        RECT 237.920 -199.245 240.815 -198.850 ;
        RECT 237.920 -201.020 238.315 -199.245 ;
        RECT 237.790 -201.505 238.370 -201.020 ;
        RECT 247.925 -201.660 250.120 -201.425 ;
        RECT 240.935 -201.740 241.420 -201.710 ;
        RECT 240.935 -202.010 246.480 -201.740 ;
        RECT 247.925 -201.845 248.160 -201.660 ;
        RECT 240.935 -202.040 241.420 -202.010 ;
        RECT 235.060 -204.045 238.600 -203.480 ;
        RECT 233.125 -204.720 233.355 -204.220 ;
        RECT 233.615 -204.865 233.845 -204.220 ;
        RECT 234.105 -204.720 234.335 -204.220 ;
        RECT 234.595 -204.865 234.825 -204.220 ;
        RECT 233.125 -205.095 236.310 -204.865 ;
        RECT 233.125 -205.875 233.355 -205.095 ;
        RECT 233.615 -205.105 234.825 -205.095 ;
        RECT 234.105 -205.875 234.335 -205.105 ;
        RECT 235.085 -205.875 235.315 -205.095 ;
        RECT 225.085 -210.370 225.315 -208.870 ;
        RECT 223.320 -211.345 224.305 -211.075 ;
        RECT 213.170 -213.395 214.855 -211.740 ;
        RECT 224.595 -213.050 224.825 -211.555 ;
        RECT 224.590 -213.235 224.825 -213.050 ;
        RECT 225.085 -213.055 225.315 -211.555 ;
        RECT 225.575 -213.235 225.805 -211.555 ;
        RECT 226.065 -213.055 226.295 -208.870 ;
        RECT 228.130 -209.645 228.360 -208.865 ;
        RECT 229.110 -209.635 229.340 -208.865 ;
        RECT 228.620 -209.645 229.830 -209.635 ;
        RECT 230.090 -209.645 230.320 -208.865 ;
        RECT 228.130 -209.875 231.315 -209.645 ;
        RECT 228.130 -210.520 228.360 -210.020 ;
        RECT 228.620 -210.520 228.850 -209.875 ;
        RECT 229.110 -210.520 229.340 -210.020 ;
        RECT 229.600 -210.520 229.830 -209.875 ;
        RECT 232.320 -211.425 232.550 -208.425 ;
        RECT 233.375 -211.425 233.605 -208.425 ;
        RECT 233.865 -211.425 234.095 -208.425 ;
        RECT 234.355 -211.425 234.585 -208.425 ;
        RECT 235.415 -211.425 235.645 -208.425 ;
        RECT 226.555 -213.235 226.785 -211.555 ;
        RECT 236.570 -212.080 237.095 -211.720 ;
        RECT 236.600 -212.495 236.925 -212.080 ;
        RECT 231.825 -212.820 236.925 -212.495 ;
        RECT 224.590 -213.470 226.785 -213.235 ;
        RECT 232.320 -214.485 232.550 -212.985 ;
        RECT 232.810 -214.485 233.040 -212.985 ;
        RECT 233.300 -214.485 233.530 -212.985 ;
        RECT 234.510 -214.485 234.740 -212.985 ;
        RECT 235.000 -214.485 235.230 -212.985 ;
        RECT 190.900 -215.395 212.625 -214.985 ;
        RECT 238.035 -215.025 238.600 -204.045 ;
        RECT 242.125 -204.210 242.775 -203.460 ;
        RECT 243.555 -203.730 243.785 -202.730 ;
        RECT 244.045 -203.870 244.275 -202.730 ;
        RECT 244.535 -203.730 244.765 -202.730 ;
        RECT 245.025 -203.870 245.255 -202.730 ;
        RECT 246.210 -203.460 246.480 -202.010 ;
        RECT 247.930 -203.340 248.160 -201.845 ;
        RECT 248.420 -203.340 248.650 -201.840 ;
        RECT 248.910 -203.340 249.140 -201.660 ;
        RECT 246.210 -203.730 247.850 -203.460 ;
        RECT 243.555 -204.100 246.740 -203.870 ;
        RECT 247.580 -204.005 247.850 -203.730 ;
        RECT 242.375 -211.230 242.645 -204.210 ;
        RECT 243.555 -205.380 243.785 -204.100 ;
        RECT 244.045 -204.110 245.255 -204.100 ;
        RECT 244.535 -205.380 244.765 -204.110 ;
        RECT 245.515 -205.380 245.745 -204.100 ;
        RECT 247.450 -204.295 248.245 -204.005 ;
        RECT 248.420 -206.025 248.650 -204.525 ;
        RECT 249.400 -206.025 249.630 -201.840 ;
        RECT 249.890 -203.340 250.120 -201.660 ;
        RECT 253.400 -204.200 256.940 -203.635 ;
        RECT 251.465 -204.875 251.695 -204.375 ;
        RECT 251.955 -205.020 252.185 -204.375 ;
        RECT 252.445 -204.875 252.675 -204.375 ;
        RECT 252.935 -205.020 253.165 -204.375 ;
        RECT 251.465 -205.250 254.650 -205.020 ;
        RECT 251.465 -206.030 251.695 -205.250 ;
        RECT 251.955 -205.260 253.165 -205.250 ;
        RECT 252.445 -206.030 252.675 -205.260 ;
        RECT 253.425 -206.030 253.655 -205.250 ;
        RECT 243.425 -210.525 243.655 -209.025 ;
        RECT 241.660 -211.500 242.645 -211.230 ;
        RECT 242.935 -213.205 243.165 -211.710 ;
        RECT 242.930 -213.390 243.165 -213.205 ;
        RECT 243.425 -213.210 243.655 -211.710 ;
        RECT 243.915 -213.390 244.145 -211.710 ;
        RECT 244.405 -213.210 244.635 -209.025 ;
        RECT 246.470 -209.800 246.700 -209.020 ;
        RECT 247.450 -209.790 247.680 -209.020 ;
        RECT 246.960 -209.800 248.170 -209.790 ;
        RECT 248.430 -209.800 248.660 -209.020 ;
        RECT 246.470 -210.030 249.655 -209.800 ;
        RECT 246.470 -210.675 246.700 -210.175 ;
        RECT 246.960 -210.675 247.190 -210.030 ;
        RECT 247.450 -210.675 247.680 -210.175 ;
        RECT 247.940 -210.675 248.170 -210.030 ;
        RECT 250.660 -211.580 250.890 -208.580 ;
        RECT 251.715 -211.580 251.945 -208.580 ;
        RECT 252.205 -211.580 252.435 -208.580 ;
        RECT 252.695 -211.580 252.925 -208.580 ;
        RECT 253.755 -211.580 253.985 -208.580 ;
        RECT 244.895 -213.390 245.125 -211.710 ;
        RECT 254.910 -212.235 255.435 -211.875 ;
        RECT 254.940 -212.650 255.265 -212.235 ;
        RECT 250.165 -212.975 255.265 -212.650 ;
        RECT 242.930 -213.625 245.125 -213.390 ;
        RECT 250.660 -214.640 250.890 -213.140 ;
        RECT 251.150 -214.640 251.380 -213.140 ;
        RECT 251.640 -214.640 251.870 -213.140 ;
        RECT 252.850 -214.640 253.080 -213.140 ;
        RECT 253.340 -214.640 253.570 -213.140 ;
        RECT 190.920 -215.550 212.625 -215.395 ;
        RECT 235.215 -215.180 238.600 -215.025 ;
        RECT 256.375 -215.180 256.940 -204.200 ;
        RECT 257.490 -211.045 258.620 -172.675 ;
        RECT 261.775 -182.695 301.705 -181.400 ;
        RECT 261.775 -200.715 263.070 -182.695 ;
        RECT 265.755 -184.150 266.985 -183.670 ;
        RECT 275.615 -184.070 277.810 -183.835 ;
        RECT 265.755 -184.420 274.170 -184.150 ;
        RECT 275.615 -184.255 275.850 -184.070 ;
        RECT 265.755 -184.770 266.985 -184.420 ;
        RECT 269.815 -186.620 270.465 -185.870 ;
        RECT 271.245 -186.140 271.475 -185.140 ;
        RECT 271.735 -186.280 271.965 -185.140 ;
        RECT 272.225 -186.140 272.455 -185.140 ;
        RECT 272.715 -186.280 272.945 -185.140 ;
        RECT 273.900 -185.870 274.170 -184.420 ;
        RECT 275.620 -185.750 275.850 -184.255 ;
        RECT 276.110 -185.750 276.340 -184.250 ;
        RECT 276.600 -185.750 276.830 -184.070 ;
        RECT 273.900 -186.140 275.540 -185.870 ;
        RECT 271.245 -186.510 274.430 -186.280 ;
        RECT 275.270 -186.415 275.540 -186.140 ;
        RECT 270.065 -193.640 270.335 -186.620 ;
        RECT 271.245 -187.790 271.475 -186.510 ;
        RECT 271.735 -186.520 272.945 -186.510 ;
        RECT 272.225 -187.790 272.455 -186.520 ;
        RECT 273.205 -187.790 273.435 -186.510 ;
        RECT 275.140 -186.705 275.935 -186.415 ;
        RECT 276.110 -188.435 276.340 -186.935 ;
        RECT 277.090 -188.435 277.320 -184.250 ;
        RECT 277.580 -185.750 277.810 -184.070 ;
        RECT 281.090 -186.610 284.630 -186.045 ;
        RECT 279.155 -187.285 279.385 -186.785 ;
        RECT 279.645 -187.430 279.875 -186.785 ;
        RECT 280.135 -187.285 280.365 -186.785 ;
        RECT 280.625 -187.430 280.855 -186.785 ;
        RECT 279.155 -187.660 282.340 -187.430 ;
        RECT 279.155 -188.440 279.385 -187.660 ;
        RECT 279.645 -187.670 280.855 -187.660 ;
        RECT 280.135 -188.440 280.365 -187.670 ;
        RECT 281.115 -188.440 281.345 -187.660 ;
        RECT 271.115 -192.935 271.345 -191.435 ;
        RECT 269.350 -193.910 270.335 -193.640 ;
        RECT 270.625 -195.615 270.855 -194.120 ;
        RECT 270.620 -195.800 270.855 -195.615 ;
        RECT 271.115 -195.620 271.345 -194.120 ;
        RECT 271.605 -195.800 271.835 -194.120 ;
        RECT 272.095 -195.620 272.325 -191.435 ;
        RECT 274.160 -192.210 274.390 -191.430 ;
        RECT 275.140 -192.200 275.370 -191.430 ;
        RECT 274.650 -192.210 275.860 -192.200 ;
        RECT 276.120 -192.210 276.350 -191.430 ;
        RECT 274.160 -192.440 277.345 -192.210 ;
        RECT 274.160 -193.085 274.390 -192.585 ;
        RECT 274.650 -193.085 274.880 -192.440 ;
        RECT 275.140 -193.085 275.370 -192.585 ;
        RECT 275.630 -193.085 275.860 -192.440 ;
        RECT 278.350 -193.990 278.580 -190.990 ;
        RECT 279.405 -193.990 279.635 -190.990 ;
        RECT 279.895 -193.990 280.125 -190.990 ;
        RECT 280.385 -193.990 280.615 -190.990 ;
        RECT 281.445 -193.990 281.675 -190.990 ;
        RECT 272.585 -195.800 272.815 -194.120 ;
        RECT 282.600 -194.645 283.125 -194.285 ;
        RECT 282.630 -195.060 282.955 -194.645 ;
        RECT 277.855 -195.385 282.955 -195.060 ;
        RECT 270.620 -196.035 272.815 -195.800 ;
        RECT 278.350 -197.050 278.580 -195.550 ;
        RECT 278.840 -197.050 279.070 -195.550 ;
        RECT 279.330 -197.050 279.560 -195.550 ;
        RECT 280.540 -197.050 280.770 -195.550 ;
        RECT 281.030 -197.050 281.260 -195.550 ;
        RECT 282.195 -197.590 282.760 -197.585 ;
        RECT 284.065 -197.590 284.630 -186.610 ;
        RECT 288.310 -192.780 288.540 -190.280 ;
        RECT 289.655 -192.780 289.885 -190.280 ;
        RECT 290.145 -192.780 290.375 -190.280 ;
        RECT 290.635 -192.780 290.865 -190.280 ;
        RECT 291.285 -192.780 291.515 -190.280 ;
        RECT 292.915 -192.780 293.145 -190.280 ;
        RECT 294.055 -191.780 294.285 -190.280 ;
        RECT 287.155 -193.580 287.845 -193.560 ;
        RECT 291.185 -193.580 291.875 -193.560 ;
        RECT 293.110 -193.580 293.380 -193.215 ;
        RECT 287.155 -193.800 293.380 -193.580 ;
        RECT 287.155 -193.830 287.845 -193.800 ;
        RECT 291.185 -193.830 291.875 -193.800 ;
        RECT 293.110 -193.905 293.380 -193.800 ;
        RECT 293.970 -193.980 294.300 -193.920 ;
        RECT 300.410 -193.980 301.705 -182.695 ;
        RECT 303.460 -182.980 304.565 -169.890 ;
        RECT 305.720 -182.795 345.640 -181.605 ;
        RECT 302.945 -184.550 304.825 -182.980 ;
        RECT 286.350 -195.515 286.865 -195.060 ;
        RECT 281.245 -198.155 284.630 -197.590 ;
        RECT 261.775 -201.415 267.815 -200.715 ;
        RECT 275.575 -201.335 277.770 -201.100 ;
        RECT 261.775 -201.685 274.130 -201.415 ;
        RECT 275.575 -201.520 275.810 -201.335 ;
        RECT 261.775 -202.010 267.815 -201.685 ;
        RECT 269.775 -203.885 270.425 -203.135 ;
        RECT 271.205 -203.405 271.435 -202.405 ;
        RECT 271.695 -203.545 271.925 -202.405 ;
        RECT 272.185 -203.405 272.415 -202.405 ;
        RECT 272.675 -203.545 272.905 -202.405 ;
        RECT 273.860 -203.135 274.130 -201.685 ;
        RECT 275.580 -203.015 275.810 -201.520 ;
        RECT 276.070 -203.015 276.300 -201.515 ;
        RECT 276.560 -203.015 276.790 -201.335 ;
        RECT 273.860 -203.405 275.500 -203.135 ;
        RECT 271.205 -203.775 274.390 -203.545 ;
        RECT 275.230 -203.680 275.500 -203.405 ;
        RECT 270.025 -210.905 270.295 -203.885 ;
        RECT 271.205 -205.055 271.435 -203.775 ;
        RECT 271.695 -203.785 272.905 -203.775 ;
        RECT 272.185 -205.055 272.415 -203.785 ;
        RECT 273.165 -205.055 273.395 -203.775 ;
        RECT 275.100 -203.970 275.895 -203.680 ;
        RECT 276.070 -205.700 276.300 -204.200 ;
        RECT 277.050 -205.700 277.280 -201.515 ;
        RECT 277.540 -203.015 277.770 -201.335 ;
        RECT 282.195 -203.310 282.760 -198.155 ;
        RECT 286.410 -198.680 286.805 -195.515 ;
        RECT 287.820 -196.760 288.050 -195.260 ;
        RECT 288.310 -196.760 288.540 -195.260 ;
        RECT 290.170 -196.760 290.400 -194.260 ;
        RECT 290.660 -196.760 290.890 -194.260 ;
        RECT 291.285 -196.760 291.515 -194.260 ;
        RECT 291.775 -196.760 292.005 -194.260 ;
        RECT 292.425 -196.760 292.655 -194.260 ;
        RECT 292.915 -196.760 293.145 -194.260 ;
        RECT 293.405 -196.760 293.635 -194.260 ;
        RECT 293.970 -194.290 302.080 -193.980 ;
        RECT 293.970 -194.335 294.300 -194.290 ;
        RECT 294.055 -196.760 294.285 -195.260 ;
        RECT 294.545 -196.760 294.775 -195.260 ;
        RECT 283.910 -199.075 286.805 -198.680 ;
        RECT 283.910 -200.850 284.305 -199.075 ;
        RECT 283.780 -201.335 284.360 -200.850 ;
        RECT 293.915 -201.490 296.110 -201.255 ;
        RECT 286.925 -201.570 287.410 -201.540 ;
        RECT 286.925 -201.840 292.470 -201.570 ;
        RECT 293.915 -201.675 294.150 -201.490 ;
        RECT 286.925 -201.870 287.410 -201.840 ;
        RECT 281.050 -203.875 284.590 -203.310 ;
        RECT 279.115 -204.550 279.345 -204.050 ;
        RECT 279.605 -204.695 279.835 -204.050 ;
        RECT 280.095 -204.550 280.325 -204.050 ;
        RECT 280.585 -204.695 280.815 -204.050 ;
        RECT 279.115 -204.925 282.300 -204.695 ;
        RECT 279.115 -205.705 279.345 -204.925 ;
        RECT 279.605 -204.935 280.815 -204.925 ;
        RECT 280.095 -205.705 280.325 -204.935 ;
        RECT 281.075 -205.705 281.305 -204.925 ;
        RECT 271.075 -210.200 271.305 -208.700 ;
        RECT 257.380 -213.545 258.870 -211.045 ;
        RECT 269.310 -211.175 270.295 -210.905 ;
        RECT 270.585 -212.880 270.815 -211.385 ;
        RECT 270.580 -213.065 270.815 -212.880 ;
        RECT 271.075 -212.885 271.305 -211.385 ;
        RECT 271.565 -213.065 271.795 -211.385 ;
        RECT 272.055 -212.885 272.285 -208.700 ;
        RECT 274.120 -209.475 274.350 -208.695 ;
        RECT 275.100 -209.465 275.330 -208.695 ;
        RECT 274.610 -209.475 275.820 -209.465 ;
        RECT 276.080 -209.475 276.310 -208.695 ;
        RECT 274.120 -209.705 277.305 -209.475 ;
        RECT 274.120 -210.350 274.350 -209.850 ;
        RECT 274.610 -210.350 274.840 -209.705 ;
        RECT 275.100 -210.350 275.330 -209.850 ;
        RECT 275.590 -210.350 275.820 -209.705 ;
        RECT 278.310 -211.255 278.540 -208.255 ;
        RECT 279.365 -211.255 279.595 -208.255 ;
        RECT 279.855 -211.255 280.085 -208.255 ;
        RECT 280.345 -211.255 280.575 -208.255 ;
        RECT 281.405 -211.255 281.635 -208.255 ;
        RECT 272.545 -213.065 272.775 -211.385 ;
        RECT 282.560 -211.910 283.085 -211.550 ;
        RECT 282.590 -212.325 282.915 -211.910 ;
        RECT 277.815 -212.650 282.915 -212.325 ;
        RECT 270.580 -213.300 272.775 -213.065 ;
        RECT 278.310 -214.315 278.540 -212.815 ;
        RECT 278.800 -214.315 279.030 -212.815 ;
        RECT 279.290 -214.315 279.520 -212.815 ;
        RECT 280.500 -214.315 280.730 -212.815 ;
        RECT 280.990 -214.315 281.220 -212.815 ;
        RECT 284.025 -214.855 284.590 -203.875 ;
        RECT 288.115 -204.040 288.765 -203.290 ;
        RECT 289.545 -203.560 289.775 -202.560 ;
        RECT 290.035 -203.700 290.265 -202.560 ;
        RECT 290.525 -203.560 290.755 -202.560 ;
        RECT 291.015 -203.700 291.245 -202.560 ;
        RECT 292.200 -203.290 292.470 -201.840 ;
        RECT 293.920 -203.170 294.150 -201.675 ;
        RECT 294.410 -203.170 294.640 -201.670 ;
        RECT 294.900 -203.170 295.130 -201.490 ;
        RECT 292.200 -203.560 293.840 -203.290 ;
        RECT 289.545 -203.930 292.730 -203.700 ;
        RECT 293.570 -203.835 293.840 -203.560 ;
        RECT 288.365 -211.060 288.635 -204.040 ;
        RECT 289.545 -205.210 289.775 -203.930 ;
        RECT 290.035 -203.940 291.245 -203.930 ;
        RECT 290.525 -205.210 290.755 -203.940 ;
        RECT 291.505 -205.210 291.735 -203.930 ;
        RECT 293.440 -204.125 294.235 -203.835 ;
        RECT 294.410 -205.855 294.640 -204.355 ;
        RECT 295.390 -205.855 295.620 -201.670 ;
        RECT 295.880 -203.170 296.110 -201.490 ;
        RECT 299.390 -204.030 302.930 -203.465 ;
        RECT 297.455 -204.705 297.685 -204.205 ;
        RECT 297.945 -204.850 298.175 -204.205 ;
        RECT 298.435 -204.705 298.665 -204.205 ;
        RECT 298.925 -204.850 299.155 -204.205 ;
        RECT 297.455 -205.080 300.640 -204.850 ;
        RECT 297.455 -205.860 297.685 -205.080 ;
        RECT 297.945 -205.090 299.155 -205.080 ;
        RECT 298.435 -205.860 298.665 -205.090 ;
        RECT 299.415 -205.860 299.645 -205.080 ;
        RECT 289.415 -210.355 289.645 -208.855 ;
        RECT 287.650 -211.330 288.635 -211.060 ;
        RECT 288.925 -213.035 289.155 -211.540 ;
        RECT 288.920 -213.220 289.155 -213.035 ;
        RECT 289.415 -213.040 289.645 -211.540 ;
        RECT 289.905 -213.220 290.135 -211.540 ;
        RECT 290.395 -213.040 290.625 -208.855 ;
        RECT 292.460 -209.630 292.690 -208.850 ;
        RECT 293.440 -209.620 293.670 -208.850 ;
        RECT 292.950 -209.630 294.160 -209.620 ;
        RECT 294.420 -209.630 294.650 -208.850 ;
        RECT 292.460 -209.860 295.645 -209.630 ;
        RECT 292.460 -210.505 292.690 -210.005 ;
        RECT 292.950 -210.505 293.180 -209.860 ;
        RECT 293.440 -210.505 293.670 -210.005 ;
        RECT 293.930 -210.505 294.160 -209.860 ;
        RECT 296.650 -211.410 296.880 -208.410 ;
        RECT 297.705 -211.410 297.935 -208.410 ;
        RECT 298.195 -211.410 298.425 -208.410 ;
        RECT 298.685 -211.410 298.915 -208.410 ;
        RECT 299.745 -211.410 299.975 -208.410 ;
        RECT 290.885 -213.220 291.115 -211.540 ;
        RECT 300.900 -212.065 301.425 -211.705 ;
        RECT 300.930 -212.480 301.255 -212.065 ;
        RECT 296.155 -212.805 301.255 -212.480 ;
        RECT 288.920 -213.455 291.115 -213.220 ;
        RECT 296.650 -214.470 296.880 -212.970 ;
        RECT 297.140 -214.470 297.370 -212.970 ;
        RECT 297.630 -214.470 297.860 -212.970 ;
        RECT 298.840 -214.470 299.070 -212.970 ;
        RECT 299.330 -214.470 299.560 -212.970 ;
        RECT 235.215 -215.590 256.940 -215.180 ;
        RECT 281.205 -215.010 284.590 -214.855 ;
        RECT 302.365 -215.010 302.930 -204.030 ;
        RECT 303.460 -211.735 304.565 -184.550 ;
        RECT 305.720 -200.415 306.910 -182.795 ;
        RECT 310.950 -183.820 312.200 -183.320 ;
        RECT 319.385 -183.740 321.580 -183.505 ;
        RECT 310.950 -184.090 317.940 -183.820 ;
        RECT 319.385 -183.925 319.620 -183.740 ;
        RECT 310.950 -184.465 312.200 -184.090 ;
        RECT 313.585 -186.290 314.235 -185.540 ;
        RECT 315.015 -185.810 315.245 -184.810 ;
        RECT 315.505 -185.950 315.735 -184.810 ;
        RECT 315.995 -185.810 316.225 -184.810 ;
        RECT 316.485 -185.950 316.715 -184.810 ;
        RECT 317.670 -185.540 317.940 -184.090 ;
        RECT 319.390 -185.420 319.620 -183.925 ;
        RECT 319.880 -185.420 320.110 -183.920 ;
        RECT 320.370 -185.420 320.600 -183.740 ;
        RECT 317.670 -185.810 319.310 -185.540 ;
        RECT 315.015 -186.180 318.200 -185.950 ;
        RECT 319.040 -186.085 319.310 -185.810 ;
        RECT 313.835 -193.310 314.105 -186.290 ;
        RECT 315.015 -187.460 315.245 -186.180 ;
        RECT 315.505 -186.190 316.715 -186.180 ;
        RECT 315.995 -187.460 316.225 -186.190 ;
        RECT 316.975 -187.460 317.205 -186.180 ;
        RECT 318.910 -186.375 319.705 -186.085 ;
        RECT 319.880 -188.105 320.110 -186.605 ;
        RECT 320.860 -188.105 321.090 -183.920 ;
        RECT 321.350 -185.420 321.580 -183.740 ;
        RECT 324.860 -186.280 328.400 -185.715 ;
        RECT 322.925 -186.955 323.155 -186.455 ;
        RECT 323.415 -187.100 323.645 -186.455 ;
        RECT 323.905 -186.955 324.135 -186.455 ;
        RECT 324.395 -187.100 324.625 -186.455 ;
        RECT 322.925 -187.330 326.110 -187.100 ;
        RECT 322.925 -188.110 323.155 -187.330 ;
        RECT 323.415 -187.340 324.625 -187.330 ;
        RECT 323.905 -188.110 324.135 -187.340 ;
        RECT 324.885 -188.110 325.115 -187.330 ;
        RECT 314.885 -192.605 315.115 -191.105 ;
        RECT 313.120 -193.580 314.105 -193.310 ;
        RECT 314.395 -195.285 314.625 -193.790 ;
        RECT 314.390 -195.470 314.625 -195.285 ;
        RECT 314.885 -195.290 315.115 -193.790 ;
        RECT 315.375 -195.470 315.605 -193.790 ;
        RECT 315.865 -195.290 316.095 -191.105 ;
        RECT 317.930 -191.880 318.160 -191.100 ;
        RECT 318.910 -191.870 319.140 -191.100 ;
        RECT 318.420 -191.880 319.630 -191.870 ;
        RECT 319.890 -191.880 320.120 -191.100 ;
        RECT 317.930 -192.110 321.115 -191.880 ;
        RECT 317.930 -192.755 318.160 -192.255 ;
        RECT 318.420 -192.755 318.650 -192.110 ;
        RECT 318.910 -192.755 319.140 -192.255 ;
        RECT 319.400 -192.755 319.630 -192.110 ;
        RECT 322.120 -193.660 322.350 -190.660 ;
        RECT 323.175 -193.660 323.405 -190.660 ;
        RECT 323.665 -193.660 323.895 -190.660 ;
        RECT 324.155 -193.660 324.385 -190.660 ;
        RECT 325.215 -193.660 325.445 -190.660 ;
        RECT 316.355 -195.470 316.585 -193.790 ;
        RECT 326.370 -194.315 326.895 -193.955 ;
        RECT 326.400 -194.730 326.725 -194.315 ;
        RECT 321.625 -195.055 326.725 -194.730 ;
        RECT 314.390 -195.705 316.585 -195.470 ;
        RECT 322.120 -196.720 322.350 -195.220 ;
        RECT 322.610 -196.720 322.840 -195.220 ;
        RECT 323.100 -196.720 323.330 -195.220 ;
        RECT 324.310 -196.720 324.540 -195.220 ;
        RECT 324.800 -196.720 325.030 -195.220 ;
        RECT 325.965 -197.260 326.530 -197.255 ;
        RECT 327.835 -197.260 328.400 -186.280 ;
        RECT 332.080 -192.450 332.310 -189.950 ;
        RECT 333.425 -192.450 333.655 -189.950 ;
        RECT 333.915 -192.450 334.145 -189.950 ;
        RECT 334.405 -192.450 334.635 -189.950 ;
        RECT 335.055 -192.450 335.285 -189.950 ;
        RECT 336.685 -192.450 336.915 -189.950 ;
        RECT 337.825 -191.450 338.055 -189.950 ;
        RECT 330.925 -193.250 331.615 -193.230 ;
        RECT 334.955 -193.250 335.645 -193.230 ;
        RECT 336.880 -193.250 337.150 -192.885 ;
        RECT 330.925 -193.470 337.150 -193.250 ;
        RECT 330.925 -193.500 331.615 -193.470 ;
        RECT 334.955 -193.500 335.645 -193.470 ;
        RECT 336.880 -193.575 337.150 -193.470 ;
        RECT 337.740 -193.650 338.070 -193.590 ;
        RECT 344.450 -193.650 345.640 -182.795 ;
        RECT 347.225 -183.005 348.110 -167.095 ;
        RECT 349.650 -182.835 391.590 -181.335 ;
        RECT 346.825 -184.460 348.515 -183.005 ;
        RECT 330.120 -195.185 330.635 -194.730 ;
        RECT 325.015 -197.825 328.400 -197.260 ;
        RECT 305.720 -201.085 311.400 -200.415 ;
        RECT 319.345 -201.005 321.540 -200.770 ;
        RECT 305.720 -201.355 317.900 -201.085 ;
        RECT 319.345 -201.190 319.580 -201.005 ;
        RECT 305.720 -201.605 311.400 -201.355 ;
        RECT 313.545 -203.555 314.195 -202.805 ;
        RECT 314.975 -203.075 315.205 -202.075 ;
        RECT 315.465 -203.215 315.695 -202.075 ;
        RECT 315.955 -203.075 316.185 -202.075 ;
        RECT 316.445 -203.215 316.675 -202.075 ;
        RECT 317.630 -202.805 317.900 -201.355 ;
        RECT 319.350 -202.685 319.580 -201.190 ;
        RECT 319.840 -202.685 320.070 -201.185 ;
        RECT 320.330 -202.685 320.560 -201.005 ;
        RECT 317.630 -203.075 319.270 -202.805 ;
        RECT 314.975 -203.445 318.160 -203.215 ;
        RECT 319.000 -203.350 319.270 -203.075 ;
        RECT 313.795 -210.575 314.065 -203.555 ;
        RECT 314.975 -204.725 315.205 -203.445 ;
        RECT 315.465 -203.455 316.675 -203.445 ;
        RECT 315.955 -204.725 316.185 -203.455 ;
        RECT 316.935 -204.725 317.165 -203.445 ;
        RECT 318.870 -203.640 319.665 -203.350 ;
        RECT 319.840 -205.370 320.070 -203.870 ;
        RECT 320.820 -205.370 321.050 -201.185 ;
        RECT 321.310 -202.685 321.540 -201.005 ;
        RECT 325.965 -202.980 326.530 -197.825 ;
        RECT 330.180 -198.350 330.575 -195.185 ;
        RECT 331.590 -196.430 331.820 -194.930 ;
        RECT 332.080 -196.430 332.310 -194.930 ;
        RECT 333.940 -196.430 334.170 -193.930 ;
        RECT 334.430 -196.430 334.660 -193.930 ;
        RECT 335.055 -196.430 335.285 -193.930 ;
        RECT 335.545 -196.430 335.775 -193.930 ;
        RECT 336.195 -196.430 336.425 -193.930 ;
        RECT 336.685 -196.430 336.915 -193.930 ;
        RECT 337.175 -196.430 337.405 -193.930 ;
        RECT 337.740 -193.960 345.850 -193.650 ;
        RECT 337.740 -194.005 338.070 -193.960 ;
        RECT 337.825 -196.430 338.055 -194.930 ;
        RECT 338.315 -196.430 338.545 -194.930 ;
        RECT 327.680 -198.745 330.575 -198.350 ;
        RECT 327.680 -200.520 328.075 -198.745 ;
        RECT 327.550 -201.005 328.130 -200.520 ;
        RECT 337.685 -201.160 339.880 -200.925 ;
        RECT 330.695 -201.240 331.180 -201.210 ;
        RECT 330.695 -201.510 336.240 -201.240 ;
        RECT 337.685 -201.345 337.920 -201.160 ;
        RECT 330.695 -201.540 331.180 -201.510 ;
        RECT 324.820 -203.545 328.360 -202.980 ;
        RECT 322.885 -204.220 323.115 -203.720 ;
        RECT 323.375 -204.365 323.605 -203.720 ;
        RECT 323.865 -204.220 324.095 -203.720 ;
        RECT 324.355 -204.365 324.585 -203.720 ;
        RECT 322.885 -204.595 326.070 -204.365 ;
        RECT 322.885 -205.375 323.115 -204.595 ;
        RECT 323.375 -204.605 324.585 -204.595 ;
        RECT 323.865 -205.375 324.095 -204.605 ;
        RECT 324.845 -205.375 325.075 -204.595 ;
        RECT 314.845 -209.870 315.075 -208.370 ;
        RECT 313.080 -210.845 314.065 -210.575 ;
        RECT 303.190 -213.230 304.650 -211.735 ;
        RECT 314.355 -212.550 314.585 -211.055 ;
        RECT 314.350 -212.735 314.585 -212.550 ;
        RECT 314.845 -212.555 315.075 -211.055 ;
        RECT 315.335 -212.735 315.565 -211.055 ;
        RECT 315.825 -212.555 316.055 -208.370 ;
        RECT 317.890 -209.145 318.120 -208.365 ;
        RECT 318.870 -209.135 319.100 -208.365 ;
        RECT 318.380 -209.145 319.590 -209.135 ;
        RECT 319.850 -209.145 320.080 -208.365 ;
        RECT 317.890 -209.375 321.075 -209.145 ;
        RECT 317.890 -210.020 318.120 -209.520 ;
        RECT 318.380 -210.020 318.610 -209.375 ;
        RECT 318.870 -210.020 319.100 -209.520 ;
        RECT 319.360 -210.020 319.590 -209.375 ;
        RECT 322.080 -210.925 322.310 -207.925 ;
        RECT 323.135 -210.925 323.365 -207.925 ;
        RECT 323.625 -210.925 323.855 -207.925 ;
        RECT 324.115 -210.925 324.345 -207.925 ;
        RECT 325.175 -210.925 325.405 -207.925 ;
        RECT 316.315 -212.735 316.545 -211.055 ;
        RECT 326.330 -211.580 326.855 -211.220 ;
        RECT 326.360 -211.995 326.685 -211.580 ;
        RECT 321.585 -212.320 326.685 -211.995 ;
        RECT 314.350 -212.970 316.545 -212.735 ;
        RECT 322.080 -213.985 322.310 -212.485 ;
        RECT 322.570 -213.985 322.800 -212.485 ;
        RECT 323.060 -213.985 323.290 -212.485 ;
        RECT 324.270 -213.985 324.500 -212.485 ;
        RECT 324.760 -213.985 324.990 -212.485 ;
        RECT 327.795 -214.525 328.360 -203.545 ;
        RECT 331.885 -203.710 332.535 -202.960 ;
        RECT 333.315 -203.230 333.545 -202.230 ;
        RECT 333.805 -203.370 334.035 -202.230 ;
        RECT 334.295 -203.230 334.525 -202.230 ;
        RECT 334.785 -203.370 335.015 -202.230 ;
        RECT 335.970 -202.960 336.240 -201.510 ;
        RECT 337.690 -202.840 337.920 -201.345 ;
        RECT 338.180 -202.840 338.410 -201.340 ;
        RECT 338.670 -202.840 338.900 -201.160 ;
        RECT 335.970 -203.230 337.610 -202.960 ;
        RECT 333.315 -203.600 336.500 -203.370 ;
        RECT 337.340 -203.505 337.610 -203.230 ;
        RECT 332.135 -210.730 332.405 -203.710 ;
        RECT 333.315 -204.880 333.545 -203.600 ;
        RECT 333.805 -203.610 335.015 -203.600 ;
        RECT 334.295 -204.880 334.525 -203.610 ;
        RECT 335.275 -204.880 335.505 -203.600 ;
        RECT 337.210 -203.795 338.005 -203.505 ;
        RECT 338.180 -205.525 338.410 -204.025 ;
        RECT 339.160 -205.525 339.390 -201.340 ;
        RECT 339.650 -202.840 339.880 -201.160 ;
        RECT 343.160 -203.700 346.700 -203.135 ;
        RECT 341.225 -204.375 341.455 -203.875 ;
        RECT 341.715 -204.520 341.945 -203.875 ;
        RECT 342.205 -204.375 342.435 -203.875 ;
        RECT 342.695 -204.520 342.925 -203.875 ;
        RECT 341.225 -204.750 344.410 -204.520 ;
        RECT 341.225 -205.530 341.455 -204.750 ;
        RECT 341.715 -204.760 342.925 -204.750 ;
        RECT 342.205 -205.530 342.435 -204.760 ;
        RECT 343.185 -205.530 343.415 -204.750 ;
        RECT 333.185 -210.025 333.415 -208.525 ;
        RECT 331.420 -211.000 332.405 -210.730 ;
        RECT 332.695 -212.705 332.925 -211.210 ;
        RECT 332.690 -212.890 332.925 -212.705 ;
        RECT 333.185 -212.710 333.415 -211.210 ;
        RECT 333.675 -212.890 333.905 -211.210 ;
        RECT 334.165 -212.710 334.395 -208.525 ;
        RECT 336.230 -209.300 336.460 -208.520 ;
        RECT 337.210 -209.290 337.440 -208.520 ;
        RECT 336.720 -209.300 337.930 -209.290 ;
        RECT 338.190 -209.300 338.420 -208.520 ;
        RECT 336.230 -209.530 339.415 -209.300 ;
        RECT 336.230 -210.175 336.460 -209.675 ;
        RECT 336.720 -210.175 336.950 -209.530 ;
        RECT 337.210 -210.175 337.440 -209.675 ;
        RECT 337.700 -210.175 337.930 -209.530 ;
        RECT 340.420 -211.080 340.650 -208.080 ;
        RECT 341.475 -211.080 341.705 -208.080 ;
        RECT 341.965 -211.080 342.195 -208.080 ;
        RECT 342.455 -211.080 342.685 -208.080 ;
        RECT 343.515 -211.080 343.745 -208.080 ;
        RECT 334.655 -212.890 334.885 -211.210 ;
        RECT 344.670 -211.735 345.195 -211.375 ;
        RECT 344.700 -212.150 345.025 -211.735 ;
        RECT 339.925 -212.475 345.025 -212.150 ;
        RECT 332.690 -213.125 334.885 -212.890 ;
        RECT 340.420 -214.140 340.650 -212.640 ;
        RECT 340.910 -214.140 341.140 -212.640 ;
        RECT 341.400 -214.140 341.630 -212.640 ;
        RECT 342.610 -214.140 342.840 -212.640 ;
        RECT 343.100 -214.140 343.330 -212.640 ;
        RECT 281.205 -215.420 302.930 -215.010 ;
        RECT 324.975 -214.680 328.360 -214.525 ;
        RECT 346.135 -214.680 346.700 -203.700 ;
        RECT 347.225 -211.445 348.110 -184.460 ;
        RECT 349.650 -200.085 351.150 -182.835 ;
        RECT 356.765 -183.735 358.105 -183.280 ;
        RECT 365.150 -183.655 367.345 -183.420 ;
        RECT 356.765 -184.005 363.705 -183.735 ;
        RECT 365.150 -183.840 365.385 -183.655 ;
        RECT 356.765 -184.480 358.105 -184.005 ;
        RECT 359.350 -186.205 360.000 -185.455 ;
        RECT 360.780 -185.725 361.010 -184.725 ;
        RECT 361.270 -185.865 361.500 -184.725 ;
        RECT 361.760 -185.725 361.990 -184.725 ;
        RECT 362.250 -185.865 362.480 -184.725 ;
        RECT 363.435 -185.455 363.705 -184.005 ;
        RECT 365.155 -185.335 365.385 -183.840 ;
        RECT 365.645 -185.335 365.875 -183.835 ;
        RECT 366.135 -185.335 366.365 -183.655 ;
        RECT 363.435 -185.725 365.075 -185.455 ;
        RECT 360.780 -186.095 363.965 -185.865 ;
        RECT 364.805 -186.000 365.075 -185.725 ;
        RECT 359.600 -193.225 359.870 -186.205 ;
        RECT 360.780 -187.375 361.010 -186.095 ;
        RECT 361.270 -186.105 362.480 -186.095 ;
        RECT 361.760 -187.375 361.990 -186.105 ;
        RECT 362.740 -187.375 362.970 -186.095 ;
        RECT 364.675 -186.290 365.470 -186.000 ;
        RECT 365.645 -188.020 365.875 -186.520 ;
        RECT 366.625 -188.020 366.855 -183.835 ;
        RECT 367.115 -185.335 367.345 -183.655 ;
        RECT 370.625 -186.195 374.165 -185.630 ;
        RECT 368.690 -186.870 368.920 -186.370 ;
        RECT 369.180 -187.015 369.410 -186.370 ;
        RECT 369.670 -186.870 369.900 -186.370 ;
        RECT 370.160 -187.015 370.390 -186.370 ;
        RECT 368.690 -187.245 371.875 -187.015 ;
        RECT 368.690 -188.025 368.920 -187.245 ;
        RECT 369.180 -187.255 370.390 -187.245 ;
        RECT 369.670 -188.025 369.900 -187.255 ;
        RECT 370.650 -188.025 370.880 -187.245 ;
        RECT 360.650 -192.520 360.880 -191.020 ;
        RECT 358.885 -193.495 359.870 -193.225 ;
        RECT 360.160 -195.200 360.390 -193.705 ;
        RECT 360.155 -195.385 360.390 -195.200 ;
        RECT 360.650 -195.205 360.880 -193.705 ;
        RECT 361.140 -195.385 361.370 -193.705 ;
        RECT 361.630 -195.205 361.860 -191.020 ;
        RECT 363.695 -191.795 363.925 -191.015 ;
        RECT 364.675 -191.785 364.905 -191.015 ;
        RECT 364.185 -191.795 365.395 -191.785 ;
        RECT 365.655 -191.795 365.885 -191.015 ;
        RECT 363.695 -192.025 366.880 -191.795 ;
        RECT 363.695 -192.670 363.925 -192.170 ;
        RECT 364.185 -192.670 364.415 -192.025 ;
        RECT 364.675 -192.670 364.905 -192.170 ;
        RECT 365.165 -192.670 365.395 -192.025 ;
        RECT 367.885 -193.575 368.115 -190.575 ;
        RECT 368.940 -193.575 369.170 -190.575 ;
        RECT 369.430 -193.575 369.660 -190.575 ;
        RECT 369.920 -193.575 370.150 -190.575 ;
        RECT 370.980 -193.575 371.210 -190.575 ;
        RECT 362.120 -195.385 362.350 -193.705 ;
        RECT 372.135 -194.230 372.660 -193.870 ;
        RECT 372.165 -194.645 372.490 -194.230 ;
        RECT 367.390 -194.970 372.490 -194.645 ;
        RECT 360.155 -195.620 362.350 -195.385 ;
        RECT 367.885 -196.635 368.115 -195.135 ;
        RECT 368.375 -196.635 368.605 -195.135 ;
        RECT 368.865 -196.635 369.095 -195.135 ;
        RECT 370.075 -196.635 370.305 -195.135 ;
        RECT 370.565 -196.635 370.795 -195.135 ;
        RECT 371.730 -197.175 372.295 -197.170 ;
        RECT 373.600 -197.175 374.165 -186.195 ;
        RECT 377.845 -192.365 378.075 -189.865 ;
        RECT 379.190 -192.365 379.420 -189.865 ;
        RECT 379.680 -192.365 379.910 -189.865 ;
        RECT 380.170 -192.365 380.400 -189.865 ;
        RECT 380.820 -192.365 381.050 -189.865 ;
        RECT 382.450 -192.365 382.680 -189.865 ;
        RECT 383.590 -191.365 383.820 -189.865 ;
        RECT 376.690 -193.165 377.380 -193.145 ;
        RECT 380.720 -193.165 381.410 -193.145 ;
        RECT 382.645 -193.165 382.915 -192.800 ;
        RECT 376.690 -193.385 382.915 -193.165 ;
        RECT 376.690 -193.415 377.380 -193.385 ;
        RECT 380.720 -193.415 381.410 -193.385 ;
        RECT 382.645 -193.490 382.915 -193.385 ;
        RECT 383.505 -193.565 383.835 -193.505 ;
        RECT 390.055 -193.565 391.590 -182.835 ;
        RECT 375.885 -195.100 376.400 -194.645 ;
        RECT 370.780 -197.740 374.165 -197.175 ;
        RECT 349.650 -201.000 357.100 -200.085 ;
        RECT 365.110 -200.920 367.305 -200.685 ;
        RECT 349.650 -201.270 363.665 -201.000 ;
        RECT 365.110 -201.105 365.345 -200.920 ;
        RECT 349.650 -201.585 357.100 -201.270 ;
        RECT 359.310 -203.470 359.960 -202.720 ;
        RECT 360.740 -202.990 360.970 -201.990 ;
        RECT 361.230 -203.130 361.460 -201.990 ;
        RECT 361.720 -202.990 361.950 -201.990 ;
        RECT 362.210 -203.130 362.440 -201.990 ;
        RECT 363.395 -202.720 363.665 -201.270 ;
        RECT 365.115 -202.600 365.345 -201.105 ;
        RECT 365.605 -202.600 365.835 -201.100 ;
        RECT 366.095 -202.600 366.325 -200.920 ;
        RECT 363.395 -202.990 365.035 -202.720 ;
        RECT 360.740 -203.360 363.925 -203.130 ;
        RECT 364.765 -203.265 365.035 -202.990 ;
        RECT 359.560 -210.490 359.830 -203.470 ;
        RECT 360.740 -204.640 360.970 -203.360 ;
        RECT 361.230 -203.370 362.440 -203.360 ;
        RECT 361.720 -204.640 361.950 -203.370 ;
        RECT 362.700 -204.640 362.930 -203.360 ;
        RECT 364.635 -203.555 365.430 -203.265 ;
        RECT 365.605 -205.285 365.835 -203.785 ;
        RECT 366.585 -205.285 366.815 -201.100 ;
        RECT 367.075 -202.600 367.305 -200.920 ;
        RECT 371.730 -202.895 372.295 -197.740 ;
        RECT 375.945 -198.265 376.340 -195.100 ;
        RECT 377.355 -196.345 377.585 -194.845 ;
        RECT 377.845 -196.345 378.075 -194.845 ;
        RECT 379.705 -196.345 379.935 -193.845 ;
        RECT 380.195 -196.345 380.425 -193.845 ;
        RECT 380.820 -196.345 381.050 -193.845 ;
        RECT 381.310 -196.345 381.540 -193.845 ;
        RECT 381.960 -196.345 382.190 -193.845 ;
        RECT 382.450 -196.345 382.680 -193.845 ;
        RECT 382.940 -196.345 383.170 -193.845 ;
        RECT 383.505 -193.875 391.615 -193.565 ;
        RECT 383.505 -193.920 383.835 -193.875 ;
        RECT 383.590 -196.345 383.820 -194.845 ;
        RECT 384.080 -196.345 384.310 -194.845 ;
        RECT 373.445 -198.660 376.340 -198.265 ;
        RECT 373.445 -200.435 373.840 -198.660 ;
        RECT 373.315 -200.920 373.895 -200.435 ;
        RECT 383.450 -201.075 385.645 -200.840 ;
        RECT 376.460 -201.155 376.945 -201.125 ;
        RECT 376.460 -201.425 382.005 -201.155 ;
        RECT 383.450 -201.260 383.685 -201.075 ;
        RECT 376.460 -201.455 376.945 -201.425 ;
        RECT 370.585 -203.460 374.125 -202.895 ;
        RECT 368.650 -204.135 368.880 -203.635 ;
        RECT 369.140 -204.280 369.370 -203.635 ;
        RECT 369.630 -204.135 369.860 -203.635 ;
        RECT 370.120 -204.280 370.350 -203.635 ;
        RECT 368.650 -204.510 371.835 -204.280 ;
        RECT 368.650 -205.290 368.880 -204.510 ;
        RECT 369.140 -204.520 370.350 -204.510 ;
        RECT 369.630 -205.290 369.860 -204.520 ;
        RECT 370.610 -205.290 370.840 -204.510 ;
        RECT 360.610 -209.785 360.840 -208.285 ;
        RECT 358.845 -210.760 359.830 -210.490 ;
        RECT 347.015 -212.965 348.320 -211.445 ;
        RECT 360.120 -212.465 360.350 -210.970 ;
        RECT 360.115 -212.650 360.350 -212.465 ;
        RECT 360.610 -212.470 360.840 -210.970 ;
        RECT 361.100 -212.650 361.330 -210.970 ;
        RECT 361.590 -212.470 361.820 -208.285 ;
        RECT 363.655 -209.060 363.885 -208.280 ;
        RECT 364.635 -209.050 364.865 -208.280 ;
        RECT 364.145 -209.060 365.355 -209.050 ;
        RECT 365.615 -209.060 365.845 -208.280 ;
        RECT 363.655 -209.290 366.840 -209.060 ;
        RECT 363.655 -209.935 363.885 -209.435 ;
        RECT 364.145 -209.935 364.375 -209.290 ;
        RECT 364.635 -209.935 364.865 -209.435 ;
        RECT 365.125 -209.935 365.355 -209.290 ;
        RECT 367.845 -210.840 368.075 -207.840 ;
        RECT 368.900 -210.840 369.130 -207.840 ;
        RECT 369.390 -210.840 369.620 -207.840 ;
        RECT 369.880 -210.840 370.110 -207.840 ;
        RECT 370.940 -210.840 371.170 -207.840 ;
        RECT 362.080 -212.650 362.310 -210.970 ;
        RECT 372.095 -211.495 372.620 -211.135 ;
        RECT 372.125 -211.910 372.450 -211.495 ;
        RECT 367.350 -212.235 372.450 -211.910 ;
        RECT 360.115 -212.885 362.310 -212.650 ;
        RECT 367.845 -213.900 368.075 -212.400 ;
        RECT 368.335 -213.900 368.565 -212.400 ;
        RECT 368.825 -213.900 369.055 -212.400 ;
        RECT 370.035 -213.900 370.265 -212.400 ;
        RECT 370.525 -213.900 370.755 -212.400 ;
        RECT 373.560 -214.440 374.125 -203.460 ;
        RECT 377.650 -203.625 378.300 -202.875 ;
        RECT 379.080 -203.145 379.310 -202.145 ;
        RECT 379.570 -203.285 379.800 -202.145 ;
        RECT 380.060 -203.145 380.290 -202.145 ;
        RECT 380.550 -203.285 380.780 -202.145 ;
        RECT 381.735 -202.875 382.005 -201.425 ;
        RECT 383.455 -202.755 383.685 -201.260 ;
        RECT 383.945 -202.755 384.175 -201.255 ;
        RECT 384.435 -202.755 384.665 -201.075 ;
        RECT 381.735 -203.145 383.375 -202.875 ;
        RECT 379.080 -203.515 382.265 -203.285 ;
        RECT 383.105 -203.420 383.375 -203.145 ;
        RECT 377.900 -210.645 378.170 -203.625 ;
        RECT 379.080 -204.795 379.310 -203.515 ;
        RECT 379.570 -203.525 380.780 -203.515 ;
        RECT 380.060 -204.795 380.290 -203.525 ;
        RECT 381.040 -204.795 381.270 -203.515 ;
        RECT 382.975 -203.710 383.770 -203.420 ;
        RECT 383.945 -205.440 384.175 -203.940 ;
        RECT 384.925 -205.440 385.155 -201.255 ;
        RECT 385.415 -202.755 385.645 -201.075 ;
        RECT 388.925 -203.615 392.465 -203.050 ;
        RECT 386.990 -204.290 387.220 -203.790 ;
        RECT 387.480 -204.435 387.710 -203.790 ;
        RECT 387.970 -204.290 388.200 -203.790 ;
        RECT 388.460 -204.435 388.690 -203.790 ;
        RECT 386.990 -204.665 390.175 -204.435 ;
        RECT 386.990 -205.445 387.220 -204.665 ;
        RECT 387.480 -204.675 388.690 -204.665 ;
        RECT 387.970 -205.445 388.200 -204.675 ;
        RECT 388.950 -205.445 389.180 -204.665 ;
        RECT 378.950 -209.940 379.180 -208.440 ;
        RECT 377.185 -210.915 378.170 -210.645 ;
        RECT 378.460 -212.620 378.690 -211.125 ;
        RECT 378.455 -212.805 378.690 -212.620 ;
        RECT 378.950 -212.625 379.180 -211.125 ;
        RECT 379.440 -212.805 379.670 -211.125 ;
        RECT 379.930 -212.625 380.160 -208.440 ;
        RECT 381.995 -209.215 382.225 -208.435 ;
        RECT 382.975 -209.205 383.205 -208.435 ;
        RECT 382.485 -209.215 383.695 -209.205 ;
        RECT 383.955 -209.215 384.185 -208.435 ;
        RECT 381.995 -209.445 385.180 -209.215 ;
        RECT 381.995 -210.090 382.225 -209.590 ;
        RECT 382.485 -210.090 382.715 -209.445 ;
        RECT 382.975 -210.090 383.205 -209.590 ;
        RECT 383.465 -210.090 383.695 -209.445 ;
        RECT 386.185 -210.995 386.415 -207.995 ;
        RECT 387.240 -210.995 387.470 -207.995 ;
        RECT 387.730 -210.995 387.960 -207.995 ;
        RECT 388.220 -210.995 388.450 -207.995 ;
        RECT 389.280 -210.995 389.510 -207.995 ;
        RECT 380.420 -212.805 380.650 -211.125 ;
        RECT 390.435 -211.650 390.960 -211.290 ;
        RECT 390.465 -212.065 390.790 -211.650 ;
        RECT 385.690 -212.390 390.790 -212.065 ;
        RECT 378.455 -213.040 380.650 -212.805 ;
        RECT 386.185 -214.055 386.415 -212.555 ;
        RECT 386.675 -214.055 386.905 -212.555 ;
        RECT 387.165 -214.055 387.395 -212.555 ;
        RECT 388.375 -214.055 388.605 -212.555 ;
        RECT 388.865 -214.055 389.095 -212.555 ;
        RECT 324.975 -215.090 346.700 -214.680 ;
        RECT 370.740 -214.595 374.125 -214.440 ;
        RECT 391.900 -214.595 392.465 -203.615 ;
        RECT 392.895 -213.065 394.450 -164.845 ;
        RECT 395.775 -182.425 438.370 -181.330 ;
        RECT 395.775 -200.615 396.870 -182.425 ;
        RECT 403.040 -183.545 404.515 -182.970 ;
        RECT 411.970 -183.465 414.165 -183.230 ;
        RECT 403.040 -183.815 410.525 -183.545 ;
        RECT 411.970 -183.650 412.205 -183.465 ;
        RECT 403.040 -184.335 404.515 -183.815 ;
        RECT 406.170 -186.015 406.820 -185.265 ;
        RECT 407.600 -185.535 407.830 -184.535 ;
        RECT 408.090 -185.675 408.320 -184.535 ;
        RECT 408.580 -185.535 408.810 -184.535 ;
        RECT 409.070 -185.675 409.300 -184.535 ;
        RECT 410.255 -185.265 410.525 -183.815 ;
        RECT 411.975 -185.145 412.205 -183.650 ;
        RECT 412.465 -185.145 412.695 -183.645 ;
        RECT 412.955 -185.145 413.185 -183.465 ;
        RECT 410.255 -185.535 411.895 -185.265 ;
        RECT 407.600 -185.905 410.785 -185.675 ;
        RECT 411.625 -185.810 411.895 -185.535 ;
        RECT 406.420 -193.035 406.690 -186.015 ;
        RECT 407.600 -187.185 407.830 -185.905 ;
        RECT 408.090 -185.915 409.300 -185.905 ;
        RECT 408.580 -187.185 408.810 -185.915 ;
        RECT 409.560 -187.185 409.790 -185.905 ;
        RECT 411.495 -186.100 412.290 -185.810 ;
        RECT 412.465 -187.830 412.695 -186.330 ;
        RECT 413.445 -187.830 413.675 -183.645 ;
        RECT 413.935 -185.145 414.165 -183.465 ;
        RECT 417.445 -186.005 420.985 -185.440 ;
        RECT 415.510 -186.680 415.740 -186.180 ;
        RECT 416.000 -186.825 416.230 -186.180 ;
        RECT 416.490 -186.680 416.720 -186.180 ;
        RECT 416.980 -186.825 417.210 -186.180 ;
        RECT 415.510 -187.055 418.695 -186.825 ;
        RECT 415.510 -187.835 415.740 -187.055 ;
        RECT 416.000 -187.065 417.210 -187.055 ;
        RECT 416.490 -187.835 416.720 -187.065 ;
        RECT 417.470 -187.835 417.700 -187.055 ;
        RECT 407.470 -192.330 407.700 -190.830 ;
        RECT 405.705 -193.305 406.690 -193.035 ;
        RECT 406.980 -195.010 407.210 -193.515 ;
        RECT 406.975 -195.195 407.210 -195.010 ;
        RECT 407.470 -195.015 407.700 -193.515 ;
        RECT 407.960 -195.195 408.190 -193.515 ;
        RECT 408.450 -195.015 408.680 -190.830 ;
        RECT 410.515 -191.605 410.745 -190.825 ;
        RECT 411.495 -191.595 411.725 -190.825 ;
        RECT 411.005 -191.605 412.215 -191.595 ;
        RECT 412.475 -191.605 412.705 -190.825 ;
        RECT 410.515 -191.835 413.700 -191.605 ;
        RECT 410.515 -192.480 410.745 -191.980 ;
        RECT 411.005 -192.480 411.235 -191.835 ;
        RECT 411.495 -192.480 411.725 -191.980 ;
        RECT 411.985 -192.480 412.215 -191.835 ;
        RECT 414.705 -193.385 414.935 -190.385 ;
        RECT 415.760 -193.385 415.990 -190.385 ;
        RECT 416.250 -193.385 416.480 -190.385 ;
        RECT 416.740 -193.385 416.970 -190.385 ;
        RECT 417.800 -193.385 418.030 -190.385 ;
        RECT 408.940 -195.195 409.170 -193.515 ;
        RECT 418.955 -194.040 419.480 -193.680 ;
        RECT 418.985 -194.455 419.310 -194.040 ;
        RECT 414.210 -194.780 419.310 -194.455 ;
        RECT 406.975 -195.430 409.170 -195.195 ;
        RECT 414.705 -196.445 414.935 -194.945 ;
        RECT 415.195 -196.445 415.425 -194.945 ;
        RECT 415.685 -196.445 415.915 -194.945 ;
        RECT 416.895 -196.445 417.125 -194.945 ;
        RECT 417.385 -196.445 417.615 -194.945 ;
        RECT 418.550 -196.985 419.115 -196.980 ;
        RECT 420.420 -196.985 420.985 -186.005 ;
        RECT 424.665 -192.175 424.895 -189.675 ;
        RECT 426.010 -192.175 426.240 -189.675 ;
        RECT 426.500 -192.175 426.730 -189.675 ;
        RECT 426.990 -192.175 427.220 -189.675 ;
        RECT 427.640 -192.175 427.870 -189.675 ;
        RECT 429.270 -192.175 429.500 -189.675 ;
        RECT 430.410 -191.175 430.640 -189.675 ;
        RECT 423.510 -192.975 424.200 -192.955 ;
        RECT 427.540 -192.975 428.230 -192.955 ;
        RECT 429.465 -192.975 429.735 -192.610 ;
        RECT 423.510 -193.195 429.735 -192.975 ;
        RECT 423.510 -193.225 424.200 -193.195 ;
        RECT 427.540 -193.225 428.230 -193.195 ;
        RECT 429.465 -193.300 429.735 -193.195 ;
        RECT 430.325 -193.375 430.655 -193.315 ;
        RECT 437.275 -193.375 438.370 -182.425 ;
        RECT 422.705 -194.910 423.220 -194.455 ;
        RECT 417.600 -197.550 420.985 -196.985 ;
        RECT 395.775 -200.810 404.670 -200.615 ;
        RECT 411.930 -200.730 414.125 -200.495 ;
        RECT 395.775 -201.080 410.485 -200.810 ;
        RECT 411.930 -200.915 412.165 -200.730 ;
        RECT 395.775 -201.710 404.670 -201.080 ;
        RECT 406.130 -203.280 406.780 -202.530 ;
        RECT 407.560 -202.800 407.790 -201.800 ;
        RECT 408.050 -202.940 408.280 -201.800 ;
        RECT 408.540 -202.800 408.770 -201.800 ;
        RECT 409.030 -202.940 409.260 -201.800 ;
        RECT 410.215 -202.530 410.485 -201.080 ;
        RECT 411.935 -202.410 412.165 -200.915 ;
        RECT 412.425 -202.410 412.655 -200.910 ;
        RECT 412.915 -202.410 413.145 -200.730 ;
        RECT 410.215 -202.800 411.855 -202.530 ;
        RECT 407.560 -203.170 410.745 -202.940 ;
        RECT 411.585 -203.075 411.855 -202.800 ;
        RECT 406.380 -210.300 406.650 -203.280 ;
        RECT 407.560 -204.450 407.790 -203.170 ;
        RECT 408.050 -203.180 409.260 -203.170 ;
        RECT 408.540 -204.450 408.770 -203.180 ;
        RECT 409.520 -204.450 409.750 -203.170 ;
        RECT 411.455 -203.365 412.250 -203.075 ;
        RECT 412.425 -205.095 412.655 -203.595 ;
        RECT 413.405 -205.095 413.635 -200.910 ;
        RECT 413.895 -202.410 414.125 -200.730 ;
        RECT 418.550 -202.705 419.115 -197.550 ;
        RECT 422.765 -198.075 423.160 -194.910 ;
        RECT 424.175 -196.155 424.405 -194.655 ;
        RECT 424.665 -196.155 424.895 -194.655 ;
        RECT 426.525 -196.155 426.755 -193.655 ;
        RECT 427.015 -196.155 427.245 -193.655 ;
        RECT 427.640 -196.155 427.870 -193.655 ;
        RECT 428.130 -196.155 428.360 -193.655 ;
        RECT 428.780 -196.155 429.010 -193.655 ;
        RECT 429.270 -196.155 429.500 -193.655 ;
        RECT 429.760 -196.155 429.990 -193.655 ;
        RECT 430.325 -193.685 438.435 -193.375 ;
        RECT 430.325 -193.730 430.655 -193.685 ;
        RECT 430.410 -196.155 430.640 -194.655 ;
        RECT 430.900 -196.155 431.130 -194.655 ;
        RECT 420.265 -198.470 423.160 -198.075 ;
        RECT 420.265 -200.245 420.660 -198.470 ;
        RECT 420.135 -200.730 420.715 -200.245 ;
        RECT 430.270 -200.885 432.465 -200.650 ;
        RECT 423.280 -200.965 423.765 -200.935 ;
        RECT 423.280 -201.235 428.825 -200.965 ;
        RECT 430.270 -201.070 430.505 -200.885 ;
        RECT 423.280 -201.265 423.765 -201.235 ;
        RECT 417.405 -203.270 420.945 -202.705 ;
        RECT 415.470 -203.945 415.700 -203.445 ;
        RECT 415.960 -204.090 416.190 -203.445 ;
        RECT 416.450 -203.945 416.680 -203.445 ;
        RECT 416.940 -204.090 417.170 -203.445 ;
        RECT 415.470 -204.320 418.655 -204.090 ;
        RECT 415.470 -205.100 415.700 -204.320 ;
        RECT 415.960 -204.330 417.170 -204.320 ;
        RECT 416.450 -205.100 416.680 -204.330 ;
        RECT 417.430 -205.100 417.660 -204.320 ;
        RECT 407.430 -209.595 407.660 -208.095 ;
        RECT 405.665 -210.570 406.650 -210.300 ;
        RECT 406.940 -212.275 407.170 -210.780 ;
        RECT 406.935 -212.460 407.170 -212.275 ;
        RECT 407.430 -212.280 407.660 -210.780 ;
        RECT 407.920 -212.460 408.150 -210.780 ;
        RECT 408.410 -212.280 408.640 -208.095 ;
        RECT 410.475 -208.870 410.705 -208.090 ;
        RECT 411.455 -208.860 411.685 -208.090 ;
        RECT 410.965 -208.870 412.175 -208.860 ;
        RECT 412.435 -208.870 412.665 -208.090 ;
        RECT 410.475 -209.100 413.660 -208.870 ;
        RECT 410.475 -209.745 410.705 -209.245 ;
        RECT 410.965 -209.745 411.195 -209.100 ;
        RECT 411.455 -209.745 411.685 -209.245 ;
        RECT 411.945 -209.745 412.175 -209.100 ;
        RECT 414.665 -210.650 414.895 -207.650 ;
        RECT 415.720 -210.650 415.950 -207.650 ;
        RECT 416.210 -210.650 416.440 -207.650 ;
        RECT 416.700 -210.650 416.930 -207.650 ;
        RECT 417.760 -210.650 417.990 -207.650 ;
        RECT 408.900 -212.460 409.130 -210.780 ;
        RECT 418.915 -211.305 419.440 -210.945 ;
        RECT 418.945 -211.720 419.270 -211.305 ;
        RECT 414.170 -212.045 419.270 -211.720 ;
        RECT 406.935 -212.695 409.130 -212.460 ;
        RECT 414.665 -213.710 414.895 -212.210 ;
        RECT 415.155 -213.710 415.385 -212.210 ;
        RECT 415.645 -213.710 415.875 -212.210 ;
        RECT 416.855 -213.710 417.085 -212.210 ;
        RECT 417.345 -213.710 417.575 -212.210 ;
        RECT 420.380 -214.250 420.945 -203.270 ;
        RECT 424.470 -203.435 425.120 -202.685 ;
        RECT 425.900 -202.955 426.130 -201.955 ;
        RECT 426.390 -203.095 426.620 -201.955 ;
        RECT 426.880 -202.955 427.110 -201.955 ;
        RECT 427.370 -203.095 427.600 -201.955 ;
        RECT 428.555 -202.685 428.825 -201.235 ;
        RECT 430.275 -202.565 430.505 -201.070 ;
        RECT 430.765 -202.565 430.995 -201.065 ;
        RECT 431.255 -202.565 431.485 -200.885 ;
        RECT 428.555 -202.955 430.195 -202.685 ;
        RECT 425.900 -203.325 429.085 -203.095 ;
        RECT 429.925 -203.230 430.195 -202.955 ;
        RECT 424.720 -210.455 424.990 -203.435 ;
        RECT 425.900 -204.605 426.130 -203.325 ;
        RECT 426.390 -203.335 427.600 -203.325 ;
        RECT 426.880 -204.605 427.110 -203.335 ;
        RECT 427.860 -204.605 428.090 -203.325 ;
        RECT 429.795 -203.520 430.590 -203.230 ;
        RECT 430.765 -205.250 430.995 -203.750 ;
        RECT 431.745 -205.250 431.975 -201.065 ;
        RECT 432.235 -202.565 432.465 -200.885 ;
        RECT 435.745 -203.425 439.285 -202.860 ;
        RECT 433.810 -204.100 434.040 -203.600 ;
        RECT 434.300 -204.245 434.530 -203.600 ;
        RECT 434.790 -204.100 435.020 -203.600 ;
        RECT 435.280 -204.245 435.510 -203.600 ;
        RECT 433.810 -204.475 436.995 -204.245 ;
        RECT 433.810 -205.255 434.040 -204.475 ;
        RECT 434.300 -204.485 435.510 -204.475 ;
        RECT 434.790 -205.255 435.020 -204.485 ;
        RECT 435.770 -205.255 436.000 -204.475 ;
        RECT 425.770 -209.750 426.000 -208.250 ;
        RECT 424.005 -210.725 424.990 -210.455 ;
        RECT 425.280 -212.430 425.510 -210.935 ;
        RECT 425.275 -212.615 425.510 -212.430 ;
        RECT 425.770 -212.435 426.000 -210.935 ;
        RECT 426.260 -212.615 426.490 -210.935 ;
        RECT 426.750 -212.435 426.980 -208.250 ;
        RECT 428.815 -209.025 429.045 -208.245 ;
        RECT 429.795 -209.015 430.025 -208.245 ;
        RECT 429.305 -209.025 430.515 -209.015 ;
        RECT 430.775 -209.025 431.005 -208.245 ;
        RECT 428.815 -209.255 432.000 -209.025 ;
        RECT 428.815 -209.900 429.045 -209.400 ;
        RECT 429.305 -209.900 429.535 -209.255 ;
        RECT 429.795 -209.900 430.025 -209.400 ;
        RECT 430.285 -209.900 430.515 -209.255 ;
        RECT 433.005 -210.805 433.235 -207.805 ;
        RECT 434.060 -210.805 434.290 -207.805 ;
        RECT 434.550 -210.805 434.780 -207.805 ;
        RECT 435.040 -210.805 435.270 -207.805 ;
        RECT 436.100 -210.805 436.330 -207.805 ;
        RECT 427.240 -212.615 427.470 -210.935 ;
        RECT 437.255 -211.460 437.780 -211.100 ;
        RECT 437.285 -211.875 437.610 -211.460 ;
        RECT 432.510 -212.200 437.610 -211.875 ;
        RECT 425.275 -212.850 427.470 -212.615 ;
        RECT 433.005 -213.865 433.235 -212.365 ;
        RECT 433.495 -213.865 433.725 -212.365 ;
        RECT 433.985 -213.865 434.215 -212.365 ;
        RECT 435.195 -213.865 435.425 -212.365 ;
        RECT 435.685 -213.865 435.915 -212.365 ;
        RECT 370.740 -215.005 392.465 -214.595 ;
        RECT 417.560 -214.405 420.945 -214.250 ;
        RECT 438.720 -214.405 439.285 -203.425 ;
        RECT 440.550 -211.225 441.970 -160.180 ;
        RECT 440.400 -212.940 442.195 -211.225 ;
        RECT 417.560 -214.815 439.285 -214.405 ;
        RECT 417.580 -214.970 439.285 -214.815 ;
        RECT 324.995 -215.245 346.700 -215.090 ;
        RECT 370.760 -215.160 392.465 -215.005 ;
        RECT 281.225 -215.575 302.930 -215.420 ;
        RECT 235.235 -215.745 256.940 -215.590 ;
        RECT 211.375 -218.615 212.960 -218.200 ;
        RECT 132.875 -219.520 176.875 -218.615 ;
        RECT 211.375 -219.520 410.125 -218.615 ;
        RECT 211.375 -219.655 212.960 -219.520 ;
        RECT 211.160 -224.115 213.005 -222.230 ;
        RECT 217.760 -223.720 410.125 -222.295 ;
        RECT 211.205 -233.055 212.705 -224.115 ;
        RECT 123.815 -234.555 212.705 -233.055 ;
        RECT 217.760 -235.770 219.185 -223.720 ;
        RECT 122.790 -236.065 219.185 -235.770 ;
        RECT 121.475 -236.670 219.185 -236.065 ;
        RECT 122.790 -237.195 219.185 -236.670 ;
        RECT 67.380 -250.735 445.485 -249.315 ;
        RECT -143.200 -261.510 -141.200 -261.280 ;
        RECT -143.200 -262.100 -141.200 -261.870 ;
        RECT -143.200 -262.690 -141.200 -262.460 ;
        RECT -147.680 -302.970 -145.405 -263.080 ;
        RECT -143.200 -263.280 -141.200 -263.050 ;
        RECT -143.200 -263.870 -141.200 -263.640 ;
        RECT -76.015 -264.185 46.025 -263.235 ;
        RECT -143.200 -264.460 -141.200 -264.230 ;
        RECT -143.200 -265.050 -141.200 -264.820 ;
        RECT -143.200 -265.640 -141.200 -265.410 ;
        RECT -143.200 -266.230 -141.200 -266.000 ;
        RECT -143.200 -266.820 -141.200 -266.590 ;
        RECT -143.200 -267.410 -141.200 -267.180 ;
        RECT -143.200 -268.000 -141.200 -267.770 ;
        RECT -143.200 -268.590 -141.200 -268.360 ;
        RECT -143.200 -269.180 -141.200 -268.950 ;
        RECT -143.200 -269.770 -141.200 -269.540 ;
        RECT -143.200 -270.360 -141.200 -270.130 ;
        RECT -106.225 -270.430 -105.995 -269.430 ;
        RECT -105.245 -270.430 -105.015 -269.430 ;
        RECT -104.265 -270.430 -104.035 -269.430 ;
        RECT -100.575 -270.430 -100.345 -269.430 ;
        RECT -76.015 -269.630 -75.065 -264.185 ;
        RECT -68.230 -266.495 -68.000 -265.495 ;
        RECT -67.250 -266.495 -67.020 -265.495 ;
        RECT -66.270 -266.495 -66.040 -265.495 ;
        RECT -65.120 -266.760 -64.835 -265.585 ;
        RECT -64.045 -266.495 -63.815 -265.495 ;
        RECT -63.065 -266.495 -62.835 -265.495 ;
        RECT -62.085 -266.495 -61.855 -265.495 ;
        RECT -60.990 -266.070 -60.760 -265.570 ;
        RECT -60.500 -266.070 -60.270 -265.570 ;
        RECT -60.010 -266.070 -59.780 -265.570 ;
        RECT -59.520 -266.070 -59.290 -265.570 ;
        RECT -59.030 -266.070 -58.800 -265.570 ;
        RECT -58.540 -266.070 -58.310 -265.570 ;
        RECT -58.050 -266.070 -57.820 -265.570 ;
        RECT -57.560 -266.070 -57.330 -265.570 ;
        RECT -54.730 -266.495 -54.500 -265.495 ;
        RECT -53.750 -266.495 -53.520 -265.495 ;
        RECT -52.770 -266.495 -52.540 -265.495 ;
        RECT -60.975 -266.760 -60.130 -266.710 ;
        RECT -65.120 -267.045 -60.130 -266.760 ;
        RECT -51.620 -266.760 -51.335 -265.585 ;
        RECT -50.545 -266.495 -50.315 -265.495 ;
        RECT -49.565 -266.495 -49.335 -265.495 ;
        RECT -48.585 -266.495 -48.355 -265.495 ;
        RECT -47.490 -266.070 -47.260 -265.570 ;
        RECT -47.000 -266.070 -46.770 -265.570 ;
        RECT -46.510 -266.070 -46.280 -265.570 ;
        RECT -46.020 -266.070 -45.790 -265.570 ;
        RECT -45.530 -266.070 -45.300 -265.570 ;
        RECT -45.040 -266.070 -44.810 -265.570 ;
        RECT -44.550 -266.070 -44.320 -265.570 ;
        RECT -44.060 -266.070 -43.830 -265.570 ;
        RECT -47.475 -266.760 -46.630 -266.710 ;
        RECT -55.915 -266.870 -55.615 -266.840 ;
        RECT -57.090 -266.975 -56.885 -266.970 ;
        RECT -60.975 -267.080 -60.130 -267.045 ;
        RECT -68.720 -267.895 -68.490 -267.395 ;
        RECT -68.230 -267.895 -68.000 -267.395 ;
        RECT -67.740 -267.895 -67.510 -267.395 ;
        RECT -67.250 -267.895 -67.020 -267.395 ;
        RECT -66.760 -267.895 -66.530 -267.395 ;
        RECT -66.270 -267.895 -66.040 -267.395 ;
        RECT -67.550 -269.010 -66.865 -268.710 ;
        RECT -69.290 -269.300 -68.990 -269.065 ;
        RECT -70.600 -269.620 -68.990 -269.300 ;
        RECT -143.200 -270.950 -141.200 -270.720 ;
        RECT -143.200 -271.540 -141.200 -271.310 ;
        RECT -96.230 -271.540 -96.000 -270.040 ;
        RECT -98.265 -271.815 -97.580 -271.730 ;
        RECT -143.200 -272.130 -141.200 -271.900 ;
        RECT -98.405 -272.020 -97.580 -271.815 ;
        RECT -143.200 -272.720 -141.200 -272.490 ;
        RECT -143.200 -273.310 -141.200 -273.080 ;
        RECT -143.200 -273.900 -141.200 -273.670 ;
        RECT -106.715 -273.965 -106.485 -272.465 ;
        RECT -106.225 -273.965 -105.995 -272.465 ;
        RECT -105.735 -273.965 -105.505 -272.465 ;
        RECT -105.165 -273.970 -104.935 -272.470 ;
        RECT -104.675 -273.970 -104.445 -272.470 ;
        RECT -104.185 -273.970 -103.955 -272.470 ;
        RECT -103.620 -273.970 -103.390 -272.470 ;
        RECT -103.130 -273.970 -102.900 -272.470 ;
        RECT -102.640 -273.970 -102.410 -272.470 ;
        RECT -101.065 -273.970 -100.835 -272.970 ;
        RECT -100.575 -273.550 -100.345 -272.970 ;
        RECT -100.575 -273.725 -98.780 -273.550 ;
        RECT -100.575 -273.970 -100.345 -273.725 ;
        RECT -143.200 -274.490 -141.200 -274.260 ;
        RECT -143.200 -275.080 -141.200 -274.850 ;
        RECT -143.200 -275.670 -141.200 -275.440 ;
        RECT -143.200 -276.260 -141.200 -276.030 ;
        RECT -143.200 -276.850 -141.200 -276.620 ;
        RECT -143.200 -277.440 -141.200 -277.210 ;
        RECT -143.200 -278.030 -141.200 -277.800 ;
        RECT -143.200 -278.620 -141.200 -278.390 ;
        RECT -143.200 -279.210 -141.200 -278.980 ;
        RECT -143.200 -280.390 -141.200 -280.160 ;
        RECT -139.885 -280.910 -139.515 -280.335 ;
        RECT -139.885 -281.140 -137.160 -280.910 ;
        RECT -143.200 -281.570 -141.200 -281.340 ;
        RECT -139.885 -282.090 -139.515 -281.140 ;
        RECT -139.885 -282.320 -137.160 -282.090 ;
        RECT -143.200 -282.750 -141.200 -282.520 ;
        RECT -139.885 -283.270 -139.515 -282.320 ;
        RECT -139.885 -283.500 -137.160 -283.270 ;
        RECT -143.200 -283.930 -141.200 -283.700 ;
        RECT -139.885 -284.450 -139.515 -283.500 ;
        RECT -139.885 -284.680 -137.160 -284.450 ;
        RECT -143.200 -285.110 -141.200 -284.880 ;
        RECT -139.885 -285.630 -139.515 -284.680 ;
        RECT -139.885 -285.860 -137.160 -285.630 ;
        RECT -143.200 -286.290 -141.200 -286.060 ;
        RECT -139.885 -286.810 -139.515 -285.860 ;
        RECT -139.885 -287.040 -137.160 -286.810 ;
        RECT -143.200 -287.470 -141.200 -287.240 ;
        RECT -139.885 -287.990 -139.515 -287.040 ;
        RECT -139.885 -288.220 -137.160 -287.990 ;
        RECT -143.200 -288.650 -141.200 -288.420 ;
        RECT -143.200 -289.205 -140.525 -289.010 ;
        RECT -139.885 -289.170 -139.515 -288.220 ;
        RECT -139.885 -289.205 -137.160 -289.170 ;
        RECT -143.200 -289.240 -137.160 -289.205 ;
        RECT -140.755 -289.400 -137.160 -289.240 ;
        RECT -140.755 -289.435 -139.515 -289.400 ;
        RECT -143.200 -289.830 -141.200 -289.600 ;
        RECT -140.755 -290.190 -140.525 -289.435 ;
        RECT -139.885 -290.060 -139.515 -289.435 ;
        RECT -143.200 -290.420 -140.525 -290.190 ;
        RECT -143.200 -291.010 -141.200 -290.780 ;
        RECT -140.755 -291.370 -140.525 -290.420 ;
        RECT -143.200 -291.600 -140.525 -291.370 ;
        RECT -143.200 -292.190 -141.200 -291.960 ;
        RECT -140.755 -292.550 -140.525 -291.600 ;
        RECT -143.200 -292.780 -140.525 -292.550 ;
        RECT -139.885 -291.000 -139.515 -290.365 ;
        RECT -139.885 -291.230 -137.160 -291.000 ;
        RECT -139.885 -292.180 -139.515 -291.230 ;
        RECT -139.885 -292.410 -137.160 -292.180 ;
        RECT -143.200 -293.370 -141.200 -293.140 ;
        RECT -139.885 -293.360 -139.515 -292.410 ;
        RECT -139.885 -293.590 -137.160 -293.360 ;
        RECT -143.200 -293.960 -140.585 -293.730 ;
        RECT -140.815 -294.115 -140.585 -293.960 ;
        RECT -139.885 -294.115 -139.515 -293.590 ;
        RECT -143.200 -294.550 -141.200 -294.320 ;
        RECT -140.815 -294.345 -139.515 -294.115 ;
        RECT -140.815 -294.910 -140.585 -294.345 ;
        RECT -143.200 -295.140 -140.585 -294.910 ;
        RECT -139.885 -294.540 -139.515 -294.345 ;
        RECT -139.885 -294.770 -137.160 -294.540 ;
        RECT -139.885 -295.415 -139.515 -294.770 ;
        RECT -143.200 -295.730 -141.200 -295.500 ;
        RECT -139.885 -296.090 -139.515 -295.720 ;
        RECT -143.200 -296.320 -139.515 -296.090 ;
        RECT -139.885 -296.370 -139.515 -296.320 ;
        RECT -139.885 -296.600 -137.160 -296.370 ;
        RECT -143.200 -296.910 -141.200 -296.680 ;
        RECT -139.885 -297.550 -139.515 -296.600 ;
        RECT -139.885 -297.780 -137.160 -297.550 ;
        RECT -139.885 -297.805 -139.515 -297.780 ;
        RECT -136.610 -302.970 -134.050 -302.265 ;
        RECT -147.680 -305.245 -134.050 -302.970 ;
        RECT -136.610 -305.390 -134.050 -305.245 ;
        RECT -109.855 -317.995 -109.550 -275.160 ;
        RECT -110.200 -318.000 -109.550 -317.995 ;
        RECT -110.200 -318.165 -109.545 -318.000 ;
        RECT -110.195 -318.590 -109.545 -318.165 ;
        RECT -109.285 -318.635 -108.965 -282.520 ;
        RECT -109.295 -319.495 -108.965 -318.635 ;
        RECT -109.400 -319.500 -108.965 -319.495 ;
        RECT -108.560 -304.875 -108.260 -280.365 ;
        RECT -105.940 -281.085 -105.710 -279.585 ;
        RECT -106.430 -283.765 -106.200 -282.270 ;
        RECT -106.435 -283.950 -106.200 -283.765 ;
        RECT -105.940 -283.770 -105.710 -282.270 ;
        RECT -105.450 -283.950 -105.220 -282.270 ;
        RECT -104.960 -283.770 -104.730 -279.585 ;
        RECT -102.895 -280.360 -102.665 -279.580 ;
        RECT -101.915 -280.350 -101.685 -279.580 ;
        RECT -102.405 -280.360 -101.195 -280.350 ;
        RECT -100.935 -280.360 -100.705 -279.580 ;
        RECT -102.895 -280.590 -99.710 -280.360 ;
        RECT -102.895 -281.235 -102.665 -280.735 ;
        RECT -102.405 -281.235 -102.175 -280.590 ;
        RECT -101.915 -281.235 -101.685 -280.735 ;
        RECT -101.425 -281.235 -101.195 -280.590 ;
        RECT -98.955 -281.395 -98.780 -273.725 ;
        RECT -98.405 -275.570 -98.225 -272.020 ;
        RECT -96.720 -274.220 -96.490 -272.725 ;
        RECT -96.725 -274.405 -96.490 -274.220 ;
        RECT -96.230 -274.225 -96.000 -272.725 ;
        RECT -95.740 -274.405 -95.510 -272.725 ;
        RECT -95.250 -274.225 -95.020 -270.040 ;
        RECT -93.185 -270.815 -92.955 -270.035 ;
        RECT -92.205 -270.805 -91.975 -270.035 ;
        RECT -92.695 -270.815 -91.485 -270.805 ;
        RECT -91.225 -270.815 -90.995 -270.035 ;
        RECT -77.920 -270.195 -74.535 -269.630 ;
        RECT -93.185 -271.045 -90.000 -270.815 ;
        RECT -93.185 -271.690 -92.955 -271.190 ;
        RECT -92.695 -271.690 -92.465 -271.045 ;
        RECT -92.205 -271.690 -91.975 -271.190 ;
        RECT -91.715 -271.690 -91.485 -271.045 ;
        RECT -89.585 -271.170 -88.855 -270.880 ;
        RECT -89.585 -271.300 -89.180 -271.170 ;
        RECT -91.145 -271.475 -89.180 -271.300 ;
        RECT -94.760 -274.405 -94.530 -272.725 ;
        RECT -96.725 -274.640 -94.530 -274.405 ;
        RECT -98.415 -276.230 -98.150 -275.570 ;
        RECT -91.145 -276.825 -90.970 -271.475 ;
        RECT -88.545 -271.985 -86.350 -271.750 ;
        RECT -88.545 -272.170 -88.310 -271.985 ;
        RECT -88.540 -273.665 -88.310 -272.170 ;
        RECT -88.050 -273.665 -87.820 -272.165 ;
        RECT -87.560 -273.665 -87.330 -271.985 ;
        RECT -89.815 -274.145 -88.830 -273.875 ;
        RECT -98.625 -277.000 -90.970 -276.825 ;
        RECT -98.625 -280.740 -98.450 -277.000 ;
        RECT -97.075 -280.110 -96.845 -279.110 ;
        RECT -96.095 -280.110 -95.865 -279.110 ;
        RECT -95.115 -280.110 -94.885 -279.110 ;
        RECT -91.425 -280.110 -91.195 -279.110 ;
        RECT -98.625 -280.970 -98.205 -280.740 ;
        RECT -104.470 -283.950 -104.240 -282.270 ;
        RECT -100.050 -282.565 -99.760 -281.880 ;
        RECT -98.980 -282.080 -98.690 -281.395 ;
        RECT -98.495 -281.425 -98.205 -280.970 ;
        RECT -89.100 -281.165 -88.830 -274.145 ;
        RECT -88.050 -276.350 -87.820 -274.850 ;
        RECT -87.070 -276.350 -86.840 -272.165 ;
        RECT -86.580 -273.665 -86.350 -271.985 ;
        RECT -80.815 -272.235 -80.585 -270.735 ;
        RECT -80.325 -272.235 -80.095 -270.735 ;
        RECT -79.835 -272.235 -79.605 -270.735 ;
        RECT -78.625 -272.235 -78.395 -270.735 ;
        RECT -78.135 -272.235 -77.905 -270.735 ;
        RECT -81.310 -272.725 -76.210 -272.400 ;
        RECT -76.535 -273.140 -76.210 -272.725 ;
        RECT -76.565 -273.500 -76.040 -273.140 ;
        RECT -85.005 -275.200 -84.775 -274.700 ;
        RECT -84.515 -275.345 -84.285 -274.700 ;
        RECT -84.025 -275.200 -83.795 -274.700 ;
        RECT -83.535 -275.345 -83.305 -274.700 ;
        RECT -85.005 -275.575 -81.820 -275.345 ;
        RECT -85.005 -276.355 -84.775 -275.575 ;
        RECT -84.515 -275.585 -83.305 -275.575 ;
        RECT -84.025 -276.355 -83.795 -275.585 ;
        RECT -83.045 -276.355 -82.815 -275.575 ;
        RECT -80.815 -276.795 -80.585 -273.795 ;
        RECT -79.760 -276.795 -79.530 -273.795 ;
        RECT -79.270 -276.795 -79.040 -273.795 ;
        RECT -78.780 -276.795 -78.550 -273.795 ;
        RECT -77.720 -276.795 -77.490 -273.795 ;
        RECT -89.350 -281.915 -88.700 -281.165 ;
        RECT -87.920 -281.275 -87.690 -279.995 ;
        RECT -86.940 -281.265 -86.710 -279.995 ;
        RECT -87.430 -281.275 -86.220 -281.265 ;
        RECT -85.960 -281.275 -85.730 -279.995 ;
        RECT -83.055 -280.850 -82.825 -279.350 ;
        RECT -87.920 -281.505 -84.735 -281.275 ;
        RECT -84.025 -281.370 -83.230 -281.080 ;
        RECT -97.565 -283.645 -97.335 -282.145 ;
        RECT -97.075 -283.645 -96.845 -282.145 ;
        RECT -96.585 -283.645 -96.355 -282.145 ;
        RECT -96.015 -283.650 -95.785 -282.150 ;
        RECT -95.525 -283.650 -95.295 -282.150 ;
        RECT -95.035 -283.650 -94.805 -282.150 ;
        RECT -94.470 -283.650 -94.240 -282.150 ;
        RECT -93.980 -283.650 -93.750 -282.150 ;
        RECT -93.490 -283.650 -93.260 -282.150 ;
        RECT -87.920 -282.645 -87.690 -281.645 ;
        RECT -87.430 -282.645 -87.200 -281.505 ;
        RECT -86.940 -282.645 -86.710 -281.645 ;
        RECT -86.450 -282.645 -86.220 -281.505 ;
        RECT -83.895 -281.645 -83.625 -281.370 ;
        RECT -85.265 -281.915 -83.625 -281.645 ;
        RECT -91.915 -283.650 -91.685 -282.650 ;
        RECT -91.425 -283.650 -91.195 -282.650 ;
        RECT -85.265 -283.365 -84.995 -281.915 ;
        RECT -90.480 -283.635 -84.995 -283.365 ;
        RECT -83.545 -283.530 -83.315 -282.035 ;
        RECT -106.435 -284.185 -104.240 -283.950 ;
        RECT -90.420 -287.205 -89.220 -283.635 ;
        RECT -83.550 -283.715 -83.315 -283.530 ;
        RECT -83.055 -283.535 -82.825 -282.035 ;
        RECT -82.565 -283.715 -82.335 -282.035 ;
        RECT -82.075 -283.535 -81.845 -279.350 ;
        RECT -80.010 -280.125 -79.780 -279.345 ;
        RECT -79.030 -280.115 -78.800 -279.345 ;
        RECT -79.520 -280.125 -78.310 -280.115 ;
        RECT -78.050 -280.125 -77.820 -279.345 ;
        RECT -80.010 -280.355 -76.825 -280.125 ;
        RECT -80.010 -281.000 -79.780 -280.500 ;
        RECT -79.520 -281.000 -79.290 -280.355 ;
        RECT -79.030 -281.000 -78.800 -280.500 ;
        RECT -78.540 -281.000 -78.310 -280.355 ;
        RECT -75.100 -281.175 -74.535 -270.195 ;
        RECT -70.600 -279.200 -70.280 -269.620 ;
        RECT -69.290 -269.750 -68.990 -269.620 ;
        RECT -67.475 -270.100 -67.000 -269.010 ;
        RECT -65.425 -269.600 -65.125 -267.265 ;
        RECT -57.565 -267.275 -56.880 -266.975 ;
        RECT -55.915 -267.170 -55.200 -266.870 ;
        RECT -51.620 -267.045 -46.630 -266.760 ;
        RECT -47.475 -267.080 -46.630 -267.045 ;
        RECT -64.535 -267.895 -64.305 -267.395 ;
        RECT -64.045 -267.895 -63.815 -267.395 ;
        RECT -63.555 -267.895 -63.325 -267.395 ;
        RECT -63.065 -267.895 -62.835 -267.395 ;
        RECT -62.575 -267.895 -62.345 -267.395 ;
        RECT -62.085 -267.895 -61.855 -267.395 ;
        RECT -60.990 -268.145 -60.760 -267.645 ;
        RECT -60.500 -268.145 -60.270 -267.645 ;
        RECT -60.010 -268.145 -59.780 -267.645 ;
        RECT -59.520 -268.145 -59.290 -267.645 ;
        RECT -59.030 -268.145 -58.800 -267.645 ;
        RECT -58.540 -268.145 -58.310 -267.645 ;
        RECT -58.050 -268.145 -57.820 -267.645 ;
        RECT -57.560 -268.145 -57.330 -267.645 ;
        RECT -65.605 -269.900 -64.945 -269.600 ;
        RECT -57.090 -269.700 -56.885 -267.275 ;
        RECT -56.740 -269.455 -56.055 -269.155 ;
        RECT -64.540 -269.940 -56.885 -269.700 ;
        RECT -67.595 -270.400 -66.935 -270.100 ;
        RECT -68.720 -271.185 -68.490 -270.685 ;
        RECT -68.230 -271.185 -68.000 -270.685 ;
        RECT -67.740 -271.185 -67.510 -270.685 ;
        RECT -67.250 -271.185 -67.020 -270.685 ;
        RECT -66.760 -271.185 -66.530 -270.685 ;
        RECT -66.270 -271.185 -66.040 -270.685 ;
        RECT -64.540 -270.710 -64.300 -269.940 ;
        RECT -64.530 -270.935 -64.300 -270.710 ;
        RECT -64.040 -270.935 -63.810 -270.435 ;
        RECT -63.580 -270.530 -63.275 -269.940 ;
        RECT -63.550 -270.935 -63.320 -270.530 ;
        RECT -63.060 -270.935 -62.830 -270.435 ;
        RECT -62.600 -270.540 -62.295 -269.940 ;
        RECT -62.570 -270.935 -62.340 -270.540 ;
        RECT -62.080 -270.935 -61.850 -270.435 ;
        RECT -61.645 -270.530 -61.340 -269.940 ;
        RECT -61.590 -270.935 -61.360 -270.530 ;
        RECT -61.100 -270.935 -60.870 -270.435 ;
        RECT -60.005 -271.185 -59.775 -270.685 ;
        RECT -59.515 -271.185 -59.285 -270.685 ;
        RECT -59.025 -271.185 -58.795 -270.685 ;
        RECT -58.535 -271.185 -58.305 -270.685 ;
        RECT -58.045 -271.185 -57.815 -270.685 ;
        RECT -57.555 -271.185 -57.325 -270.685 ;
        RECT -61.730 -271.535 -60.885 -271.500 ;
        RECT -61.730 -271.820 -56.740 -271.535 ;
        RECT -56.495 -271.695 -56.195 -269.455 ;
        RECT -55.915 -270.910 -55.615 -267.170 ;
        RECT -44.120 -267.285 -43.350 -266.985 ;
        RECT -55.220 -267.895 -54.990 -267.395 ;
        RECT -54.730 -267.895 -54.500 -267.395 ;
        RECT -54.240 -267.895 -54.010 -267.395 ;
        RECT -53.750 -267.895 -53.520 -267.395 ;
        RECT -53.260 -267.895 -53.030 -267.395 ;
        RECT -52.770 -267.895 -52.540 -267.395 ;
        RECT -54.565 -269.040 -53.880 -268.740 ;
        RECT -54.510 -270.080 -54.035 -269.040 ;
        RECT -51.865 -269.160 -51.565 -267.340 ;
        RECT -51.035 -267.895 -50.805 -267.395 ;
        RECT -50.545 -267.895 -50.315 -267.395 ;
        RECT -50.055 -267.895 -49.825 -267.395 ;
        RECT -49.565 -267.895 -49.335 -267.395 ;
        RECT -49.075 -267.895 -48.845 -267.395 ;
        RECT -48.585 -267.895 -48.355 -267.395 ;
        RECT -47.490 -268.145 -47.260 -267.645 ;
        RECT -47.000 -268.145 -46.770 -267.645 ;
        RECT -46.510 -268.145 -46.280 -267.645 ;
        RECT -46.020 -268.145 -45.790 -267.645 ;
        RECT -45.530 -268.145 -45.300 -267.645 ;
        RECT -45.040 -268.145 -44.810 -267.645 ;
        RECT -44.550 -268.145 -44.320 -267.645 ;
        RECT -44.060 -268.145 -43.830 -267.645 ;
        RECT -43.580 -268.660 -43.350 -267.285 ;
        RECT -47.445 -268.885 -43.350 -268.660 ;
        RECT -47.445 -268.890 -43.390 -268.885 ;
        RECT -52.010 -269.460 -51.350 -269.160 ;
        RECT -47.445 -269.720 -47.215 -268.890 ;
        RECT -41.375 -269.040 -40.715 -268.740 ;
        RECT -41.290 -269.365 -40.815 -269.040 ;
        RECT -38.615 -269.365 -38.140 -264.185 ;
        RECT -37.400 -268.545 -37.170 -265.545 ;
        RECT -36.340 -268.545 -36.110 -265.545 ;
        RECT -35.850 -268.545 -35.620 -265.545 ;
        RECT -35.360 -268.545 -35.130 -265.545 ;
        RECT -34.305 -268.545 -34.075 -265.545 ;
        RECT -30.250 -267.525 -30.020 -266.525 ;
        RECT -29.760 -267.525 -29.530 -266.525 ;
        RECT -29.270 -267.525 -29.040 -266.525 ;
        RECT -28.670 -267.525 -28.440 -266.525 ;
        RECT -28.180 -267.525 -27.950 -266.525 ;
        RECT -27.690 -267.525 -27.460 -266.525 ;
        RECT -25.880 -267.525 -25.650 -266.525 ;
        RECT -24.900 -267.525 -24.670 -266.525 ;
        RECT -23.350 -267.525 -23.120 -266.525 ;
        RECT -21.805 -267.525 -21.575 -266.525 ;
        RECT -17.750 -267.525 -17.520 -266.525 ;
        RECT -17.260 -267.525 -17.030 -266.525 ;
        RECT -16.770 -267.525 -16.540 -266.525 ;
        RECT -16.170 -267.525 -15.940 -266.525 ;
        RECT -15.680 -267.525 -15.450 -266.525 ;
        RECT -15.190 -267.525 -14.960 -266.525 ;
        RECT -13.380 -267.525 -13.150 -266.525 ;
        RECT -12.400 -267.525 -12.170 -266.525 ;
        RECT -10.850 -267.525 -10.620 -266.525 ;
        RECT -9.305 -267.525 -9.075 -266.525 ;
        RECT -5.250 -267.525 -5.020 -266.525 ;
        RECT -4.760 -267.525 -4.530 -266.525 ;
        RECT -4.270 -267.525 -4.040 -266.525 ;
        RECT -3.670 -267.525 -3.440 -266.525 ;
        RECT -3.180 -267.525 -2.950 -266.525 ;
        RECT -2.690 -267.525 -2.460 -266.525 ;
        RECT -0.880 -267.525 -0.650 -266.525 ;
        RECT 0.100 -267.525 0.330 -266.525 ;
        RECT 1.650 -267.525 1.880 -266.525 ;
        RECT 3.195 -267.525 3.425 -266.525 ;
        RECT 7.250 -267.525 7.480 -266.525 ;
        RECT 7.740 -267.525 7.970 -266.525 ;
        RECT 8.230 -267.525 8.460 -266.525 ;
        RECT 8.830 -267.525 9.060 -266.525 ;
        RECT 9.320 -267.525 9.550 -266.525 ;
        RECT 9.810 -267.525 10.040 -266.525 ;
        RECT 11.620 -267.525 11.850 -266.525 ;
        RECT 12.600 -267.525 12.830 -266.525 ;
        RECT 14.150 -267.525 14.380 -266.525 ;
        RECT 15.695 -267.525 15.925 -266.525 ;
        RECT 19.750 -267.525 19.980 -266.525 ;
        RECT 20.240 -267.525 20.470 -266.525 ;
        RECT 20.730 -267.525 20.960 -266.525 ;
        RECT 21.330 -267.525 21.560 -266.525 ;
        RECT 21.820 -267.525 22.050 -266.525 ;
        RECT 22.310 -267.525 22.540 -266.525 ;
        RECT 24.120 -267.525 24.350 -266.525 ;
        RECT 25.100 -267.525 25.330 -266.525 ;
        RECT 26.650 -267.525 26.880 -266.525 ;
        RECT 28.195 -267.525 28.425 -266.525 ;
        RECT 34.750 -267.525 34.980 -266.525 ;
        RECT 35.240 -267.525 35.470 -266.525 ;
        RECT 35.730 -267.525 35.960 -266.525 ;
        RECT 36.330 -267.525 36.560 -266.525 ;
        RECT 36.820 -267.525 37.050 -266.525 ;
        RECT 37.310 -267.525 37.540 -266.525 ;
        RECT 39.120 -267.525 39.350 -266.525 ;
        RECT 40.100 -267.525 40.330 -266.525 ;
        RECT 41.650 -267.525 41.880 -266.525 ;
        RECT 43.195 -267.525 43.425 -266.525 ;
        RECT -24.435 -268.165 -23.740 -268.075 ;
        RECT -21.360 -268.165 -20.665 -268.105 ;
        RECT -11.935 -268.165 -11.240 -268.075 ;
        RECT -8.860 -268.165 -8.165 -268.105 ;
        RECT 0.565 -268.165 1.260 -268.075 ;
        RECT 3.640 -268.165 4.335 -268.105 ;
        RECT 13.065 -268.165 13.760 -268.075 ;
        RECT 16.140 -268.165 16.835 -268.105 ;
        RECT 25.565 -268.165 26.260 -268.075 ;
        RECT 28.640 -268.165 29.335 -268.105 ;
        RECT 40.565 -268.165 41.260 -268.075 ;
        RECT 43.640 -268.165 44.335 -268.105 ;
        RECT 47.145 -268.165 48.145 -266.405 ;
        RECT -30.225 -268.360 -29.530 -268.295 ;
        RECT -24.435 -268.305 -19.910 -268.165 ;
        RECT -24.435 -268.345 -23.740 -268.305 ;
        RECT -30.225 -268.500 -28.455 -268.360 ;
        RECT -21.360 -268.375 -20.665 -268.305 ;
        RECT -30.225 -268.565 -29.530 -268.500 ;
        RECT -51.015 -269.950 -47.215 -269.720 ;
        RECT -42.990 -269.890 -42.330 -269.590 ;
        RECT -41.290 -269.840 -38.140 -269.365 ;
        RECT -54.600 -270.380 -53.915 -270.080 ;
        RECT -51.015 -270.435 -50.785 -269.950 ;
        RECT -50.040 -270.435 -49.830 -269.950 ;
        RECT -49.065 -270.435 -48.855 -269.950 ;
        RECT -48.085 -270.435 -47.875 -269.950 ;
        RECT -55.920 -271.135 -55.615 -270.910 ;
        RECT -55.920 -271.570 -55.620 -271.135 ;
        RECT -55.220 -271.185 -54.990 -270.685 ;
        RECT -54.730 -271.185 -54.500 -270.685 ;
        RECT -54.240 -271.185 -54.010 -270.685 ;
        RECT -53.750 -271.185 -53.520 -270.685 ;
        RECT -53.260 -271.185 -53.030 -270.685 ;
        RECT -52.770 -271.185 -52.540 -270.685 ;
        RECT -51.030 -270.935 -50.785 -270.435 ;
        RECT -50.540 -270.935 -50.310 -270.435 ;
        RECT -50.050 -270.935 -49.820 -270.435 ;
        RECT -49.560 -270.935 -49.330 -270.435 ;
        RECT -49.070 -270.935 -48.840 -270.435 ;
        RECT -48.580 -270.935 -48.350 -270.435 ;
        RECT -48.090 -270.935 -47.860 -270.435 ;
        RECT -47.600 -270.935 -47.370 -270.435 ;
        RECT -46.505 -271.185 -46.275 -270.685 ;
        RECT -46.015 -271.185 -45.785 -270.685 ;
        RECT -45.525 -271.185 -45.295 -270.685 ;
        RECT -45.035 -271.185 -44.805 -270.685 ;
        RECT -44.545 -271.185 -44.315 -270.685 ;
        RECT -44.055 -271.185 -43.825 -270.685 ;
        RECT -42.825 -271.030 -42.535 -269.890 ;
        RECT -41.290 -270.085 -40.815 -269.840 ;
        RECT -41.465 -270.385 -40.780 -270.085 ;
        RECT -48.230 -271.535 -47.385 -271.500 ;
        RECT -61.730 -271.870 -60.885 -271.820 ;
        RECT -68.720 -273.085 -68.490 -272.085 ;
        RECT -67.740 -273.085 -67.510 -272.085 ;
        RECT -66.760 -273.085 -66.530 -272.085 ;
        RECT -64.530 -272.850 -64.300 -272.510 ;
        RECT -64.530 -273.010 -64.275 -272.850 ;
        RECT -64.040 -273.010 -63.810 -272.510 ;
        RECT -63.550 -272.725 -63.320 -272.510 ;
        RECT -64.525 -273.425 -64.275 -273.010 ;
        RECT -63.570 -273.425 -63.315 -272.725 ;
        RECT -63.060 -273.010 -62.830 -272.510 ;
        RECT -62.570 -272.820 -62.340 -272.510 ;
        RECT -62.570 -273.425 -62.315 -272.820 ;
        RECT -62.080 -273.010 -61.850 -272.510 ;
        RECT -61.590 -272.820 -61.360 -272.510 ;
        RECT -61.600 -273.425 -61.345 -272.820 ;
        RECT -61.100 -273.010 -60.870 -272.510 ;
        RECT -60.005 -273.085 -59.775 -272.085 ;
        RECT -59.025 -273.085 -58.795 -272.085 ;
        RECT -58.045 -273.085 -57.815 -272.085 ;
        RECT -57.025 -272.995 -56.740 -271.820 ;
        RECT -48.230 -271.820 -43.240 -271.535 ;
        RECT -42.835 -271.690 -42.535 -271.030 ;
        RECT -42.095 -271.185 -41.865 -270.685 ;
        RECT -41.605 -271.185 -41.375 -270.685 ;
        RECT -41.115 -271.185 -40.885 -270.685 ;
        RECT -40.625 -271.185 -40.395 -270.685 ;
        RECT -40.135 -271.185 -39.905 -270.685 ;
        RECT -39.645 -271.185 -39.415 -270.685 ;
        RECT -48.230 -271.870 -47.385 -271.820 ;
        RECT -55.220 -273.085 -54.990 -272.085 ;
        RECT -54.240 -273.085 -54.010 -272.085 ;
        RECT -53.260 -273.085 -53.030 -272.085 ;
        RECT -51.030 -273.010 -50.800 -272.510 ;
        RECT -50.540 -273.010 -50.310 -272.510 ;
        RECT -50.050 -273.010 -49.820 -272.510 ;
        RECT -49.560 -273.010 -49.330 -272.510 ;
        RECT -49.070 -273.010 -48.840 -272.510 ;
        RECT -48.580 -273.010 -48.350 -272.510 ;
        RECT -48.090 -273.010 -47.860 -272.510 ;
        RECT -47.600 -273.010 -47.370 -272.510 ;
        RECT -46.505 -273.085 -46.275 -272.085 ;
        RECT -45.525 -273.085 -45.295 -272.085 ;
        RECT -44.545 -273.085 -44.315 -272.085 ;
        RECT -43.525 -273.425 -43.240 -271.820 ;
        RECT -42.095 -273.085 -41.865 -272.085 ;
        RECT -41.115 -273.085 -40.885 -272.085 ;
        RECT -40.135 -273.085 -39.905 -272.085 ;
        RECT -64.525 -273.710 -43.240 -273.425 ;
        RECT -38.615 -274.510 -38.140 -269.840 ;
        RECT -36.985 -271.605 -36.755 -270.105 ;
        RECT -36.495 -271.605 -36.265 -270.105 ;
        RECT -35.285 -271.605 -35.055 -270.105 ;
        RECT -34.795 -271.605 -34.565 -270.105 ;
        RECT -34.305 -271.605 -34.075 -270.105 ;
        RECT -52.975 -275.075 -38.135 -274.510 ;
        RECT -63.600 -276.865 -61.405 -276.630 ;
        RECT -63.600 -277.050 -63.365 -276.865 ;
        RECT -63.595 -278.545 -63.365 -277.050 ;
        RECT -63.105 -278.545 -62.875 -277.045 ;
        RECT -62.615 -278.545 -62.385 -276.865 ;
        RECT -66.290 -279.200 -65.360 -278.990 ;
        RECT -70.600 -279.520 -65.360 -279.200 ;
        RECT -66.290 -279.760 -65.360 -279.520 ;
        RECT -78.075 -281.740 -74.535 -281.175 ;
        RECT -63.105 -281.230 -62.875 -279.730 ;
        RECT -62.125 -281.230 -61.895 -277.045 ;
        RECT -61.635 -278.545 -61.405 -276.865 ;
        RECT -55.870 -277.115 -55.640 -275.615 ;
        RECT -55.380 -277.115 -55.150 -275.615 ;
        RECT -54.890 -277.115 -54.660 -275.615 ;
        RECT -53.680 -277.115 -53.450 -275.615 ;
        RECT -53.190 -277.115 -52.960 -275.615 ;
        RECT -56.365 -277.605 -51.265 -277.280 ;
        RECT -51.590 -278.020 -51.265 -277.605 ;
        RECT -51.620 -278.380 -51.095 -278.020 ;
        RECT -60.060 -280.080 -59.830 -279.580 ;
        RECT -59.570 -280.225 -59.340 -279.580 ;
        RECT -59.080 -280.080 -58.850 -279.580 ;
        RECT -58.590 -280.225 -58.360 -279.580 ;
        RECT -60.060 -280.455 -56.875 -280.225 ;
        RECT -60.060 -281.235 -59.830 -280.455 ;
        RECT -59.570 -280.465 -58.360 -280.455 ;
        RECT -59.080 -281.235 -58.850 -280.465 ;
        RECT -58.100 -281.235 -57.870 -280.455 ;
        RECT -55.870 -281.675 -55.640 -278.675 ;
        RECT -54.815 -281.675 -54.585 -278.675 ;
        RECT -54.325 -281.675 -54.095 -278.675 ;
        RECT -53.835 -281.675 -53.605 -278.675 ;
        RECT -52.775 -281.675 -52.545 -278.675 ;
        RECT -81.585 -283.715 -81.355 -282.035 ;
        RECT -83.550 -283.950 -81.355 -283.715 ;
        RECT -78.490 -285.495 -77.150 -284.170 ;
        RECT -78.245 -288.270 -77.305 -285.495 ;
        RECT -78.465 -289.595 -77.125 -288.270 ;
        RECT -75.100 -294.630 -74.535 -281.740 ;
        RECT -62.975 -286.155 -62.745 -284.875 ;
        RECT -61.995 -286.145 -61.765 -284.875 ;
        RECT -62.485 -286.155 -61.275 -286.145 ;
        RECT -61.015 -286.155 -60.785 -284.875 ;
        RECT -58.110 -285.730 -57.880 -284.230 ;
        RECT -77.920 -295.195 -74.535 -294.630 ;
        RECT -105.615 -298.555 -105.385 -295.555 ;
        RECT -104.555 -298.555 -104.325 -295.555 ;
        RECT -104.065 -298.555 -103.835 -295.555 ;
        RECT -103.575 -298.555 -103.345 -295.555 ;
        RECT -103.010 -298.555 -102.780 -295.555 ;
        RECT -102.520 -298.555 -102.290 -295.555 ;
        RECT -102.030 -298.555 -101.800 -295.555 ;
        RECT -99.585 -297.200 -99.355 -295.200 ;
        RECT -98.530 -297.200 -98.300 -295.200 ;
        RECT -98.040 -297.200 -97.810 -295.200 ;
        RECT -97.550 -297.200 -97.320 -295.200 ;
        RECT -95.060 -297.205 -94.830 -295.205 ;
        RECT -94.005 -297.205 -93.775 -295.205 ;
        RECT -93.515 -297.205 -93.285 -295.205 ;
        RECT -93.025 -297.205 -92.795 -295.205 ;
        RECT -88.545 -296.985 -86.350 -296.750 ;
        RECT -88.545 -297.170 -88.310 -296.985 ;
        RECT -96.365 -298.015 -96.075 -297.330 ;
        RECT -100.570 -298.200 -100.280 -298.180 ;
        RECT -100.575 -298.865 -100.280 -298.200 ;
        RECT -97.490 -298.440 -96.805 -298.150 ;
        RECT -101.925 -300.185 -101.240 -299.895 ;
        RECT -105.615 -301.375 -105.385 -300.375 ;
        RECT -105.125 -301.375 -104.895 -300.375 ;
        RECT -104.635 -301.375 -104.405 -300.375 ;
        RECT -104.145 -301.375 -103.915 -300.375 ;
        RECT -106.285 -302.605 -102.265 -301.855 ;
        RECT -106.225 -304.665 -105.790 -302.605 ;
        RECT -105.325 -304.665 -104.890 -302.605 ;
        RECT -104.460 -304.665 -104.025 -302.605 ;
        RECT -103.540 -304.665 -103.105 -302.605 ;
        RECT -102.915 -304.665 -102.480 -302.605 ;
        RECT -107.350 -304.875 -102.435 -304.665 ;
        RECT -108.560 -305.175 -102.435 -304.875 ;
        RECT -109.400 -320.115 -108.785 -319.500 ;
        RECT -108.560 -321.335 -108.260 -305.175 ;
        RECT -107.350 -305.240 -102.435 -305.175 ;
        RECT -101.865 -305.175 -101.415 -300.185 ;
        RECT -100.575 -302.950 -100.360 -298.865 ;
        RECT -99.585 -299.660 -99.355 -298.660 ;
        RECT -99.095 -299.660 -98.865 -298.660 ;
        RECT -98.605 -299.660 -98.375 -298.660 ;
        RECT -100.580 -303.635 -100.290 -302.950 ;
        RECT -101.865 -305.625 -100.280 -305.175 ;
        RECT -107.300 -307.105 -107.070 -306.105 ;
        RECT -106.810 -307.105 -106.580 -306.105 ;
        RECT -105.235 -307.605 -105.005 -306.105 ;
        RECT -104.745 -307.605 -104.515 -306.105 ;
        RECT -104.255 -307.605 -104.025 -306.105 ;
        RECT -103.690 -307.605 -103.460 -306.105 ;
        RECT -103.200 -307.605 -102.970 -306.105 ;
        RECT -102.710 -307.605 -102.480 -306.105 ;
        RECT -102.140 -307.610 -101.910 -306.110 ;
        RECT -101.650 -307.610 -101.420 -306.110 ;
        RECT -101.160 -307.610 -100.930 -306.110 ;
        RECT -100.730 -308.565 -100.280 -305.625 ;
        RECT -97.035 -308.290 -96.860 -298.440 ;
        RECT -96.365 -303.345 -96.190 -298.015 ;
        RECT -95.980 -298.875 -95.690 -298.190 ;
        RECT -92.835 -298.445 -92.150 -298.155 ;
        RECT -96.475 -304.030 -96.185 -303.345 ;
        RECT -95.980 -303.730 -95.805 -298.875 ;
        RECT -95.060 -299.665 -94.830 -298.665 ;
        RECT -94.570 -299.665 -94.340 -298.665 ;
        RECT -94.080 -299.665 -93.850 -298.665 ;
        RECT -96.010 -304.415 -95.720 -303.730 ;
        RECT -97.075 -308.975 -96.785 -308.290 ;
        RECT -92.410 -308.720 -92.235 -298.445 ;
        RECT -88.540 -298.665 -88.310 -297.170 ;
        RECT -88.050 -298.665 -87.820 -297.165 ;
        RECT -87.560 -298.665 -87.330 -296.985 ;
        RECT -89.815 -299.145 -88.830 -298.875 ;
        RECT -91.530 -299.935 -90.945 -299.320 ;
        RECT -92.025 -306.960 -91.735 -306.275 ;
        RECT -92.450 -309.405 -92.160 -308.720 ;
        RECT -107.300 -310.645 -107.070 -309.645 ;
        RECT -103.610 -310.645 -103.380 -309.645 ;
        RECT -102.630 -310.645 -102.400 -309.645 ;
        RECT -101.650 -310.645 -101.420 -309.645 ;
        RECT -107.295 -312.000 -107.080 -310.645 ;
        RECT -107.545 -312.580 -106.755 -312.000 ;
        RECT -92.020 -312.140 -91.825 -306.960 ;
        RECT -91.515 -311.255 -91.055 -299.935 ;
        RECT -89.100 -306.165 -88.830 -299.145 ;
        RECT -88.050 -301.350 -87.820 -299.850 ;
        RECT -87.070 -301.350 -86.840 -297.165 ;
        RECT -86.580 -298.665 -86.350 -296.985 ;
        RECT -80.815 -297.235 -80.585 -295.735 ;
        RECT -80.325 -297.235 -80.095 -295.735 ;
        RECT -79.835 -297.235 -79.605 -295.735 ;
        RECT -78.625 -297.235 -78.395 -295.735 ;
        RECT -78.135 -297.235 -77.905 -295.735 ;
        RECT -81.310 -297.725 -76.210 -297.400 ;
        RECT -76.535 -298.140 -76.210 -297.725 ;
        RECT -76.565 -298.500 -76.040 -298.140 ;
        RECT -85.005 -300.200 -84.775 -299.700 ;
        RECT -84.515 -300.345 -84.285 -299.700 ;
        RECT -84.025 -300.200 -83.795 -299.700 ;
        RECT -83.535 -300.345 -83.305 -299.700 ;
        RECT -85.005 -300.575 -81.820 -300.345 ;
        RECT -85.005 -301.355 -84.775 -300.575 ;
        RECT -84.515 -300.585 -83.305 -300.575 ;
        RECT -84.025 -301.355 -83.795 -300.585 ;
        RECT -83.045 -301.355 -82.815 -300.575 ;
        RECT -80.815 -301.795 -80.585 -298.795 ;
        RECT -79.760 -301.795 -79.530 -298.795 ;
        RECT -79.270 -301.795 -79.040 -298.795 ;
        RECT -78.780 -301.795 -78.550 -298.795 ;
        RECT -77.720 -301.795 -77.490 -298.795 ;
        RECT -89.350 -306.915 -88.700 -306.165 ;
        RECT -87.920 -306.275 -87.690 -304.995 ;
        RECT -86.940 -306.265 -86.710 -304.995 ;
        RECT -87.430 -306.275 -86.220 -306.265 ;
        RECT -85.960 -306.275 -85.730 -304.995 ;
        RECT -83.055 -305.850 -82.825 -304.350 ;
        RECT -87.920 -306.505 -84.735 -306.275 ;
        RECT -84.025 -306.370 -83.230 -306.080 ;
        RECT -87.920 -307.645 -87.690 -306.645 ;
        RECT -87.430 -307.645 -87.200 -306.505 ;
        RECT -86.940 -307.645 -86.710 -306.645 ;
        RECT -86.450 -307.645 -86.220 -306.505 ;
        RECT -83.895 -306.645 -83.625 -306.370 ;
        RECT -85.265 -306.915 -83.625 -306.645 ;
        RECT -85.265 -308.365 -84.995 -306.915 ;
        RECT -90.480 -308.635 -84.995 -308.365 ;
        RECT -83.545 -308.530 -83.315 -307.035 ;
        RECT -90.480 -309.985 -90.210 -308.635 ;
        RECT -83.550 -308.715 -83.315 -308.530 ;
        RECT -83.055 -308.535 -82.825 -307.035 ;
        RECT -82.565 -308.715 -82.335 -307.035 ;
        RECT -82.075 -308.535 -81.845 -304.350 ;
        RECT -80.010 -305.125 -79.780 -304.345 ;
        RECT -79.030 -305.115 -78.800 -304.345 ;
        RECT -79.520 -305.125 -78.310 -305.115 ;
        RECT -78.050 -305.125 -77.820 -304.345 ;
        RECT -80.010 -305.355 -76.825 -305.125 ;
        RECT -80.010 -306.000 -79.780 -305.500 ;
        RECT -79.520 -306.000 -79.290 -305.355 ;
        RECT -79.030 -306.000 -78.800 -305.500 ;
        RECT -78.540 -306.000 -78.310 -305.355 ;
        RECT -75.100 -306.175 -74.535 -295.195 ;
        RECT -73.770 -298.155 -72.730 -286.175 ;
        RECT -62.975 -286.385 -59.790 -286.155 ;
        RECT -59.080 -286.250 -58.285 -285.960 ;
        RECT -62.975 -287.525 -62.745 -286.525 ;
        RECT -62.485 -287.525 -62.255 -286.385 ;
        RECT -61.995 -287.525 -61.765 -286.525 ;
        RECT -61.505 -287.525 -61.275 -286.385 ;
        RECT -58.950 -286.525 -58.680 -286.250 ;
        RECT -60.320 -286.795 -58.680 -286.525 ;
        RECT -60.320 -288.245 -60.050 -286.795 ;
        RECT -70.890 -288.515 -60.050 -288.245 ;
        RECT -58.600 -288.410 -58.370 -286.915 ;
        RECT -70.890 -293.935 -70.620 -288.515 ;
        RECT -58.605 -288.595 -58.370 -288.410 ;
        RECT -58.110 -288.415 -57.880 -286.915 ;
        RECT -57.620 -288.595 -57.390 -286.915 ;
        RECT -57.130 -288.415 -56.900 -284.230 ;
        RECT -55.065 -285.005 -54.835 -284.225 ;
        RECT -54.085 -284.995 -53.855 -284.225 ;
        RECT -54.575 -285.005 -53.365 -284.995 ;
        RECT -53.105 -285.005 -52.875 -284.225 ;
        RECT -55.065 -285.235 -51.880 -285.005 ;
        RECT -55.065 -285.880 -54.835 -285.380 ;
        RECT -54.575 -285.880 -54.345 -285.235 ;
        RECT -54.085 -285.880 -53.855 -285.380 ;
        RECT -53.595 -285.880 -53.365 -285.235 ;
        RECT -50.155 -286.055 -49.590 -275.075 ;
        RECT -53.130 -286.620 -49.590 -286.055 ;
        RECT -56.640 -288.595 -56.410 -286.915 ;
        RECT -58.605 -288.830 -56.410 -288.595 ;
        RECT -68.230 -291.130 -68.000 -290.130 ;
        RECT -67.250 -291.130 -67.020 -290.130 ;
        RECT -66.270 -291.130 -66.040 -290.130 ;
        RECT -65.120 -291.395 -64.835 -290.220 ;
        RECT -64.045 -291.130 -63.815 -290.130 ;
        RECT -63.065 -291.130 -62.835 -290.130 ;
        RECT -62.085 -291.130 -61.855 -290.130 ;
        RECT -60.990 -290.705 -60.760 -290.205 ;
        RECT -60.500 -290.705 -60.270 -290.205 ;
        RECT -60.010 -290.705 -59.780 -290.205 ;
        RECT -59.520 -290.705 -59.290 -290.205 ;
        RECT -59.030 -290.705 -58.800 -290.205 ;
        RECT -58.540 -290.705 -58.310 -290.205 ;
        RECT -58.050 -290.705 -57.820 -290.205 ;
        RECT -57.560 -290.705 -57.330 -290.205 ;
        RECT -54.730 -291.130 -54.500 -290.130 ;
        RECT -53.750 -291.130 -53.520 -290.130 ;
        RECT -52.770 -291.130 -52.540 -290.130 ;
        RECT -60.975 -291.395 -60.130 -291.345 ;
        RECT -65.120 -291.680 -60.130 -291.395 ;
        RECT -51.620 -291.395 -51.335 -290.220 ;
        RECT -50.545 -291.130 -50.315 -290.130 ;
        RECT -49.565 -291.130 -49.335 -290.130 ;
        RECT -48.585 -291.130 -48.355 -290.130 ;
        RECT -47.490 -290.705 -47.260 -290.205 ;
        RECT -47.000 -290.705 -46.770 -290.205 ;
        RECT -46.510 -290.705 -46.280 -290.205 ;
        RECT -46.020 -290.705 -45.790 -290.205 ;
        RECT -45.530 -290.705 -45.300 -290.205 ;
        RECT -45.040 -290.705 -44.810 -290.205 ;
        RECT -44.550 -290.705 -44.320 -290.205 ;
        RECT -44.060 -290.705 -43.830 -290.205 ;
        RECT -47.475 -291.395 -46.630 -291.345 ;
        RECT -55.915 -291.505 -55.615 -291.475 ;
        RECT -57.090 -291.610 -56.885 -291.605 ;
        RECT -60.975 -291.715 -60.130 -291.680 ;
        RECT -68.720 -292.530 -68.490 -292.030 ;
        RECT -68.230 -292.530 -68.000 -292.030 ;
        RECT -67.740 -292.530 -67.510 -292.030 ;
        RECT -67.250 -292.530 -67.020 -292.030 ;
        RECT -66.760 -292.530 -66.530 -292.030 ;
        RECT -66.270 -292.530 -66.040 -292.030 ;
        RECT -67.550 -293.645 -66.865 -293.345 ;
        RECT -69.290 -293.935 -68.990 -293.700 ;
        RECT -70.890 -294.255 -68.990 -293.935 ;
        RECT -69.290 -294.385 -68.990 -294.255 ;
        RECT -67.475 -294.735 -67.000 -293.645 ;
        RECT -65.425 -294.235 -65.125 -291.900 ;
        RECT -57.565 -291.910 -56.880 -291.610 ;
        RECT -55.915 -291.805 -55.200 -291.505 ;
        RECT -51.620 -291.680 -46.630 -291.395 ;
        RECT -47.475 -291.715 -46.630 -291.680 ;
        RECT -64.535 -292.530 -64.305 -292.030 ;
        RECT -64.045 -292.530 -63.815 -292.030 ;
        RECT -63.555 -292.530 -63.325 -292.030 ;
        RECT -63.065 -292.530 -62.835 -292.030 ;
        RECT -62.575 -292.530 -62.345 -292.030 ;
        RECT -62.085 -292.530 -61.855 -292.030 ;
        RECT -60.990 -292.780 -60.760 -292.280 ;
        RECT -60.500 -292.780 -60.270 -292.280 ;
        RECT -60.010 -292.780 -59.780 -292.280 ;
        RECT -59.520 -292.780 -59.290 -292.280 ;
        RECT -59.030 -292.780 -58.800 -292.280 ;
        RECT -58.540 -292.780 -58.310 -292.280 ;
        RECT -58.050 -292.780 -57.820 -292.280 ;
        RECT -57.560 -292.780 -57.330 -292.280 ;
        RECT -65.605 -294.535 -64.945 -294.235 ;
        RECT -57.090 -294.335 -56.885 -291.910 ;
        RECT -56.740 -294.090 -56.055 -293.790 ;
        RECT -64.540 -294.575 -56.885 -294.335 ;
        RECT -67.595 -295.035 -66.935 -294.735 ;
        RECT -68.720 -295.820 -68.490 -295.320 ;
        RECT -68.230 -295.820 -68.000 -295.320 ;
        RECT -67.740 -295.820 -67.510 -295.320 ;
        RECT -67.250 -295.820 -67.020 -295.320 ;
        RECT -66.760 -295.820 -66.530 -295.320 ;
        RECT -66.270 -295.820 -66.040 -295.320 ;
        RECT -64.540 -295.345 -64.300 -294.575 ;
        RECT -64.530 -295.570 -64.300 -295.345 ;
        RECT -64.040 -295.570 -63.810 -295.070 ;
        RECT -63.580 -295.165 -63.275 -294.575 ;
        RECT -63.550 -295.570 -63.320 -295.165 ;
        RECT -63.060 -295.570 -62.830 -295.070 ;
        RECT -62.600 -295.175 -62.295 -294.575 ;
        RECT -62.570 -295.570 -62.340 -295.175 ;
        RECT -62.080 -295.570 -61.850 -295.070 ;
        RECT -61.645 -295.165 -61.340 -294.575 ;
        RECT -61.590 -295.570 -61.360 -295.165 ;
        RECT -61.100 -295.570 -60.870 -295.070 ;
        RECT -60.005 -295.820 -59.775 -295.320 ;
        RECT -59.515 -295.820 -59.285 -295.320 ;
        RECT -59.025 -295.820 -58.795 -295.320 ;
        RECT -58.535 -295.820 -58.305 -295.320 ;
        RECT -58.045 -295.820 -57.815 -295.320 ;
        RECT -57.555 -295.820 -57.325 -295.320 ;
        RECT -61.730 -296.170 -60.885 -296.135 ;
        RECT -61.730 -296.455 -56.740 -296.170 ;
        RECT -56.495 -296.330 -56.195 -294.090 ;
        RECT -55.915 -295.545 -55.615 -291.805 ;
        RECT -44.120 -291.920 -43.350 -291.620 ;
        RECT -55.220 -292.530 -54.990 -292.030 ;
        RECT -54.730 -292.530 -54.500 -292.030 ;
        RECT -54.240 -292.530 -54.010 -292.030 ;
        RECT -53.750 -292.530 -53.520 -292.030 ;
        RECT -53.260 -292.530 -53.030 -292.030 ;
        RECT -52.770 -292.530 -52.540 -292.030 ;
        RECT -54.565 -293.675 -53.880 -293.375 ;
        RECT -54.510 -294.715 -54.035 -293.675 ;
        RECT -51.865 -293.795 -51.565 -291.975 ;
        RECT -51.035 -292.530 -50.805 -292.030 ;
        RECT -50.545 -292.530 -50.315 -292.030 ;
        RECT -50.055 -292.530 -49.825 -292.030 ;
        RECT -49.565 -292.530 -49.335 -292.030 ;
        RECT -49.075 -292.530 -48.845 -292.030 ;
        RECT -48.585 -292.530 -48.355 -292.030 ;
        RECT -47.490 -292.780 -47.260 -292.280 ;
        RECT -47.000 -292.780 -46.770 -292.280 ;
        RECT -46.510 -292.780 -46.280 -292.280 ;
        RECT -46.020 -292.780 -45.790 -292.280 ;
        RECT -45.530 -292.780 -45.300 -292.280 ;
        RECT -45.040 -292.780 -44.810 -292.280 ;
        RECT -44.550 -292.780 -44.320 -292.280 ;
        RECT -44.060 -292.780 -43.830 -292.280 ;
        RECT -43.580 -293.295 -43.350 -291.920 ;
        RECT -47.445 -293.520 -43.350 -293.295 ;
        RECT -41.290 -293.375 -40.815 -275.075 ;
        RECT -47.445 -293.525 -43.390 -293.520 ;
        RECT -52.010 -294.095 -51.350 -293.795 ;
        RECT -47.445 -294.355 -47.215 -293.525 ;
        RECT -41.375 -293.675 -40.715 -293.375 ;
        RECT -51.015 -294.585 -47.215 -294.355 ;
        RECT -42.990 -294.525 -42.330 -294.225 ;
        RECT -54.600 -295.015 -53.915 -294.715 ;
        RECT -51.015 -295.070 -50.785 -294.585 ;
        RECT -50.040 -295.070 -49.830 -294.585 ;
        RECT -49.065 -295.070 -48.855 -294.585 ;
        RECT -48.085 -295.070 -47.875 -294.585 ;
        RECT -55.920 -295.770 -55.615 -295.545 ;
        RECT -55.920 -296.205 -55.620 -295.770 ;
        RECT -55.220 -295.820 -54.990 -295.320 ;
        RECT -54.730 -295.820 -54.500 -295.320 ;
        RECT -54.240 -295.820 -54.010 -295.320 ;
        RECT -53.750 -295.820 -53.520 -295.320 ;
        RECT -53.260 -295.820 -53.030 -295.320 ;
        RECT -52.770 -295.820 -52.540 -295.320 ;
        RECT -51.030 -295.570 -50.785 -295.070 ;
        RECT -50.540 -295.570 -50.310 -295.070 ;
        RECT -50.050 -295.570 -49.820 -295.070 ;
        RECT -49.560 -295.570 -49.330 -295.070 ;
        RECT -49.070 -295.570 -48.840 -295.070 ;
        RECT -48.580 -295.570 -48.350 -295.070 ;
        RECT -48.090 -295.570 -47.860 -295.070 ;
        RECT -47.600 -295.570 -47.370 -295.070 ;
        RECT -46.505 -295.820 -46.275 -295.320 ;
        RECT -46.015 -295.820 -45.785 -295.320 ;
        RECT -45.525 -295.820 -45.295 -295.320 ;
        RECT -45.035 -295.820 -44.805 -295.320 ;
        RECT -44.545 -295.820 -44.315 -295.320 ;
        RECT -44.055 -295.820 -43.825 -295.320 ;
        RECT -42.825 -295.665 -42.535 -294.525 ;
        RECT -41.290 -294.720 -40.815 -293.675 ;
        RECT -41.465 -295.020 -40.780 -294.720 ;
        RECT -48.230 -296.170 -47.385 -296.135 ;
        RECT -61.730 -296.505 -60.885 -296.455 ;
        RECT -68.720 -297.720 -68.490 -296.720 ;
        RECT -67.740 -297.720 -67.510 -296.720 ;
        RECT -66.760 -297.720 -66.530 -296.720 ;
        RECT -64.530 -297.485 -64.300 -297.145 ;
        RECT -64.530 -297.645 -64.275 -297.485 ;
        RECT -64.040 -297.645 -63.810 -297.145 ;
        RECT -63.550 -297.360 -63.320 -297.145 ;
        RECT -64.525 -298.060 -64.275 -297.645 ;
        RECT -63.570 -298.060 -63.315 -297.360 ;
        RECT -63.060 -297.645 -62.830 -297.145 ;
        RECT -62.570 -297.455 -62.340 -297.145 ;
        RECT -62.570 -298.060 -62.315 -297.455 ;
        RECT -62.080 -297.645 -61.850 -297.145 ;
        RECT -61.590 -297.455 -61.360 -297.145 ;
        RECT -61.600 -298.060 -61.345 -297.455 ;
        RECT -61.100 -297.645 -60.870 -297.145 ;
        RECT -60.005 -297.720 -59.775 -296.720 ;
        RECT -59.025 -297.720 -58.795 -296.720 ;
        RECT -58.045 -297.720 -57.815 -296.720 ;
        RECT -57.025 -297.630 -56.740 -296.455 ;
        RECT -48.230 -296.455 -43.240 -296.170 ;
        RECT -42.835 -296.325 -42.535 -295.665 ;
        RECT -42.095 -295.820 -41.865 -295.320 ;
        RECT -41.605 -295.820 -41.375 -295.320 ;
        RECT -41.115 -295.820 -40.885 -295.320 ;
        RECT -40.625 -295.820 -40.395 -295.320 ;
        RECT -40.135 -295.820 -39.905 -295.320 ;
        RECT -39.645 -295.820 -39.415 -295.320 ;
        RECT -48.230 -296.505 -47.385 -296.455 ;
        RECT -55.220 -297.720 -54.990 -296.720 ;
        RECT -54.240 -297.720 -54.010 -296.720 ;
        RECT -53.260 -297.720 -53.030 -296.720 ;
        RECT -51.030 -297.645 -50.800 -297.145 ;
        RECT -50.540 -297.645 -50.310 -297.145 ;
        RECT -50.050 -297.645 -49.820 -297.145 ;
        RECT -49.560 -297.645 -49.330 -297.145 ;
        RECT -49.070 -297.645 -48.840 -297.145 ;
        RECT -48.580 -297.645 -48.350 -297.145 ;
        RECT -48.090 -297.645 -47.860 -297.145 ;
        RECT -47.600 -297.645 -47.370 -297.145 ;
        RECT -46.505 -297.720 -46.275 -296.720 ;
        RECT -45.525 -297.720 -45.295 -296.720 ;
        RECT -44.545 -297.720 -44.315 -296.720 ;
        RECT -43.525 -298.060 -43.240 -296.455 ;
        RECT -42.095 -297.720 -41.865 -296.720 ;
        RECT -41.115 -297.720 -40.885 -296.720 ;
        RECT -40.135 -297.720 -39.905 -296.720 ;
        RECT -64.525 -298.345 -43.240 -298.060 ;
        RECT -78.075 -306.740 -74.535 -306.175 ;
        RECT -81.585 -308.715 -81.355 -307.035 ;
        RECT -83.550 -308.950 -81.355 -308.715 ;
        RECT -38.660 -309.865 -37.780 -277.290 ;
        RECT -37.265 -293.215 -37.035 -290.215 ;
        RECT -36.205 -293.215 -35.975 -290.215 ;
        RECT -35.715 -293.215 -35.485 -290.215 ;
        RECT -35.225 -293.215 -34.995 -290.215 ;
        RECT -34.170 -293.215 -33.940 -290.215 ;
        RECT -36.850 -296.275 -36.620 -294.775 ;
        RECT -36.360 -296.275 -36.130 -294.775 ;
        RECT -35.150 -296.275 -34.920 -294.775 ;
        RECT -34.660 -296.275 -34.430 -294.775 ;
        RECT -34.170 -296.275 -33.940 -294.775 ;
        RECT -90.630 -310.665 -89.910 -309.985 ;
        RECT -38.725 -310.720 -37.725 -309.865 ;
        RECT -32.985 -311.155 -32.325 -268.795 ;
        RECT -28.595 -269.225 -28.455 -268.500 ;
        RECT -26.480 -268.490 -25.785 -268.445 ;
        RECT -22.295 -268.490 -21.615 -268.445 ;
        RECT -26.480 -268.630 -21.615 -268.490 ;
        RECT -26.480 -268.715 -25.785 -268.630 ;
        RECT -22.295 -268.675 -21.615 -268.630 ;
        RECT -28.315 -268.860 -27.620 -268.815 ;
        RECT -22.925 -268.850 -22.230 -268.845 ;
        RECT -22.925 -268.860 -20.270 -268.850 ;
        RECT -28.315 -268.990 -20.270 -268.860 ;
        RECT -28.315 -269.000 -22.230 -268.990 ;
        RECT -28.315 -269.085 -27.620 -269.000 ;
        RECT -22.925 -269.115 -22.230 -269.000 ;
        RECT -23.825 -269.225 -23.170 -269.165 ;
        RECT -28.595 -269.365 -23.170 -269.225 ;
        RECT -23.825 -269.395 -23.170 -269.365 ;
        RECT -30.250 -270.555 -30.020 -269.555 ;
        RECT -29.760 -270.555 -29.530 -269.555 ;
        RECT -28.180 -270.555 -27.950 -269.555 ;
        RECT -27.690 -270.555 -27.460 -269.555 ;
        RECT -26.370 -270.555 -26.140 -269.555 ;
        RECT -25.880 -270.555 -25.650 -269.555 ;
        RECT -24.900 -270.555 -24.670 -269.555 ;
        RECT -24.410 -270.555 -24.180 -269.555 ;
        RECT -23.350 -270.555 -23.120 -269.555 ;
        RECT -22.860 -270.555 -22.630 -269.555 ;
        RECT -21.805 -270.555 -21.575 -269.555 ;
        RECT -21.315 -270.555 -21.085 -269.555 ;
        RECT -28.065 -272.270 -27.835 -271.770 ;
        RECT -27.575 -272.270 -27.345 -271.770 ;
        RECT -27.085 -272.270 -26.855 -271.770 ;
        RECT -26.595 -272.270 -26.365 -271.770 ;
        RECT -26.105 -272.270 -25.875 -271.770 ;
        RECT -25.615 -272.270 -25.385 -271.770 ;
        RECT -20.410 -272.185 -20.270 -268.990 ;
        RECT -20.500 -272.865 -20.270 -272.185 ;
        RECT -27.575 -274.170 -27.345 -273.170 ;
        RECT -26.595 -274.170 -26.365 -273.170 ;
        RECT -25.615 -274.170 -25.385 -273.170 ;
        RECT -20.050 -274.345 -19.910 -268.305 ;
        RECT -17.725 -268.360 -17.030 -268.295 ;
        RECT -11.935 -268.305 -7.055 -268.165 ;
        RECT -11.935 -268.345 -11.240 -268.305 ;
        RECT -17.725 -268.500 -15.955 -268.360 ;
        RECT -8.860 -268.375 -8.165 -268.305 ;
        RECT -17.725 -268.565 -17.030 -268.500 ;
        RECT -16.095 -269.225 -15.955 -268.500 ;
        RECT -13.980 -268.490 -13.285 -268.445 ;
        RECT -9.795 -268.490 -9.115 -268.445 ;
        RECT -13.980 -268.630 -9.115 -268.490 ;
        RECT -13.980 -268.715 -13.285 -268.630 ;
        RECT -9.795 -268.675 -9.115 -268.630 ;
        RECT -15.815 -268.860 -15.120 -268.815 ;
        RECT -10.425 -268.850 -9.730 -268.845 ;
        RECT -10.425 -268.860 -7.485 -268.850 ;
        RECT -15.815 -268.990 -7.485 -268.860 ;
        RECT -15.815 -269.000 -9.730 -268.990 ;
        RECT -15.815 -269.085 -15.120 -269.000 ;
        RECT -10.425 -269.115 -9.730 -269.000 ;
        RECT -11.325 -269.225 -10.670 -269.165 ;
        RECT -16.095 -269.365 -10.670 -269.225 ;
        RECT -11.325 -269.395 -10.670 -269.365 ;
        RECT -18.590 -270.390 -18.360 -269.710 ;
        RECT -18.585 -273.240 -18.365 -270.390 ;
        RECT -17.750 -270.555 -17.520 -269.555 ;
        RECT -17.260 -270.555 -17.030 -269.555 ;
        RECT -15.680 -270.555 -15.450 -269.555 ;
        RECT -15.190 -270.555 -14.960 -269.555 ;
        RECT -13.870 -270.555 -13.640 -269.555 ;
        RECT -13.380 -270.555 -13.150 -269.555 ;
        RECT -12.400 -270.555 -12.170 -269.555 ;
        RECT -11.910 -270.555 -11.680 -269.555 ;
        RECT -10.850 -270.555 -10.620 -269.555 ;
        RECT -10.360 -270.555 -10.130 -269.555 ;
        RECT -9.305 -270.555 -9.075 -269.555 ;
        RECT -8.815 -270.555 -8.585 -269.555 ;
        RECT -18.590 -273.920 -18.360 -273.240 ;
        RECT -7.625 -274.010 -7.485 -268.990 ;
        RECT -7.195 -273.595 -7.055 -268.305 ;
        RECT -5.225 -268.360 -4.530 -268.295 ;
        RECT 0.565 -268.305 5.305 -268.165 ;
        RECT 0.565 -268.345 1.260 -268.305 ;
        RECT -5.225 -268.500 -3.455 -268.360 ;
        RECT 3.640 -268.375 4.335 -268.305 ;
        RECT -5.225 -268.565 -4.530 -268.500 ;
        RECT -3.595 -269.225 -3.455 -268.500 ;
        RECT -1.480 -268.490 -0.785 -268.445 ;
        RECT 2.705 -268.490 3.385 -268.445 ;
        RECT -1.480 -268.630 3.385 -268.490 ;
        RECT -1.480 -268.715 -0.785 -268.630 ;
        RECT 2.705 -268.675 3.385 -268.630 ;
        RECT -3.315 -268.860 -2.620 -268.815 ;
        RECT 2.075 -268.850 2.770 -268.845 ;
        RECT 2.075 -268.860 4.935 -268.850 ;
        RECT -3.315 -268.990 4.935 -268.860 ;
        RECT -3.315 -269.000 2.770 -268.990 ;
        RECT -3.315 -269.085 -2.620 -269.000 ;
        RECT 2.075 -269.115 2.770 -269.000 ;
        RECT 1.175 -269.225 1.830 -269.165 ;
        RECT -3.595 -269.365 1.830 -269.225 ;
        RECT 1.175 -269.395 1.830 -269.365 ;
        RECT -5.850 -270.410 -5.620 -269.730 ;
        RECT -5.845 -271.595 -5.625 -270.410 ;
        RECT -5.250 -270.555 -5.020 -269.555 ;
        RECT -4.760 -270.555 -4.530 -269.555 ;
        RECT -3.180 -270.555 -2.950 -269.555 ;
        RECT -2.690 -270.555 -2.460 -269.555 ;
        RECT -1.370 -270.555 -1.140 -269.555 ;
        RECT -0.880 -270.555 -0.650 -269.555 ;
        RECT 0.100 -270.555 0.330 -269.555 ;
        RECT 0.590 -270.555 0.820 -269.555 ;
        RECT 1.650 -270.555 1.880 -269.555 ;
        RECT 2.140 -270.555 2.370 -269.555 ;
        RECT 3.195 -270.555 3.425 -269.555 ;
        RECT 3.685 -270.555 3.915 -269.555 ;
        RECT -5.025 -271.595 -4.345 -271.590 ;
        RECT -5.850 -271.815 -4.345 -271.595 ;
        RECT -5.025 -271.820 -4.345 -271.815 ;
        RECT 4.795 -273.315 4.935 -268.990 ;
        RECT 5.165 -273.030 5.305 -268.305 ;
        RECT 7.275 -268.360 7.970 -268.295 ;
        RECT 13.065 -268.305 17.680 -268.165 ;
        RECT 13.065 -268.345 13.760 -268.305 ;
        RECT 7.275 -268.500 9.045 -268.360 ;
        RECT 16.140 -268.375 16.835 -268.305 ;
        RECT 7.275 -268.565 7.970 -268.500 ;
        RECT 8.905 -269.225 9.045 -268.500 ;
        RECT 11.020 -268.490 11.715 -268.445 ;
        RECT 15.205 -268.490 15.885 -268.445 ;
        RECT 11.020 -268.630 15.885 -268.490 ;
        RECT 11.020 -268.715 11.715 -268.630 ;
        RECT 15.205 -268.675 15.885 -268.630 ;
        RECT 9.185 -268.860 9.880 -268.815 ;
        RECT 14.575 -268.850 15.270 -268.845 ;
        RECT 14.575 -268.860 17.265 -268.850 ;
        RECT 9.185 -268.990 17.265 -268.860 ;
        RECT 9.185 -269.000 15.270 -268.990 ;
        RECT 9.185 -269.085 9.880 -269.000 ;
        RECT 14.575 -269.115 15.270 -269.000 ;
        RECT 13.675 -269.225 14.330 -269.165 ;
        RECT 8.905 -269.365 14.330 -269.225 ;
        RECT 13.675 -269.395 14.330 -269.365 ;
        RECT 6.550 -270.410 6.780 -269.730 ;
        RECT 6.555 -271.660 6.775 -270.410 ;
        RECT 7.250 -270.555 7.480 -269.555 ;
        RECT 7.740 -270.555 7.970 -269.555 ;
        RECT 9.320 -270.555 9.550 -269.555 ;
        RECT 9.810 -270.555 10.040 -269.555 ;
        RECT 11.130 -270.555 11.360 -269.555 ;
        RECT 11.620 -270.555 11.850 -269.555 ;
        RECT 12.600 -270.555 12.830 -269.555 ;
        RECT 13.090 -270.555 13.320 -269.555 ;
        RECT 14.150 -270.555 14.380 -269.555 ;
        RECT 14.640 -270.555 14.870 -269.555 ;
        RECT 15.695 -270.555 15.925 -269.555 ;
        RECT 16.185 -270.555 16.415 -269.555 ;
        RECT 7.460 -271.660 8.140 -271.655 ;
        RECT 6.555 -271.880 8.140 -271.660 ;
        RECT 7.460 -271.885 8.140 -271.880 ;
        RECT 17.125 -272.715 17.265 -268.990 ;
        RECT 17.540 -272.345 17.680 -268.305 ;
        RECT 19.775 -268.360 20.470 -268.295 ;
        RECT 25.565 -268.305 34.205 -268.165 ;
        RECT 25.565 -268.345 26.260 -268.305 ;
        RECT 19.775 -268.500 21.545 -268.360 ;
        RECT 28.640 -268.375 29.335 -268.305 ;
        RECT 19.775 -268.565 20.470 -268.500 ;
        RECT 21.405 -269.225 21.545 -268.500 ;
        RECT 23.520 -268.490 24.215 -268.445 ;
        RECT 27.705 -268.490 28.385 -268.445 ;
        RECT 23.520 -268.630 28.385 -268.490 ;
        RECT 23.520 -268.715 24.215 -268.630 ;
        RECT 27.705 -268.675 28.385 -268.630 ;
        RECT 26.175 -269.225 26.830 -269.165 ;
        RECT 21.405 -269.365 26.830 -269.225 ;
        RECT 26.175 -269.395 26.830 -269.365 ;
        RECT 18.635 -270.410 18.865 -269.730 ;
        RECT 18.640 -271.970 18.860 -270.410 ;
        RECT 19.750 -270.555 19.980 -269.555 ;
        RECT 20.240 -270.555 20.470 -269.555 ;
        RECT 21.820 -270.555 22.050 -269.555 ;
        RECT 22.310 -270.555 22.540 -269.555 ;
        RECT 23.630 -270.555 23.860 -269.555 ;
        RECT 24.120 -270.555 24.350 -269.555 ;
        RECT 25.100 -270.555 25.330 -269.555 ;
        RECT 25.590 -270.555 25.820 -269.555 ;
        RECT 26.650 -270.555 26.880 -269.555 ;
        RECT 27.140 -270.555 27.370 -269.555 ;
        RECT 28.195 -270.555 28.425 -269.555 ;
        RECT 28.685 -270.555 28.915 -269.555 ;
        RECT 33.160 -270.410 33.390 -269.730 ;
        RECT 33.165 -271.890 33.385 -270.410 ;
        RECT 34.065 -271.680 34.205 -268.305 ;
        RECT 34.775 -268.360 35.470 -268.295 ;
        RECT 40.565 -268.305 54.990 -268.165 ;
        RECT 40.565 -268.345 41.260 -268.305 ;
        RECT 34.775 -268.500 36.545 -268.360 ;
        RECT 43.640 -268.375 44.335 -268.305 ;
        RECT 34.775 -268.565 35.470 -268.500 ;
        RECT 36.405 -269.225 36.545 -268.500 ;
        RECT 38.520 -268.490 39.215 -268.445 ;
        RECT 42.705 -268.490 43.385 -268.445 ;
        RECT 38.520 -268.630 43.385 -268.490 ;
        RECT 38.520 -268.715 39.215 -268.630 ;
        RECT 42.705 -268.675 43.385 -268.630 ;
        RECT 41.175 -269.225 41.830 -269.165 ;
        RECT 36.405 -269.365 41.830 -269.225 ;
        RECT 41.175 -269.395 41.830 -269.365 ;
        RECT 34.750 -270.555 34.980 -269.555 ;
        RECT 35.240 -270.555 35.470 -269.555 ;
        RECT 36.820 -270.555 37.050 -269.555 ;
        RECT 37.310 -270.555 37.540 -269.555 ;
        RECT 38.630 -270.555 38.860 -269.555 ;
        RECT 39.120 -270.555 39.350 -269.555 ;
        RECT 40.100 -270.555 40.330 -269.555 ;
        RECT 40.590 -270.555 40.820 -269.555 ;
        RECT 41.650 -270.555 41.880 -269.555 ;
        RECT 42.140 -270.555 42.370 -269.555 ;
        RECT 43.195 -270.555 43.425 -269.555 ;
        RECT 43.685 -270.555 43.915 -269.555 ;
        RECT 48.205 -271.680 54.165 -271.095 ;
        RECT 34.065 -271.820 54.210 -271.680 ;
        RECT 18.375 -272.200 19.055 -271.970 ;
        RECT 32.900 -272.120 33.580 -271.890 ;
        RECT 17.540 -272.535 53.445 -272.345 ;
        RECT 17.125 -272.855 53.070 -272.715 ;
        RECT 5.165 -273.170 52.685 -273.030 ;
        RECT 4.795 -273.455 52.260 -273.315 ;
        RECT -7.195 -273.850 51.890 -273.595 ;
        RECT -7.625 -274.190 51.465 -274.010 ;
        RECT -20.050 -274.600 51.110 -274.345 ;
        RECT -18.575 -275.195 -17.895 -275.185 ;
        RECT 16.670 -275.195 17.350 -275.175 ;
        RECT -18.575 -275.405 17.350 -275.195 ;
        RECT -18.575 -275.415 -17.895 -275.405 ;
        RECT -30.975 -275.605 -30.295 -275.595 ;
        RECT 16.150 -275.605 16.925 -275.595 ;
        RECT -30.975 -275.815 16.925 -275.605 ;
        RECT -30.975 -275.825 -30.295 -275.815 ;
        RECT 16.150 -275.825 16.925 -275.815 ;
        RECT -29.350 -278.685 -29.120 -277.685 ;
        RECT -28.370 -278.685 -28.140 -277.685 ;
        RECT -27.390 -278.685 -27.160 -277.685 ;
        RECT -25.160 -278.260 -24.930 -277.760 ;
        RECT -24.670 -278.260 -24.440 -277.760 ;
        RECT -24.180 -278.260 -23.950 -277.760 ;
        RECT -23.690 -278.260 -23.460 -277.760 ;
        RECT -23.200 -278.260 -22.970 -277.760 ;
        RECT -22.710 -278.260 -22.480 -277.760 ;
        RECT -22.220 -278.260 -21.990 -277.760 ;
        RECT -21.730 -278.260 -21.500 -277.760 ;
        RECT -20.635 -278.685 -20.405 -277.685 ;
        RECT -19.655 -278.685 -19.425 -277.685 ;
        RECT -18.675 -278.685 -18.445 -277.685 ;
        RECT -22.360 -278.950 -21.515 -278.900 ;
        RECT -17.655 -278.950 -17.370 -277.775 ;
        RECT -15.850 -278.685 -15.620 -277.685 ;
        RECT -14.870 -278.685 -14.640 -277.685 ;
        RECT -13.890 -278.685 -13.660 -277.685 ;
        RECT -11.660 -278.260 -11.430 -277.760 ;
        RECT -11.170 -278.260 -10.940 -277.760 ;
        RECT -10.680 -278.260 -10.450 -277.760 ;
        RECT -10.190 -278.260 -9.960 -277.760 ;
        RECT -9.700 -278.260 -9.470 -277.760 ;
        RECT -9.210 -278.260 -8.980 -277.760 ;
        RECT -8.720 -278.260 -8.490 -277.760 ;
        RECT -8.230 -278.260 -8.000 -277.760 ;
        RECT -7.135 -278.685 -6.905 -277.685 ;
        RECT -6.155 -278.685 -5.925 -277.685 ;
        RECT -5.175 -278.685 -4.945 -277.685 ;
        RECT -22.360 -279.235 -17.370 -278.950 ;
        RECT -8.860 -278.950 -8.015 -278.900 ;
        RECT -4.155 -278.950 -3.870 -277.775 ;
        RECT -2.725 -278.685 -2.495 -277.685 ;
        RECT -1.745 -278.685 -1.515 -277.685 ;
        RECT -0.765 -278.685 -0.535 -277.685 ;
        RECT 1.925 -278.770 2.155 -277.770 ;
        RECT 5.615 -278.770 5.845 -277.770 ;
        RECT 6.595 -278.770 6.825 -277.770 ;
        RECT 7.575 -278.770 7.805 -277.770 ;
        RECT 8.705 -278.575 8.935 -278.565 ;
        RECT -22.360 -279.270 -21.515 -279.235 ;
        RECT -29.350 -280.085 -29.120 -279.585 ;
        RECT -28.860 -280.085 -28.630 -279.585 ;
        RECT -28.370 -280.085 -28.140 -279.585 ;
        RECT -27.880 -280.085 -27.650 -279.585 ;
        RECT -27.390 -280.085 -27.160 -279.585 ;
        RECT -26.900 -280.085 -26.670 -279.585 ;
        RECT -25.160 -280.060 -24.930 -279.835 ;
        RECT -28.225 -280.670 -27.565 -280.370 ;
        RECT -29.920 -281.150 -29.620 -281.020 ;
        RECT -31.695 -281.465 -29.620 -281.150 ;
        RECT -31.610 -281.470 -29.620 -281.465 ;
        RECT -29.920 -281.705 -29.620 -281.470 ;
        RECT -28.105 -281.760 -27.630 -280.670 ;
        RECT -25.170 -280.830 -24.930 -280.060 ;
        RECT -24.670 -280.335 -24.440 -279.835 ;
        RECT -24.180 -280.240 -23.950 -279.835 ;
        RECT -24.210 -280.830 -23.905 -280.240 ;
        RECT -23.690 -280.335 -23.460 -279.835 ;
        RECT -23.200 -280.230 -22.970 -279.835 ;
        RECT -23.230 -280.830 -22.925 -280.230 ;
        RECT -22.710 -280.335 -22.480 -279.835 ;
        RECT -22.220 -280.240 -21.990 -279.835 ;
        RECT -22.275 -280.830 -21.970 -280.240 ;
        RECT -21.730 -280.335 -21.500 -279.835 ;
        RECT -20.635 -280.085 -20.405 -279.585 ;
        RECT -20.145 -280.085 -19.915 -279.585 ;
        RECT -19.655 -280.085 -19.425 -279.585 ;
        RECT -19.165 -280.085 -18.935 -279.585 ;
        RECT -18.675 -280.085 -18.445 -279.585 ;
        RECT -18.185 -280.085 -17.955 -279.585 ;
        RECT -25.170 -281.070 -17.515 -280.830 ;
        RECT -28.180 -282.060 -27.495 -281.760 ;
        RECT -29.350 -283.375 -29.120 -282.875 ;
        RECT -28.860 -283.375 -28.630 -282.875 ;
        RECT -28.370 -283.375 -28.140 -282.875 ;
        RECT -27.880 -283.375 -27.650 -282.875 ;
        RECT -27.390 -283.375 -27.160 -282.875 ;
        RECT -26.900 -283.375 -26.670 -282.875 ;
        RECT -25.165 -283.375 -24.935 -282.875 ;
        RECT -24.675 -283.375 -24.445 -282.875 ;
        RECT -24.185 -283.375 -23.955 -282.875 ;
        RECT -23.695 -283.375 -23.465 -282.875 ;
        RECT -23.205 -283.375 -22.975 -282.875 ;
        RECT -22.715 -283.375 -22.485 -282.875 ;
        RECT -21.620 -283.125 -21.390 -282.625 ;
        RECT -21.130 -283.125 -20.900 -282.625 ;
        RECT -20.640 -283.125 -20.410 -282.625 ;
        RECT -20.150 -283.125 -19.920 -282.625 ;
        RECT -19.660 -283.125 -19.430 -282.625 ;
        RECT -19.170 -283.125 -18.940 -282.625 ;
        RECT -18.680 -283.125 -18.450 -282.625 ;
        RECT -18.190 -283.125 -17.960 -282.625 ;
        RECT -17.720 -283.495 -17.515 -281.070 ;
        RECT -17.125 -281.315 -16.825 -279.075 ;
        RECT -16.550 -279.635 -16.250 -279.200 ;
        RECT -8.860 -279.235 -3.870 -278.950 ;
        RECT -8.860 -279.270 -8.015 -279.235 ;
        RECT -16.550 -279.860 -16.245 -279.635 ;
        RECT -17.370 -281.615 -16.685 -281.315 ;
        RECT -21.605 -283.725 -20.760 -283.690 ;
        RECT -25.750 -284.010 -20.760 -283.725 ;
        RECT -18.195 -283.795 -17.510 -283.495 ;
        RECT -16.545 -283.600 -16.245 -279.860 ;
        RECT -15.850 -280.085 -15.620 -279.585 ;
        RECT -15.360 -280.085 -15.130 -279.585 ;
        RECT -14.870 -280.085 -14.640 -279.585 ;
        RECT -14.380 -280.085 -14.150 -279.585 ;
        RECT -13.890 -280.085 -13.660 -279.585 ;
        RECT -13.400 -280.085 -13.170 -279.585 ;
        RECT -11.660 -280.335 -11.415 -279.835 ;
        RECT -11.170 -280.335 -10.940 -279.835 ;
        RECT -10.680 -280.335 -10.450 -279.835 ;
        RECT -10.190 -280.335 -9.960 -279.835 ;
        RECT -9.700 -280.335 -9.470 -279.835 ;
        RECT -9.210 -280.335 -8.980 -279.835 ;
        RECT -8.720 -280.335 -8.490 -279.835 ;
        RECT -8.230 -280.335 -8.000 -279.835 ;
        RECT -7.135 -280.085 -6.905 -279.585 ;
        RECT -6.645 -280.085 -6.415 -279.585 ;
        RECT -6.155 -280.085 -5.925 -279.585 ;
        RECT -5.665 -280.085 -5.435 -279.585 ;
        RECT -5.175 -280.085 -4.945 -279.585 ;
        RECT -4.685 -280.085 -4.455 -279.585 ;
        RECT -15.230 -280.690 -14.545 -280.390 ;
        RECT -15.140 -281.730 -14.665 -280.690 ;
        RECT -11.645 -280.820 -11.415 -280.335 ;
        RECT -10.670 -280.820 -10.460 -280.335 ;
        RECT -9.695 -280.820 -9.485 -280.335 ;
        RECT -8.715 -280.820 -8.505 -280.335 ;
        RECT -11.645 -281.050 -7.845 -280.820 ;
        RECT -12.640 -281.610 -11.980 -281.310 ;
        RECT -15.195 -282.030 -14.510 -281.730 ;
        RECT -15.850 -283.375 -15.620 -282.875 ;
        RECT -15.360 -283.375 -15.130 -282.875 ;
        RECT -14.870 -283.375 -14.640 -282.875 ;
        RECT -14.380 -283.375 -14.150 -282.875 ;
        RECT -13.890 -283.375 -13.660 -282.875 ;
        RECT -13.400 -283.375 -13.170 -282.875 ;
        RECT -12.495 -283.430 -12.195 -281.610 ;
        RECT -8.075 -281.880 -7.845 -281.050 ;
        RECT -4.155 -281.420 -3.870 -279.235 ;
        RECT -3.465 -279.740 -3.165 -279.080 ;
        RECT 8.665 -279.245 8.935 -278.575 ;
        RECT 10.590 -278.615 10.820 -277.835 ;
        RECT 11.570 -278.605 11.800 -277.835 ;
        RECT 11.080 -278.615 12.290 -278.605 ;
        RECT 12.550 -278.615 12.780 -277.835 ;
        RECT 10.465 -278.845 12.780 -278.615 ;
        RECT -3.455 -280.880 -3.165 -279.740 ;
        RECT -2.725 -280.085 -2.495 -279.585 ;
        RECT -2.235 -280.085 -2.005 -279.585 ;
        RECT -1.745 -280.085 -1.515 -279.585 ;
        RECT -1.255 -280.085 -1.025 -279.585 ;
        RECT -0.765 -280.085 -0.535 -279.585 ;
        RECT -0.275 -280.085 -0.045 -279.585 ;
        RECT 1.200 -280.065 1.905 -279.800 ;
        RECT -1.445 -280.685 -0.760 -280.385 ;
        RECT -3.455 -281.170 -2.260 -280.880 ;
        RECT -2.550 -281.315 -2.260 -281.170 ;
        RECT -4.155 -281.705 -2.825 -281.420 ;
        RECT -2.570 -281.615 -1.910 -281.315 ;
        RECT -8.075 -281.885 -4.020 -281.880 ;
        RECT -8.075 -282.110 -3.980 -281.885 ;
        RECT -11.665 -283.375 -11.435 -282.875 ;
        RECT -11.175 -283.375 -10.945 -282.875 ;
        RECT -10.685 -283.375 -10.455 -282.875 ;
        RECT -10.195 -283.375 -9.965 -282.875 ;
        RECT -9.705 -283.375 -9.475 -282.875 ;
        RECT -9.215 -283.375 -8.985 -282.875 ;
        RECT -8.120 -283.125 -7.890 -282.625 ;
        RECT -7.630 -283.125 -7.400 -282.625 ;
        RECT -7.140 -283.125 -6.910 -282.625 ;
        RECT -6.650 -283.125 -6.420 -282.625 ;
        RECT -6.160 -283.125 -5.930 -282.625 ;
        RECT -5.670 -283.125 -5.440 -282.625 ;
        RECT -5.180 -283.125 -4.950 -282.625 ;
        RECT -4.690 -283.125 -4.460 -282.625 ;
        RECT -4.210 -283.485 -3.980 -282.110 ;
        RECT -3.110 -282.310 -2.825 -281.705 ;
        RECT -1.270 -281.730 -0.795 -280.685 ;
        RECT -1.355 -282.030 -0.695 -281.730 ;
        RECT 1.200 -282.310 1.485 -280.065 ;
        RECT 1.925 -282.310 2.155 -281.310 ;
        RECT 2.415 -282.310 2.645 -281.310 ;
        RECT 3.990 -282.310 4.220 -280.810 ;
        RECT 4.480 -282.310 4.710 -280.810 ;
        RECT 4.970 -282.310 5.200 -280.810 ;
        RECT 5.535 -282.310 5.765 -280.810 ;
        RECT 6.025 -282.310 6.255 -280.810 ;
        RECT 6.515 -282.310 6.745 -280.810 ;
        RECT 7.085 -282.305 7.315 -280.805 ;
        RECT 7.575 -282.305 7.805 -280.805 ;
        RECT 8.065 -282.305 8.295 -280.805 ;
        RECT -3.110 -282.595 1.485 -282.310 ;
        RECT -17.720 -283.800 -17.515 -283.795 ;
        RECT -16.545 -283.900 -15.830 -283.600 ;
        RECT -8.105 -283.725 -7.260 -283.690 ;
        RECT -16.545 -283.930 -16.245 -283.900 ;
        RECT -28.860 -285.275 -28.630 -284.275 ;
        RECT -27.880 -285.275 -27.650 -284.275 ;
        RECT -26.900 -285.275 -26.670 -284.275 ;
        RECT -25.750 -285.185 -25.465 -284.010 ;
        RECT -21.605 -284.060 -20.760 -284.010 ;
        RECT -12.250 -284.010 -7.260 -283.725 ;
        RECT -4.750 -283.785 -3.980 -283.485 ;
        RECT 8.665 -283.270 8.895 -279.245 ;
        RECT 9.110 -279.665 9.790 -279.435 ;
        RECT 11.080 -279.490 11.310 -278.845 ;
        RECT 11.570 -279.490 11.800 -278.990 ;
        RECT 12.060 -279.490 12.290 -278.845 ;
        RECT 12.550 -279.490 12.780 -278.990 ;
        RECT 9.430 -282.710 9.660 -279.665 ;
        RECT 14.125 -282.205 14.355 -280.525 ;
        RECT 14.615 -282.025 14.845 -277.840 ;
        RECT 15.595 -279.340 15.825 -277.840 ;
        RECT 18.615 -278.625 18.845 -277.845 ;
        RECT 19.595 -278.615 19.825 -277.845 ;
        RECT 19.105 -278.625 20.315 -278.615 ;
        RECT 20.575 -278.625 20.805 -277.845 ;
        RECT 18.490 -278.855 20.805 -278.625 ;
        RECT 19.105 -279.500 19.335 -278.855 ;
        RECT 19.595 -279.500 19.825 -279.000 ;
        RECT 20.085 -279.500 20.315 -278.855 ;
        RECT 20.575 -279.500 20.805 -279.000 ;
        RECT 15.105 -282.205 15.335 -280.525 ;
        RECT 15.595 -282.025 15.825 -280.525 ;
        RECT 16.085 -282.020 16.315 -280.525 ;
        RECT 16.085 -282.205 16.320 -282.020 ;
        RECT 14.125 -282.440 16.320 -282.205 ;
        RECT 22.150 -282.215 22.380 -280.535 ;
        RECT 22.640 -282.035 22.870 -277.850 ;
        RECT 23.620 -279.350 23.850 -277.850 ;
        RECT 26.735 -278.725 26.965 -277.725 ;
        RECT 30.425 -278.725 30.655 -277.725 ;
        RECT 31.405 -278.725 31.635 -277.725 ;
        RECT 32.385 -278.725 32.615 -277.725 ;
        RECT 34.800 -278.780 35.030 -277.780 ;
        RECT 35.290 -278.935 35.520 -277.780 ;
        RECT 35.780 -278.780 36.010 -277.780 ;
        RECT 36.380 -278.780 36.610 -277.780 ;
        RECT 36.870 -278.780 37.100 -277.780 ;
        RECT 37.360 -278.780 37.590 -277.780 ;
        RECT 39.170 -278.780 39.400 -277.780 ;
        RECT 40.150 -278.780 40.380 -277.780 ;
        RECT 41.700 -278.780 41.930 -277.780 ;
        RECT 43.245 -278.780 43.475 -277.780 ;
        RECT 32.760 -279.165 35.520 -278.935 ;
        RECT 32.780 -279.210 33.460 -279.165 ;
        RECT 40.615 -279.420 41.310 -279.330 ;
        RECT 43.690 -279.385 44.385 -279.360 ;
        RECT 48.345 -279.385 49.435 -279.090 ;
        RECT 43.690 -279.420 49.435 -279.385 ;
        RECT 40.615 -279.525 49.435 -279.420 ;
        RECT 34.825 -279.615 35.520 -279.550 ;
        RECT 40.615 -279.560 44.890 -279.525 ;
        RECT 48.345 -279.535 49.435 -279.525 ;
        RECT 40.615 -279.600 41.310 -279.560 ;
        RECT 34.825 -279.755 36.595 -279.615 ;
        RECT 43.690 -279.630 44.385 -279.560 ;
        RECT 34.825 -279.820 35.520 -279.755 ;
        RECT 36.455 -280.480 36.595 -279.755 ;
        RECT 38.570 -279.745 39.265 -279.700 ;
        RECT 42.755 -279.745 43.435 -279.700 ;
        RECT 38.570 -279.885 43.435 -279.745 ;
        RECT 38.570 -279.970 39.265 -279.885 ;
        RECT 42.755 -279.930 43.435 -279.885 ;
        RECT 41.225 -280.480 41.880 -280.420 ;
        RECT 23.130 -282.215 23.360 -280.535 ;
        RECT 23.620 -282.035 23.850 -280.535 ;
        RECT 24.110 -282.030 24.340 -280.535 ;
        RECT 36.455 -280.620 41.880 -280.480 ;
        RECT 41.225 -280.650 41.880 -280.620 ;
        RECT 24.110 -282.215 24.345 -282.030 ;
        RECT 22.150 -282.450 24.345 -282.215 ;
        RECT 26.735 -282.265 26.965 -281.265 ;
        RECT 27.225 -282.265 27.455 -281.265 ;
        RECT 28.800 -282.265 29.030 -280.765 ;
        RECT 29.290 -282.265 29.520 -280.765 ;
        RECT 29.780 -282.265 30.010 -280.765 ;
        RECT 30.345 -282.265 30.575 -280.765 ;
        RECT 30.835 -282.265 31.065 -280.765 ;
        RECT 31.325 -282.265 31.555 -280.765 ;
        RECT 31.895 -282.260 32.125 -280.760 ;
        RECT 32.385 -282.260 32.615 -280.760 ;
        RECT 32.875 -282.260 33.105 -280.760 ;
        RECT 34.800 -281.810 35.030 -280.810 ;
        RECT 35.290 -281.810 35.520 -280.810 ;
        RECT 36.870 -281.810 37.100 -280.810 ;
        RECT 37.360 -281.810 37.590 -280.810 ;
        RECT 38.680 -281.810 38.910 -280.810 ;
        RECT 39.170 -281.810 39.400 -280.810 ;
        RECT 40.150 -281.810 40.380 -280.810 ;
        RECT 40.640 -281.810 40.870 -280.810 ;
        RECT 41.700 -281.810 41.930 -280.810 ;
        RECT 42.190 -281.810 42.420 -280.810 ;
        RECT 43.245 -281.810 43.475 -280.810 ;
        RECT 43.735 -281.810 43.965 -280.810 ;
        RECT 9.430 -282.940 18.175 -282.710 ;
        RECT 8.665 -283.500 26.015 -283.270 ;
        RECT -24.675 -285.275 -24.445 -284.275 ;
        RECT -23.695 -285.275 -23.465 -284.275 ;
        RECT -22.715 -285.275 -22.485 -284.275 ;
        RECT -21.620 -285.200 -21.390 -284.700 ;
        RECT -21.130 -285.200 -20.900 -284.700 ;
        RECT -20.640 -285.200 -20.410 -284.700 ;
        RECT -20.150 -285.200 -19.920 -284.700 ;
        RECT -19.660 -285.200 -19.430 -284.700 ;
        RECT -19.170 -285.200 -18.940 -284.700 ;
        RECT -18.680 -285.200 -18.450 -284.700 ;
        RECT -18.190 -285.200 -17.960 -284.700 ;
        RECT -15.360 -285.275 -15.130 -284.275 ;
        RECT -14.380 -285.275 -14.150 -284.275 ;
        RECT -13.400 -285.275 -13.170 -284.275 ;
        RECT -12.250 -285.185 -11.965 -284.010 ;
        RECT -8.105 -284.060 -7.260 -284.010 ;
        RECT -11.175 -285.275 -10.945 -284.275 ;
        RECT -10.195 -285.275 -9.965 -284.275 ;
        RECT -9.215 -285.275 -8.985 -284.275 ;
        RECT -8.120 -285.200 -7.890 -284.700 ;
        RECT -7.630 -285.200 -7.400 -284.700 ;
        RECT -7.140 -285.200 -6.910 -284.700 ;
        RECT -6.650 -285.200 -6.420 -284.700 ;
        RECT -6.160 -285.200 -5.930 -284.700 ;
        RECT -5.670 -285.200 -5.440 -284.700 ;
        RECT -5.180 -285.200 -4.950 -284.700 ;
        RECT -4.690 -285.200 -4.460 -284.700 ;
        RECT -28.860 -292.465 -28.630 -291.465 ;
        RECT -27.880 -292.465 -27.650 -291.465 ;
        RECT -26.900 -292.465 -26.670 -291.465 ;
        RECT -25.750 -292.730 -25.465 -291.555 ;
        RECT -24.675 -292.465 -24.445 -291.465 ;
        RECT -23.695 -292.465 -23.465 -291.465 ;
        RECT -22.715 -292.465 -22.485 -291.465 ;
        RECT -21.620 -292.040 -21.390 -291.540 ;
        RECT -21.130 -292.040 -20.900 -291.540 ;
        RECT -20.640 -292.040 -20.410 -291.540 ;
        RECT -20.150 -292.040 -19.920 -291.540 ;
        RECT -19.660 -292.040 -19.430 -291.540 ;
        RECT -19.170 -292.040 -18.940 -291.540 ;
        RECT -18.680 -292.040 -18.450 -291.540 ;
        RECT -18.190 -292.040 -17.960 -291.540 ;
        RECT -15.360 -292.465 -15.130 -291.465 ;
        RECT -14.380 -292.465 -14.150 -291.465 ;
        RECT -13.400 -292.465 -13.170 -291.465 ;
        RECT -21.605 -292.730 -20.760 -292.680 ;
        RECT -25.750 -293.015 -20.760 -292.730 ;
        RECT -12.250 -292.730 -11.965 -291.555 ;
        RECT -11.175 -292.465 -10.945 -291.465 ;
        RECT -10.195 -292.465 -9.965 -291.465 ;
        RECT -9.215 -292.465 -8.985 -291.465 ;
        RECT -8.120 -292.040 -7.890 -291.540 ;
        RECT -7.630 -292.040 -7.400 -291.540 ;
        RECT -7.140 -292.040 -6.910 -291.540 ;
        RECT -6.650 -292.040 -6.420 -291.540 ;
        RECT -6.160 -292.040 -5.930 -291.540 ;
        RECT -5.670 -292.040 -5.440 -291.540 ;
        RECT -5.180 -292.040 -4.950 -291.540 ;
        RECT -4.690 -292.040 -4.460 -291.540 ;
        RECT -8.105 -292.730 -7.260 -292.680 ;
        RECT -16.545 -292.840 -16.245 -292.810 ;
        RECT -17.720 -292.945 -17.515 -292.940 ;
        RECT -21.605 -293.050 -20.760 -293.015 ;
        RECT -29.350 -293.865 -29.120 -293.365 ;
        RECT -28.860 -293.865 -28.630 -293.365 ;
        RECT -28.370 -293.865 -28.140 -293.365 ;
        RECT -27.880 -293.865 -27.650 -293.365 ;
        RECT -27.390 -293.865 -27.160 -293.365 ;
        RECT -26.900 -293.865 -26.670 -293.365 ;
        RECT -31.650 -295.270 -30.775 -294.175 ;
        RECT -28.180 -294.980 -27.495 -294.680 ;
        RECT -29.920 -295.270 -29.620 -295.035 ;
        RECT -31.650 -295.590 -29.620 -295.270 ;
        RECT -31.650 -295.745 -30.775 -295.590 ;
        RECT -29.920 -295.720 -29.620 -295.590 ;
        RECT -28.105 -295.920 -27.630 -294.980 ;
        RECT -26.055 -295.570 -25.755 -293.235 ;
        RECT -18.195 -293.245 -17.510 -292.945 ;
        RECT -16.545 -293.140 -15.830 -292.840 ;
        RECT -12.250 -293.015 -7.260 -292.730 ;
        RECT -8.105 -293.050 -7.260 -293.015 ;
        RECT -25.165 -293.865 -24.935 -293.365 ;
        RECT -24.675 -293.865 -24.445 -293.365 ;
        RECT -24.185 -293.865 -23.955 -293.365 ;
        RECT -23.695 -293.865 -23.465 -293.365 ;
        RECT -23.205 -293.865 -22.975 -293.365 ;
        RECT -22.715 -293.865 -22.485 -293.365 ;
        RECT -21.620 -294.115 -21.390 -293.615 ;
        RECT -21.130 -294.115 -20.900 -293.615 ;
        RECT -20.640 -294.115 -20.410 -293.615 ;
        RECT -20.150 -294.115 -19.920 -293.615 ;
        RECT -19.660 -294.115 -19.430 -293.615 ;
        RECT -19.170 -294.115 -18.940 -293.615 ;
        RECT -18.680 -294.115 -18.450 -293.615 ;
        RECT -18.190 -294.115 -17.960 -293.615 ;
        RECT -26.235 -295.870 -25.575 -295.570 ;
        RECT -17.720 -295.670 -17.515 -293.245 ;
        RECT -30.540 -296.070 -27.630 -295.920 ;
        RECT -25.170 -295.910 -17.515 -295.670 ;
        RECT -30.540 -296.370 -27.565 -296.070 ;
        RECT -30.540 -296.395 -27.630 -296.370 ;
        RECT -30.540 -296.790 -30.065 -296.395 ;
        RECT -31.615 -297.265 -30.065 -296.790 ;
        RECT -29.350 -297.155 -29.120 -296.655 ;
        RECT -28.860 -297.155 -28.630 -296.655 ;
        RECT -28.370 -297.155 -28.140 -296.655 ;
        RECT -27.880 -297.155 -27.650 -296.655 ;
        RECT -27.390 -297.155 -27.160 -296.655 ;
        RECT -26.900 -297.155 -26.670 -296.655 ;
        RECT -25.170 -296.680 -24.930 -295.910 ;
        RECT -25.160 -296.905 -24.930 -296.680 ;
        RECT -24.670 -296.905 -24.440 -296.405 ;
        RECT -24.210 -296.500 -23.905 -295.910 ;
        RECT -24.180 -296.905 -23.950 -296.500 ;
        RECT -23.690 -296.905 -23.460 -296.405 ;
        RECT -23.230 -296.510 -22.925 -295.910 ;
        RECT -23.200 -296.905 -22.970 -296.510 ;
        RECT -22.710 -296.905 -22.480 -296.405 ;
        RECT -22.275 -296.500 -21.970 -295.910 ;
        RECT -22.220 -296.905 -21.990 -296.500 ;
        RECT -21.730 -296.905 -21.500 -296.405 ;
        RECT -20.635 -297.155 -20.405 -296.655 ;
        RECT -20.145 -297.155 -19.915 -296.655 ;
        RECT -19.655 -297.155 -19.425 -296.655 ;
        RECT -19.165 -297.155 -18.935 -296.655 ;
        RECT -18.675 -297.155 -18.445 -296.655 ;
        RECT -18.185 -297.155 -17.955 -296.655 ;
        RECT -16.545 -296.880 -16.245 -293.140 ;
        RECT -4.750 -293.255 -3.980 -292.955 ;
        RECT -15.850 -293.865 -15.620 -293.365 ;
        RECT -15.360 -293.865 -15.130 -293.365 ;
        RECT -14.870 -293.865 -14.640 -293.365 ;
        RECT -14.380 -293.865 -14.150 -293.365 ;
        RECT -13.890 -293.865 -13.660 -293.365 ;
        RECT -13.400 -293.865 -13.170 -293.365 ;
        RECT -11.665 -293.865 -11.435 -293.365 ;
        RECT -11.175 -293.865 -10.945 -293.365 ;
        RECT -10.685 -293.865 -10.455 -293.365 ;
        RECT -10.195 -293.865 -9.965 -293.365 ;
        RECT -9.705 -293.865 -9.475 -293.365 ;
        RECT -9.215 -293.865 -8.985 -293.365 ;
        RECT -8.120 -294.115 -7.890 -293.615 ;
        RECT -7.630 -294.115 -7.400 -293.615 ;
        RECT -7.140 -294.115 -6.910 -293.615 ;
        RECT -6.650 -294.115 -6.420 -293.615 ;
        RECT -6.160 -294.115 -5.930 -293.615 ;
        RECT -5.670 -294.115 -5.440 -293.615 ;
        RECT -5.180 -294.115 -4.950 -293.615 ;
        RECT -4.690 -294.115 -4.460 -293.615 ;
        RECT -4.210 -294.630 -3.980 -293.255 ;
        RECT 8.665 -293.470 26.015 -293.240 ;
        RECT -15.195 -295.010 -14.510 -294.710 ;
        RECT -8.075 -294.855 -3.980 -294.630 ;
        RECT -3.110 -294.430 1.485 -294.145 ;
        RECT -8.075 -294.860 -4.020 -294.855 ;
        RECT -15.140 -296.050 -14.665 -295.010 ;
        RECT -8.075 -295.690 -7.845 -294.860 ;
        RECT -3.110 -295.035 -2.825 -294.430 ;
        RECT -2.005 -295.010 -1.345 -294.710 ;
        RECT -11.645 -295.920 -7.845 -295.690 ;
        RECT -4.155 -295.320 -2.825 -295.035 ;
        RECT -15.230 -296.350 -14.545 -296.050 ;
        RECT -11.645 -296.405 -11.415 -295.920 ;
        RECT -10.670 -296.405 -10.460 -295.920 ;
        RECT -9.695 -296.405 -9.485 -295.920 ;
        RECT -8.715 -296.405 -8.505 -295.920 ;
        RECT -16.550 -297.105 -16.245 -296.880 ;
        RECT -22.360 -297.505 -21.515 -297.470 ;
        RECT -22.360 -297.790 -17.370 -297.505 ;
        RECT -16.550 -297.540 -16.250 -297.105 ;
        RECT -15.850 -297.155 -15.620 -296.655 ;
        RECT -15.360 -297.155 -15.130 -296.655 ;
        RECT -14.870 -297.155 -14.640 -296.655 ;
        RECT -14.380 -297.155 -14.150 -296.655 ;
        RECT -13.890 -297.155 -13.660 -296.655 ;
        RECT -13.400 -297.155 -13.170 -296.655 ;
        RECT -11.660 -296.905 -11.415 -296.405 ;
        RECT -11.170 -296.905 -10.940 -296.405 ;
        RECT -10.680 -296.905 -10.450 -296.405 ;
        RECT -10.190 -296.905 -9.960 -296.405 ;
        RECT -9.700 -296.905 -9.470 -296.405 ;
        RECT -9.210 -296.905 -8.980 -296.405 ;
        RECT -8.720 -296.905 -8.490 -296.405 ;
        RECT -8.230 -296.905 -8.000 -296.405 ;
        RECT -7.135 -297.155 -6.905 -296.655 ;
        RECT -6.645 -297.155 -6.415 -296.655 ;
        RECT -6.155 -297.155 -5.925 -296.655 ;
        RECT -5.665 -297.155 -5.435 -296.655 ;
        RECT -5.175 -297.155 -4.945 -296.655 ;
        RECT -4.685 -297.155 -4.455 -296.655 ;
        RECT -8.860 -297.505 -8.015 -297.470 ;
        RECT -4.155 -297.505 -3.870 -295.320 ;
        RECT -3.620 -295.860 -2.960 -295.560 ;
        RECT -3.455 -297.000 -3.165 -295.860 ;
        RECT -1.920 -296.055 -1.445 -295.010 ;
        RECT -2.095 -296.355 -1.410 -296.055 ;
        RECT -22.360 -297.840 -21.515 -297.790 ;
        RECT -29.350 -299.055 -29.120 -298.055 ;
        RECT -28.370 -299.055 -28.140 -298.055 ;
        RECT -27.390 -299.055 -27.160 -298.055 ;
        RECT -25.160 -298.980 -24.930 -298.480 ;
        RECT -24.670 -298.980 -24.440 -298.480 ;
        RECT -24.180 -298.980 -23.950 -298.480 ;
        RECT -23.690 -298.980 -23.460 -298.480 ;
        RECT -23.200 -298.980 -22.970 -298.480 ;
        RECT -22.710 -298.980 -22.480 -298.480 ;
        RECT -22.220 -298.980 -21.990 -298.480 ;
        RECT -21.730 -298.980 -21.500 -298.480 ;
        RECT -20.635 -299.055 -20.405 -298.055 ;
        RECT -19.655 -299.055 -19.425 -298.055 ;
        RECT -18.675 -299.055 -18.445 -298.055 ;
        RECT -17.655 -298.965 -17.370 -297.790 ;
        RECT -8.860 -297.790 -3.870 -297.505 ;
        RECT -3.465 -297.660 -3.165 -297.000 ;
        RECT -2.725 -297.155 -2.495 -296.655 ;
        RECT -2.235 -297.155 -2.005 -296.655 ;
        RECT -1.745 -297.155 -1.515 -296.655 ;
        RECT -1.255 -297.155 -1.025 -296.655 ;
        RECT -0.765 -297.155 -0.535 -296.655 ;
        RECT -0.275 -297.155 -0.045 -296.655 ;
        RECT 1.200 -296.675 1.485 -294.430 ;
        RECT 1.925 -295.430 2.155 -294.430 ;
        RECT 2.415 -295.430 2.645 -294.430 ;
        RECT 3.990 -295.930 4.220 -294.430 ;
        RECT 4.480 -295.930 4.710 -294.430 ;
        RECT 4.970 -295.930 5.200 -294.430 ;
        RECT 5.535 -295.930 5.765 -294.430 ;
        RECT 6.025 -295.930 6.255 -294.430 ;
        RECT 6.515 -295.930 6.745 -294.430 ;
        RECT 7.085 -295.935 7.315 -294.435 ;
        RECT 7.575 -295.935 7.805 -294.435 ;
        RECT 8.065 -295.935 8.295 -294.435 ;
        RECT 1.200 -296.940 1.905 -296.675 ;
        RECT 8.665 -297.495 8.895 -293.470 ;
        RECT 9.430 -294.030 18.175 -293.800 ;
        RECT 9.430 -297.075 9.660 -294.030 ;
        RECT 14.125 -294.535 16.320 -294.300 ;
        RECT 14.125 -296.215 14.355 -294.535 ;
        RECT 9.110 -297.305 9.790 -297.075 ;
        RECT -8.860 -297.840 -8.015 -297.790 ;
        RECT -15.850 -299.055 -15.620 -298.055 ;
        RECT -14.870 -299.055 -14.640 -298.055 ;
        RECT -13.890 -299.055 -13.660 -298.055 ;
        RECT -11.660 -298.980 -11.430 -298.480 ;
        RECT -11.170 -298.980 -10.940 -298.480 ;
        RECT -10.680 -298.980 -10.450 -298.480 ;
        RECT -10.190 -298.980 -9.960 -298.480 ;
        RECT -9.700 -298.980 -9.470 -298.480 ;
        RECT -9.210 -298.980 -8.980 -298.480 ;
        RECT -8.720 -298.980 -8.490 -298.480 ;
        RECT -8.230 -298.980 -8.000 -298.480 ;
        RECT -7.135 -299.055 -6.905 -298.055 ;
        RECT -6.155 -299.055 -5.925 -298.055 ;
        RECT -5.175 -299.055 -4.945 -298.055 ;
        RECT -4.155 -298.965 -3.870 -297.790 ;
        RECT -2.725 -299.055 -2.495 -298.055 ;
        RECT -1.745 -299.055 -1.515 -298.055 ;
        RECT -0.765 -299.055 -0.535 -298.055 ;
        RECT 1.925 -298.970 2.155 -297.970 ;
        RECT 5.615 -298.970 5.845 -297.970 ;
        RECT 6.595 -298.970 6.825 -297.970 ;
        RECT 7.575 -298.970 7.805 -297.970 ;
        RECT 8.665 -298.165 8.935 -297.495 ;
        RECT 11.080 -297.895 11.310 -297.250 ;
        RECT 11.570 -297.750 11.800 -297.250 ;
        RECT 12.060 -297.895 12.290 -297.250 ;
        RECT 12.550 -297.750 12.780 -297.250 ;
        RECT 10.465 -298.125 12.780 -297.895 ;
        RECT 8.705 -298.175 8.935 -298.165 ;
        RECT 10.590 -298.905 10.820 -298.125 ;
        RECT 11.080 -298.135 12.290 -298.125 ;
        RECT 11.570 -298.905 11.800 -298.135 ;
        RECT 12.550 -298.905 12.780 -298.125 ;
        RECT 14.615 -298.900 14.845 -294.715 ;
        RECT 15.105 -296.215 15.335 -294.535 ;
        RECT 15.595 -296.215 15.825 -294.715 ;
        RECT 16.085 -294.720 16.320 -294.535 ;
        RECT 22.150 -294.525 24.345 -294.290 ;
        RECT 16.085 -296.215 16.315 -294.720 ;
        RECT 22.150 -296.205 22.380 -294.525 ;
        RECT 15.595 -298.900 15.825 -297.400 ;
        RECT 19.105 -297.885 19.335 -297.240 ;
        RECT 19.595 -297.740 19.825 -297.240 ;
        RECT 20.085 -297.885 20.315 -297.240 ;
        RECT 20.575 -297.740 20.805 -297.240 ;
        RECT 18.490 -298.115 20.805 -297.885 ;
        RECT 18.615 -298.895 18.845 -298.115 ;
        RECT 19.105 -298.125 20.315 -298.115 ;
        RECT 19.595 -298.895 19.825 -298.125 ;
        RECT 20.575 -298.895 20.805 -298.115 ;
        RECT 22.640 -298.890 22.870 -294.705 ;
        RECT 23.130 -296.205 23.360 -294.525 ;
        RECT 23.620 -296.205 23.850 -294.705 ;
        RECT 24.110 -294.710 24.345 -294.525 ;
        RECT 24.110 -296.205 24.340 -294.710 ;
        RECT 26.735 -295.475 26.965 -294.475 ;
        RECT 27.225 -295.475 27.455 -294.475 ;
        RECT 28.800 -295.975 29.030 -294.475 ;
        RECT 29.290 -295.975 29.520 -294.475 ;
        RECT 29.780 -295.975 30.010 -294.475 ;
        RECT 30.345 -295.975 30.575 -294.475 ;
        RECT 30.835 -295.975 31.065 -294.475 ;
        RECT 31.325 -295.975 31.555 -294.475 ;
        RECT 31.895 -295.980 32.125 -294.480 ;
        RECT 32.385 -295.980 32.615 -294.480 ;
        RECT 32.875 -295.980 33.105 -294.480 ;
        RECT 34.800 -295.930 35.030 -294.930 ;
        RECT 35.290 -295.930 35.520 -294.930 ;
        RECT 36.870 -295.930 37.100 -294.930 ;
        RECT 37.360 -295.930 37.590 -294.930 ;
        RECT 38.680 -295.930 38.910 -294.930 ;
        RECT 39.170 -295.930 39.400 -294.930 ;
        RECT 40.150 -295.930 40.380 -294.930 ;
        RECT 40.640 -295.930 40.870 -294.930 ;
        RECT 41.700 -295.930 41.930 -294.930 ;
        RECT 42.190 -295.930 42.420 -294.930 ;
        RECT 43.245 -295.930 43.475 -294.930 ;
        RECT 43.735 -295.930 43.965 -294.930 ;
        RECT 41.225 -296.120 41.880 -296.090 ;
        RECT 36.455 -296.260 41.880 -296.120 ;
        RECT 34.825 -296.985 35.520 -296.920 ;
        RECT 36.455 -296.985 36.595 -296.260 ;
        RECT 41.225 -296.320 41.880 -296.260 ;
        RECT 34.825 -297.125 36.595 -296.985 ;
        RECT 38.570 -296.855 39.265 -296.770 ;
        RECT 42.755 -296.855 43.435 -296.810 ;
        RECT 38.570 -296.995 43.435 -296.855 ;
        RECT 38.570 -297.040 39.265 -296.995 ;
        RECT 42.755 -297.040 43.435 -296.995 ;
        RECT 34.825 -297.190 35.520 -297.125 ;
        RECT 40.615 -297.180 41.310 -297.140 ;
        RECT 43.690 -297.180 44.385 -297.110 ;
        RECT 40.615 -297.215 44.890 -297.180 ;
        RECT 49.180 -297.215 49.320 -279.535 ;
        RECT 50.855 -292.990 51.110 -274.600 ;
        RECT 50.840 -293.465 51.135 -292.990 ;
        RECT 40.615 -297.320 49.320 -297.215 ;
        RECT 23.620 -298.890 23.850 -297.390 ;
        RECT 40.615 -297.410 41.310 -297.320 ;
        RECT 43.690 -297.355 49.320 -297.320 ;
        RECT 43.690 -297.380 44.385 -297.355 ;
        RECT 32.780 -297.575 33.460 -297.530 ;
        RECT 32.760 -297.805 35.520 -297.575 ;
        RECT 26.735 -299.015 26.965 -298.015 ;
        RECT 30.425 -299.015 30.655 -298.015 ;
        RECT 31.405 -299.015 31.635 -298.015 ;
        RECT 32.385 -299.015 32.615 -298.015 ;
        RECT 34.800 -298.960 35.030 -297.960 ;
        RECT 35.290 -298.960 35.520 -297.805 ;
        RECT 35.780 -298.960 36.010 -297.960 ;
        RECT 36.380 -298.960 36.610 -297.960 ;
        RECT 36.870 -298.960 37.100 -297.960 ;
        RECT 37.360 -298.960 37.590 -297.960 ;
        RECT 39.170 -298.960 39.400 -297.960 ;
        RECT 40.150 -298.960 40.380 -297.960 ;
        RECT 41.700 -298.960 41.930 -297.960 ;
        RECT 43.245 -298.960 43.475 -297.960 ;
        RECT 16.150 -300.925 16.925 -300.915 ;
        RECT -30.355 -300.960 16.925 -300.925 ;
        RECT -30.975 -301.135 16.925 -300.960 ;
        RECT -30.975 -301.190 -30.295 -301.135 ;
        RECT 16.150 -301.145 16.925 -301.135 ;
        RECT -18.575 -301.335 -17.895 -301.325 ;
        RECT -18.575 -301.545 17.350 -301.335 ;
        RECT -18.575 -301.555 -17.895 -301.545 ;
        RECT 16.670 -301.565 17.350 -301.545 ;
        RECT 50.855 -302.140 51.110 -293.465 ;
        RECT -20.050 -302.370 51.110 -302.140 ;
        RECT -20.050 -302.395 48.990 -302.370 ;
        RECT -30.250 -307.185 -30.020 -306.185 ;
        RECT -29.760 -307.185 -29.530 -306.185 ;
        RECT -28.180 -307.185 -27.950 -306.185 ;
        RECT -27.690 -307.185 -27.460 -306.185 ;
        RECT -26.370 -307.185 -26.140 -306.185 ;
        RECT -25.880 -307.185 -25.650 -306.185 ;
        RECT -24.900 -307.185 -24.670 -306.185 ;
        RECT -24.410 -307.185 -24.180 -306.185 ;
        RECT -23.350 -307.185 -23.120 -306.185 ;
        RECT -22.860 -307.185 -22.630 -306.185 ;
        RECT -21.805 -307.185 -21.575 -306.185 ;
        RECT -21.315 -307.185 -21.085 -306.185 ;
        RECT -23.825 -307.375 -23.170 -307.345 ;
        RECT -28.595 -307.515 -23.170 -307.375 ;
        RECT -30.225 -308.240 -29.530 -308.175 ;
        RECT -28.595 -308.240 -28.455 -307.515 ;
        RECT -23.825 -307.575 -23.170 -307.515 ;
        RECT -30.225 -308.380 -28.455 -308.240 ;
        RECT -26.480 -308.110 -25.785 -308.025 ;
        RECT -22.295 -308.110 -21.615 -308.065 ;
        RECT -26.480 -308.250 -21.615 -308.110 ;
        RECT -26.480 -308.295 -25.785 -308.250 ;
        RECT -22.295 -308.295 -21.615 -308.250 ;
        RECT -30.225 -308.445 -29.530 -308.380 ;
        RECT -24.435 -308.435 -23.740 -308.395 ;
        RECT -21.360 -308.435 -20.665 -308.365 ;
        RECT -20.050 -308.435 -19.910 -302.395 ;
        RECT 49.930 -302.550 50.670 -302.510 ;
        RECT 51.285 -302.550 51.465 -274.190 ;
        RECT 51.635 -296.950 51.890 -273.850 ;
        RECT 51.605 -297.645 51.950 -296.950 ;
        RECT -7.625 -302.730 51.465 -302.550 ;
        RECT -18.590 -303.500 -18.360 -302.820 ;
        RECT -18.585 -306.350 -18.365 -303.500 ;
        RECT -18.590 -307.030 -18.360 -306.350 ;
        RECT -17.750 -307.185 -17.520 -306.185 ;
        RECT -17.260 -307.185 -17.030 -306.185 ;
        RECT -15.680 -307.185 -15.450 -306.185 ;
        RECT -15.190 -307.185 -14.960 -306.185 ;
        RECT -13.870 -307.185 -13.640 -306.185 ;
        RECT -13.380 -307.185 -13.150 -306.185 ;
        RECT -12.400 -307.185 -12.170 -306.185 ;
        RECT -11.910 -307.185 -11.680 -306.185 ;
        RECT -10.850 -307.185 -10.620 -306.185 ;
        RECT -10.360 -307.185 -10.130 -306.185 ;
        RECT -9.305 -307.185 -9.075 -306.185 ;
        RECT -8.815 -307.185 -8.585 -306.185 ;
        RECT -11.325 -307.375 -10.670 -307.345 ;
        RECT -16.095 -307.515 -10.670 -307.375 ;
        RECT -24.435 -308.575 -19.910 -308.435 ;
        RECT -17.725 -308.240 -17.030 -308.175 ;
        RECT -16.095 -308.240 -15.955 -307.515 ;
        RECT -11.325 -307.575 -10.670 -307.515 ;
        RECT -15.815 -307.740 -15.120 -307.655 ;
        RECT -10.425 -307.740 -9.730 -307.625 ;
        RECT -15.815 -307.750 -9.730 -307.740 ;
        RECT -7.625 -307.750 -7.485 -302.730 ;
        RECT 49.930 -302.750 50.670 -302.730 ;
        RECT 51.635 -302.890 51.890 -297.645 ;
        RECT -15.815 -307.880 -7.485 -307.750 ;
        RECT -15.815 -307.925 -15.120 -307.880 ;
        RECT -10.425 -307.890 -7.485 -307.880 ;
        RECT -7.195 -303.045 51.890 -302.890 ;
        RECT -7.195 -303.145 48.990 -303.045 ;
        RECT 49.955 -303.080 51.890 -303.045 ;
        RECT -10.425 -307.895 -9.730 -307.890 ;
        RECT -17.725 -308.380 -15.955 -308.240 ;
        RECT -13.980 -308.110 -13.285 -308.025 ;
        RECT -9.795 -308.110 -9.115 -308.065 ;
        RECT -13.980 -308.250 -9.115 -308.110 ;
        RECT -13.980 -308.295 -13.285 -308.250 ;
        RECT -9.795 -308.295 -9.115 -308.250 ;
        RECT -17.725 -308.445 -17.030 -308.380 ;
        RECT -11.935 -308.435 -11.240 -308.395 ;
        RECT -8.860 -308.435 -8.165 -308.365 ;
        RECT -7.195 -308.435 -7.055 -303.145 ;
        RECT 49.130 -303.285 49.845 -303.195 ;
        RECT 52.120 -303.285 52.260 -273.455 ;
        RECT 52.545 -291.390 52.685 -273.170 ;
        RECT 52.445 -291.980 52.765 -291.390 ;
        RECT 4.795 -303.425 52.260 -303.285 ;
        RECT -5.025 -304.925 -4.345 -304.920 ;
        RECT -5.850 -305.145 -4.345 -304.925 ;
        RECT -5.845 -306.330 -5.625 -305.145 ;
        RECT -5.025 -305.150 -4.345 -305.145 ;
        RECT -5.850 -307.010 -5.620 -306.330 ;
        RECT -5.250 -307.185 -5.020 -306.185 ;
        RECT -4.760 -307.185 -4.530 -306.185 ;
        RECT -3.180 -307.185 -2.950 -306.185 ;
        RECT -2.690 -307.185 -2.460 -306.185 ;
        RECT -1.370 -307.185 -1.140 -306.185 ;
        RECT -0.880 -307.185 -0.650 -306.185 ;
        RECT 0.100 -307.185 0.330 -306.185 ;
        RECT 0.590 -307.185 0.820 -306.185 ;
        RECT 1.650 -307.185 1.880 -306.185 ;
        RECT 2.140 -307.185 2.370 -306.185 ;
        RECT 3.195 -307.185 3.425 -306.185 ;
        RECT 3.685 -307.185 3.915 -306.185 ;
        RECT 1.175 -307.375 1.830 -307.345 ;
        RECT -3.595 -307.515 1.830 -307.375 ;
        RECT -11.935 -308.575 -7.055 -308.435 ;
        RECT -5.225 -308.240 -4.530 -308.175 ;
        RECT -3.595 -308.240 -3.455 -307.515 ;
        RECT 1.175 -307.575 1.830 -307.515 ;
        RECT -3.315 -307.740 -2.620 -307.655 ;
        RECT 2.075 -307.740 2.770 -307.625 ;
        RECT -3.315 -307.750 2.770 -307.740 ;
        RECT 4.795 -307.750 4.935 -303.425 ;
        RECT 49.130 -303.430 49.845 -303.425 ;
        RECT 52.545 -303.570 52.685 -291.980 ;
        RECT -3.315 -307.880 4.935 -307.750 ;
        RECT -3.315 -307.925 -2.620 -307.880 ;
        RECT 2.075 -307.890 4.935 -307.880 ;
        RECT 5.165 -303.710 52.685 -303.570 ;
        RECT 2.075 -307.895 2.770 -307.890 ;
        RECT -5.225 -308.380 -3.455 -308.240 ;
        RECT -1.480 -308.110 -0.785 -308.025 ;
        RECT 2.705 -308.110 3.385 -308.065 ;
        RECT -1.480 -308.250 3.385 -308.110 ;
        RECT -1.480 -308.295 -0.785 -308.250 ;
        RECT 2.705 -308.295 3.385 -308.250 ;
        RECT -5.225 -308.445 -4.530 -308.380 ;
        RECT 0.565 -308.435 1.260 -308.395 ;
        RECT 3.640 -308.435 4.335 -308.365 ;
        RECT 5.165 -308.435 5.305 -303.710 ;
        RECT 48.500 -303.885 49.220 -303.850 ;
        RECT 52.930 -303.885 53.070 -272.855 ;
        RECT 17.125 -304.025 53.070 -303.885 ;
        RECT 53.255 -280.205 53.445 -272.535 ;
        RECT 53.255 -280.870 53.505 -280.205 ;
        RECT 7.460 -304.860 8.140 -304.855 ;
        RECT 6.555 -305.080 8.140 -304.860 ;
        RECT 6.555 -306.330 6.775 -305.080 ;
        RECT 7.460 -305.085 8.140 -305.080 ;
        RECT 6.550 -307.010 6.780 -306.330 ;
        RECT 7.250 -307.185 7.480 -306.185 ;
        RECT 7.740 -307.185 7.970 -306.185 ;
        RECT 9.320 -307.185 9.550 -306.185 ;
        RECT 9.810 -307.185 10.040 -306.185 ;
        RECT 11.130 -307.185 11.360 -306.185 ;
        RECT 11.620 -307.185 11.850 -306.185 ;
        RECT 12.600 -307.185 12.830 -306.185 ;
        RECT 13.090 -307.185 13.320 -306.185 ;
        RECT 14.150 -307.185 14.380 -306.185 ;
        RECT 14.640 -307.185 14.870 -306.185 ;
        RECT 15.695 -307.185 15.925 -306.185 ;
        RECT 16.185 -307.185 16.415 -306.185 ;
        RECT 13.675 -307.375 14.330 -307.345 ;
        RECT 8.905 -307.515 14.330 -307.375 ;
        RECT 0.565 -308.575 5.305 -308.435 ;
        RECT 7.275 -308.240 7.970 -308.175 ;
        RECT 8.905 -308.240 9.045 -307.515 ;
        RECT 13.675 -307.575 14.330 -307.515 ;
        RECT 9.185 -307.740 9.880 -307.655 ;
        RECT 14.575 -307.740 15.270 -307.625 ;
        RECT 9.185 -307.750 15.270 -307.740 ;
        RECT 17.125 -307.750 17.265 -304.025 ;
        RECT 48.500 -304.085 49.220 -304.025 ;
        RECT 53.255 -304.205 53.445 -280.870 ;
        RECT 9.185 -307.880 17.265 -307.750 ;
        RECT 9.185 -307.925 9.880 -307.880 ;
        RECT 14.575 -307.890 17.265 -307.880 ;
        RECT 17.540 -304.255 46.030 -304.205 ;
        RECT 49.430 -304.255 53.445 -304.205 ;
        RECT 17.540 -304.395 53.445 -304.255 ;
        RECT 14.575 -307.895 15.270 -307.890 ;
        RECT 7.275 -308.380 9.045 -308.240 ;
        RECT 11.020 -308.110 11.715 -308.025 ;
        RECT 15.205 -308.110 15.885 -308.065 ;
        RECT 11.020 -308.250 15.885 -308.110 ;
        RECT 11.020 -308.295 11.715 -308.250 ;
        RECT 15.205 -308.295 15.885 -308.250 ;
        RECT 7.275 -308.445 7.970 -308.380 ;
        RECT 13.065 -308.435 13.760 -308.395 ;
        RECT 16.140 -308.435 16.835 -308.365 ;
        RECT 17.540 -308.435 17.680 -304.395 ;
        RECT 18.375 -304.770 19.055 -304.540 ;
        RECT 18.640 -306.330 18.860 -304.770 ;
        RECT 32.900 -304.850 33.580 -304.620 ;
        RECT 18.635 -307.010 18.865 -306.330 ;
        RECT 19.750 -307.185 19.980 -306.185 ;
        RECT 20.240 -307.185 20.470 -306.185 ;
        RECT 21.820 -307.185 22.050 -306.185 ;
        RECT 22.310 -307.185 22.540 -306.185 ;
        RECT 23.630 -307.185 23.860 -306.185 ;
        RECT 24.120 -307.185 24.350 -306.185 ;
        RECT 25.100 -307.185 25.330 -306.185 ;
        RECT 25.590 -307.185 25.820 -306.185 ;
        RECT 26.650 -307.185 26.880 -306.185 ;
        RECT 27.140 -307.185 27.370 -306.185 ;
        RECT 28.195 -307.185 28.425 -306.185 ;
        RECT 28.685 -307.185 28.915 -306.185 ;
        RECT 33.165 -306.330 33.385 -304.850 ;
        RECT 54.070 -304.920 54.210 -271.820 ;
        RECT 34.065 -305.060 54.210 -304.920 ;
        RECT 33.160 -307.010 33.390 -306.330 ;
        RECT 26.175 -307.375 26.830 -307.345 ;
        RECT 21.405 -307.515 26.830 -307.375 ;
        RECT 13.065 -308.575 17.680 -308.435 ;
        RECT 19.775 -308.240 20.470 -308.175 ;
        RECT 21.405 -308.240 21.545 -307.515 ;
        RECT 26.175 -307.575 26.830 -307.515 ;
        RECT 19.775 -308.380 21.545 -308.240 ;
        RECT 23.520 -308.110 24.215 -308.025 ;
        RECT 27.705 -308.110 28.385 -308.065 ;
        RECT 23.520 -308.250 28.385 -308.110 ;
        RECT 23.520 -308.295 24.215 -308.250 ;
        RECT 27.705 -308.295 28.385 -308.250 ;
        RECT 19.775 -308.445 20.470 -308.380 ;
        RECT 25.565 -308.435 26.260 -308.395 ;
        RECT 28.640 -308.435 29.335 -308.365 ;
        RECT 34.065 -308.435 34.205 -305.060 ;
        RECT 34.750 -307.185 34.980 -306.185 ;
        RECT 35.240 -307.185 35.470 -306.185 ;
        RECT 36.820 -307.185 37.050 -306.185 ;
        RECT 37.310 -307.185 37.540 -306.185 ;
        RECT 38.630 -307.185 38.860 -306.185 ;
        RECT 39.120 -307.185 39.350 -306.185 ;
        RECT 40.100 -307.185 40.330 -306.185 ;
        RECT 40.590 -307.185 40.820 -306.185 ;
        RECT 41.650 -307.185 41.880 -306.185 ;
        RECT 42.140 -307.185 42.370 -306.185 ;
        RECT 43.195 -307.185 43.425 -306.185 ;
        RECT 43.685 -307.185 43.915 -306.185 ;
        RECT 41.175 -307.375 41.830 -307.345 ;
        RECT 36.405 -307.515 41.830 -307.375 ;
        RECT 25.565 -308.575 34.205 -308.435 ;
        RECT 34.775 -308.240 35.470 -308.175 ;
        RECT 36.405 -308.240 36.545 -307.515 ;
        RECT 41.175 -307.575 41.830 -307.515 ;
        RECT 34.775 -308.380 36.545 -308.240 ;
        RECT 38.520 -308.110 39.215 -308.025 ;
        RECT 42.705 -308.110 43.385 -308.065 ;
        RECT 38.520 -308.250 43.385 -308.110 ;
        RECT 38.520 -308.295 39.215 -308.250 ;
        RECT 42.705 -308.295 43.385 -308.250 ;
        RECT 34.775 -308.445 35.470 -308.380 ;
        RECT 40.565 -308.435 41.260 -308.395 ;
        RECT 43.640 -308.435 44.335 -308.365 ;
        RECT 54.850 -308.435 54.990 -268.305 ;
        RECT 40.565 -308.575 54.990 -308.435 ;
        RECT 58.060 -306.435 59.060 -276.155 ;
        RECT 67.380 -293.865 68.725 -250.735 ;
        RECT 72.340 -255.400 397.965 -253.845 ;
        RECT 67.075 -295.570 69.005 -293.865 ;
        RECT 72.340 -295.315 73.595 -255.400 ;
        RECT 75.275 -257.650 351.625 -256.765 ;
        RECT 75.275 -289.065 76.930 -257.650 ;
        RECT 80.835 -260.445 308.080 -259.340 ;
        RECT 80.835 -280.165 81.285 -260.445 ;
        RECT 87.740 -263.230 262.135 -262.100 ;
        RECT 85.780 -265.630 218.010 -264.305 ;
        RECT 84.370 -267.660 175.605 -266.415 ;
        RECT 84.500 -271.060 87.325 -271.055 ;
        RECT 83.075 -271.760 87.325 -271.060 ;
        RECT 136.500 -273.220 168.825 -272.375 ;
        RECT 82.910 -276.370 84.245 -275.980 ;
        RECT 82.910 -277.145 132.480 -276.370 ;
        RECT 82.910 -277.470 84.245 -277.145 ;
        RECT 84.225 -279.690 88.360 -278.935 ;
        RECT 104.890 -279.605 105.120 -279.105 ;
        RECT 105.380 -279.605 105.610 -279.105 ;
        RECT 105.870 -279.605 106.100 -279.105 ;
        RECT 106.360 -279.605 106.590 -279.105 ;
        RECT 106.850 -279.605 107.080 -279.105 ;
        RECT 107.340 -279.605 107.570 -279.105 ;
        RECT 107.830 -279.605 108.060 -279.105 ;
        RECT 108.320 -279.605 108.550 -279.105 ;
        RECT 109.415 -280.030 109.645 -279.030 ;
        RECT 110.395 -280.030 110.625 -279.030 ;
        RECT 111.375 -280.030 111.605 -279.030 ;
        RECT 80.815 -280.985 81.305 -280.165 ;
        RECT 74.755 -291.190 77.325 -289.065 ;
        RECT 80.835 -291.810 81.285 -280.985 ;
        RECT 94.360 -281.200 94.590 -280.200 ;
        RECT 94.850 -281.200 95.080 -280.200 ;
        RECT 95.340 -281.200 95.570 -280.200 ;
        RECT 95.830 -281.200 96.060 -280.200 ;
        RECT 107.690 -280.295 108.535 -280.245 ;
        RECT 112.395 -280.295 112.680 -279.120 ;
        RECT 113.600 -280.030 113.830 -279.030 ;
        RECT 114.580 -280.030 114.810 -279.030 ;
        RECT 115.560 -280.030 115.790 -279.030 ;
        RECT 118.390 -279.605 118.620 -279.105 ;
        RECT 118.880 -279.605 119.110 -279.105 ;
        RECT 119.370 -279.605 119.600 -279.105 ;
        RECT 119.860 -279.605 120.090 -279.105 ;
        RECT 120.350 -279.605 120.580 -279.105 ;
        RECT 120.840 -279.605 121.070 -279.105 ;
        RECT 121.330 -279.605 121.560 -279.105 ;
        RECT 121.820 -279.605 122.050 -279.105 ;
        RECT 122.915 -280.030 123.145 -279.030 ;
        RECT 123.895 -280.030 124.125 -279.030 ;
        RECT 124.875 -280.030 125.105 -279.030 ;
        RECT 104.410 -280.820 105.180 -280.520 ;
        RECT 107.690 -280.580 112.680 -280.295 ;
        RECT 121.190 -280.295 122.035 -280.245 ;
        RECT 125.895 -280.295 126.180 -279.120 ;
        RECT 127.100 -280.030 127.330 -279.030 ;
        RECT 128.080 -280.030 128.310 -279.030 ;
        RECT 129.060 -280.030 129.290 -279.030 ;
        RECT 116.675 -280.405 116.975 -280.375 ;
        RECT 107.690 -280.615 108.535 -280.580 ;
        RECT 116.260 -280.705 116.975 -280.405 ;
        RECT 117.945 -280.510 118.150 -280.505 ;
        RECT 98.540 -281.390 98.750 -281.370 ;
        RECT 98.130 -281.690 98.790 -281.390 ;
        RECT 94.360 -286.020 94.590 -283.020 ;
        RECT 95.420 -286.020 95.650 -283.020 ;
        RECT 95.910 -286.020 96.140 -283.020 ;
        RECT 96.400 -286.020 96.630 -283.020 ;
        RECT 96.965 -286.020 97.195 -283.020 ;
        RECT 97.455 -286.020 97.685 -283.020 ;
        RECT 97.945 -286.020 98.175 -283.020 ;
        RECT 83.535 -290.705 94.085 -289.725 ;
        RECT 93.105 -290.735 94.085 -290.705 ;
        RECT 93.105 -291.505 94.095 -290.735 ;
        RECT 93.070 -291.715 98.255 -291.505 ;
        RECT 80.835 -291.875 90.750 -291.810 ;
        RECT 80.835 -292.085 97.805 -291.875 ;
        RECT 80.835 -292.260 90.750 -292.085 ;
        RECT 94.335 -294.290 94.565 -293.290 ;
        RECT 94.825 -294.290 95.055 -293.290 ;
        RECT 95.315 -294.290 95.545 -293.290 ;
        RECT 96.385 -294.815 97.045 -294.515 ;
        RECT 72.260 -296.465 73.700 -295.315 ;
        RECT 96.820 -295.380 97.030 -294.815 ;
        RECT 97.595 -294.940 97.805 -292.085 ;
        RECT 98.045 -294.520 98.255 -291.715 ;
        RECT 98.540 -291.860 98.750 -281.690 ;
        RECT 98.990 -281.995 103.540 -281.710 ;
        RECT 98.990 -288.750 99.275 -281.995 ;
        RECT 101.775 -282.575 102.435 -282.275 ;
        RECT 101.875 -283.620 102.350 -282.575 ;
        RECT 103.255 -282.600 103.540 -281.995 ;
        RECT 104.410 -282.195 104.640 -280.820 ;
        RECT 104.890 -281.680 105.120 -281.180 ;
        RECT 105.380 -281.680 105.610 -281.180 ;
        RECT 105.870 -281.680 106.100 -281.180 ;
        RECT 106.360 -281.680 106.590 -281.180 ;
        RECT 106.850 -281.680 107.080 -281.180 ;
        RECT 107.340 -281.680 107.570 -281.180 ;
        RECT 107.830 -281.680 108.060 -281.180 ;
        RECT 108.320 -281.680 108.550 -281.180 ;
        RECT 109.415 -281.430 109.645 -280.930 ;
        RECT 109.905 -281.430 110.135 -280.930 ;
        RECT 110.395 -281.430 110.625 -280.930 ;
        RECT 110.885 -281.430 111.115 -280.930 ;
        RECT 111.375 -281.430 111.605 -280.930 ;
        RECT 111.865 -281.430 112.095 -280.930 ;
        RECT 113.600 -281.430 113.830 -280.930 ;
        RECT 114.090 -281.430 114.320 -280.930 ;
        RECT 114.580 -281.430 114.810 -280.930 ;
        RECT 115.070 -281.430 115.300 -280.930 ;
        RECT 115.560 -281.430 115.790 -280.930 ;
        RECT 116.050 -281.430 116.280 -280.930 ;
        RECT 104.410 -282.420 108.505 -282.195 ;
        RECT 104.450 -282.425 108.505 -282.420 ;
        RECT 103.255 -282.885 104.585 -282.600 ;
        RECT 103.390 -283.425 104.050 -283.125 ;
        RECT 101.840 -283.920 102.525 -283.620 ;
        RECT 100.475 -284.720 100.705 -284.220 ;
        RECT 100.965 -284.720 101.195 -284.220 ;
        RECT 101.455 -284.720 101.685 -284.220 ;
        RECT 101.945 -284.720 102.175 -284.220 ;
        RECT 102.435 -284.720 102.665 -284.220 ;
        RECT 102.925 -284.720 103.155 -284.220 ;
        RECT 103.595 -284.565 103.885 -283.425 ;
        RECT 103.595 -285.225 103.895 -284.565 ;
        RECT 104.300 -285.070 104.585 -282.885 ;
        RECT 108.275 -283.255 108.505 -282.425 ;
        RECT 114.940 -282.575 115.625 -282.275 ;
        RECT 108.275 -283.485 112.075 -283.255 ;
        RECT 108.935 -283.970 109.145 -283.485 ;
        RECT 109.915 -283.970 110.125 -283.485 ;
        RECT 110.890 -283.970 111.100 -283.485 ;
        RECT 111.845 -283.970 112.075 -283.485 ;
        RECT 115.095 -283.615 115.570 -282.575 ;
        RECT 114.975 -283.915 115.660 -283.615 ;
        RECT 104.885 -284.720 105.115 -284.220 ;
        RECT 105.375 -284.720 105.605 -284.220 ;
        RECT 105.865 -284.720 106.095 -284.220 ;
        RECT 106.355 -284.720 106.585 -284.220 ;
        RECT 106.845 -284.720 107.075 -284.220 ;
        RECT 107.335 -284.720 107.565 -284.220 ;
        RECT 108.430 -284.470 108.660 -283.970 ;
        RECT 108.920 -284.470 109.150 -283.970 ;
        RECT 109.410 -284.470 109.640 -283.970 ;
        RECT 109.900 -284.470 110.130 -283.970 ;
        RECT 110.390 -284.470 110.620 -283.970 ;
        RECT 110.880 -284.470 111.110 -283.970 ;
        RECT 111.370 -284.470 111.600 -283.970 ;
        RECT 111.845 -284.470 112.090 -283.970 ;
        RECT 113.600 -284.720 113.830 -284.220 ;
        RECT 114.090 -284.720 114.320 -284.220 ;
        RECT 114.580 -284.720 114.810 -284.220 ;
        RECT 115.070 -284.720 115.300 -284.220 ;
        RECT 115.560 -284.720 115.790 -284.220 ;
        RECT 116.050 -284.720 116.280 -284.220 ;
        RECT 116.675 -284.445 116.975 -280.705 ;
        RECT 117.940 -280.810 118.625 -280.510 ;
        RECT 121.190 -280.580 126.180 -280.295 ;
        RECT 121.190 -280.615 122.035 -280.580 ;
        RECT 117.945 -283.235 118.150 -280.810 ;
        RECT 118.390 -281.680 118.620 -281.180 ;
        RECT 118.880 -281.680 119.110 -281.180 ;
        RECT 119.370 -281.680 119.600 -281.180 ;
        RECT 119.860 -281.680 120.090 -281.180 ;
        RECT 120.350 -281.680 120.580 -281.180 ;
        RECT 120.840 -281.680 121.070 -281.180 ;
        RECT 121.330 -281.680 121.560 -281.180 ;
        RECT 121.820 -281.680 122.050 -281.180 ;
        RECT 122.915 -281.430 123.145 -280.930 ;
        RECT 123.405 -281.430 123.635 -280.930 ;
        RECT 123.895 -281.430 124.125 -280.930 ;
        RECT 124.385 -281.430 124.615 -280.930 ;
        RECT 124.875 -281.430 125.105 -280.930 ;
        RECT 125.365 -281.430 125.595 -280.930 ;
        RECT 126.185 -283.135 126.485 -280.800 ;
        RECT 127.100 -281.430 127.330 -280.930 ;
        RECT 127.590 -281.430 127.820 -280.930 ;
        RECT 128.080 -281.430 128.310 -280.930 ;
        RECT 128.570 -281.430 128.800 -280.930 ;
        RECT 129.060 -281.430 129.290 -280.930 ;
        RECT 129.550 -281.430 129.780 -280.930 ;
        RECT 127.925 -282.545 128.610 -282.245 ;
        RECT 117.945 -283.475 125.600 -283.235 ;
        RECT 126.005 -283.435 126.665 -283.135 ;
        RECT 116.675 -284.670 116.980 -284.445 ;
        RECT 108.445 -285.070 109.290 -285.035 ;
        RECT 104.300 -285.355 109.290 -285.070 ;
        RECT 116.680 -285.105 116.980 -284.670 ;
        RECT 118.385 -284.720 118.615 -284.220 ;
        RECT 118.875 -284.720 119.105 -284.220 ;
        RECT 119.365 -284.720 119.595 -284.220 ;
        RECT 119.855 -284.720 120.085 -284.220 ;
        RECT 120.345 -284.720 120.575 -284.220 ;
        RECT 120.835 -284.720 121.065 -284.220 ;
        RECT 121.930 -284.470 122.160 -283.970 ;
        RECT 122.400 -284.065 122.705 -283.475 ;
        RECT 122.420 -284.470 122.650 -284.065 ;
        RECT 122.910 -284.470 123.140 -283.970 ;
        RECT 123.355 -284.075 123.660 -283.475 ;
        RECT 123.400 -284.470 123.630 -284.075 ;
        RECT 123.890 -284.470 124.120 -283.970 ;
        RECT 124.335 -284.065 124.640 -283.475 ;
        RECT 124.380 -284.470 124.610 -284.065 ;
        RECT 124.870 -284.470 125.100 -283.970 ;
        RECT 125.360 -284.245 125.600 -283.475 ;
        RECT 128.060 -283.635 128.535 -282.545 ;
        RECT 130.050 -282.835 130.350 -282.600 ;
        RECT 130.050 -283.155 131.395 -282.835 ;
        RECT 130.050 -283.285 130.780 -283.155 ;
        RECT 127.995 -283.935 128.655 -283.635 ;
        RECT 125.360 -284.470 125.590 -284.245 ;
        RECT 127.100 -284.720 127.330 -284.220 ;
        RECT 127.590 -284.720 127.820 -284.220 ;
        RECT 128.080 -284.720 128.310 -284.220 ;
        RECT 128.570 -284.720 128.800 -284.220 ;
        RECT 129.060 -284.720 129.290 -284.220 ;
        RECT 129.550 -284.720 129.780 -284.220 ;
        RECT 121.945 -285.070 122.790 -285.035 ;
        RECT 100.965 -286.620 101.195 -285.620 ;
        RECT 101.945 -286.620 102.175 -285.620 ;
        RECT 102.925 -286.620 103.155 -285.620 ;
        RECT 104.300 -286.530 104.585 -285.355 ;
        RECT 108.445 -285.405 109.290 -285.355 ;
        RECT 117.800 -285.355 122.790 -285.070 ;
        RECT 105.375 -286.620 105.605 -285.620 ;
        RECT 106.355 -286.620 106.585 -285.620 ;
        RECT 107.335 -286.620 107.565 -285.620 ;
        RECT 108.430 -286.545 108.660 -286.045 ;
        RECT 108.920 -286.545 109.150 -286.045 ;
        RECT 109.410 -286.545 109.640 -286.045 ;
        RECT 109.900 -286.545 110.130 -286.045 ;
        RECT 110.390 -286.545 110.620 -286.045 ;
        RECT 110.880 -286.545 111.110 -286.045 ;
        RECT 111.370 -286.545 111.600 -286.045 ;
        RECT 111.860 -286.545 112.090 -286.045 ;
        RECT 114.090 -286.620 114.320 -285.620 ;
        RECT 115.070 -286.620 115.300 -285.620 ;
        RECT 116.050 -286.620 116.280 -285.620 ;
        RECT 117.800 -286.530 118.085 -285.355 ;
        RECT 121.945 -285.405 122.790 -285.355 ;
        RECT 118.875 -286.620 119.105 -285.620 ;
        RECT 119.855 -286.620 120.085 -285.620 ;
        RECT 120.835 -286.620 121.065 -285.620 ;
        RECT 121.930 -286.545 122.160 -286.045 ;
        RECT 122.420 -286.545 122.650 -286.045 ;
        RECT 122.910 -286.545 123.140 -286.045 ;
        RECT 123.400 -286.545 123.630 -286.045 ;
        RECT 123.890 -286.545 124.120 -286.045 ;
        RECT 124.380 -286.545 124.610 -286.045 ;
        RECT 124.870 -286.545 125.100 -286.045 ;
        RECT 125.360 -286.545 125.590 -286.045 ;
        RECT 127.590 -286.620 127.820 -285.620 ;
        RECT 128.570 -286.620 128.800 -285.620 ;
        RECT 129.550 -286.620 129.780 -285.620 ;
        RECT 130.330 -287.505 130.780 -283.285 ;
        RECT 110.620 -287.955 130.780 -287.505 ;
        RECT 110.620 -288.410 111.420 -287.955 ;
        RECT 98.990 -289.035 115.350 -288.750 ;
        RECT 110.605 -289.985 111.405 -289.325 ;
        RECT 98.540 -292.070 102.390 -291.860 ;
        RECT 110.090 -291.900 110.750 -291.600 ;
        RECT 99.065 -294.290 99.295 -293.290 ;
        RECT 99.555 -294.290 99.785 -293.290 ;
        RECT 100.045 -294.290 100.275 -293.290 ;
        RECT 98.625 -294.520 99.285 -294.485 ;
        RECT 98.045 -294.730 99.285 -294.520 ;
        RECT 98.625 -294.785 99.285 -294.730 ;
        RECT 99.740 -294.940 100.400 -294.885 ;
        RECT 97.595 -295.150 100.400 -294.940 ;
        RECT 99.740 -295.185 100.400 -295.150 ;
        RECT 101.565 -295.380 101.865 -295.230 ;
        RECT 96.820 -295.590 101.865 -295.380 ;
        RECT 94.335 -297.750 94.565 -295.750 ;
        RECT 95.390 -297.750 95.620 -295.750 ;
        RECT 95.880 -297.750 96.110 -295.750 ;
        RECT 96.370 -297.750 96.600 -295.750 ;
        RECT 99.065 -297.750 99.295 -295.750 ;
        RECT 100.120 -297.750 100.350 -295.750 ;
        RECT 100.610 -297.750 100.840 -295.750 ;
        RECT 101.100 -297.750 101.330 -295.750 ;
        RECT 101.565 -295.890 101.865 -295.590 ;
        RECT 102.180 -296.480 102.390 -292.070 ;
        RECT 103.155 -294.885 103.385 -293.385 ;
        RECT 103.645 -294.885 103.875 -293.385 ;
        RECT 104.135 -294.885 104.365 -293.385 ;
        RECT 104.705 -294.880 104.935 -293.380 ;
        RECT 105.195 -294.880 105.425 -293.380 ;
        RECT 105.685 -294.880 105.915 -293.380 ;
        RECT 106.250 -294.880 106.480 -293.380 ;
        RECT 106.740 -294.880 106.970 -293.380 ;
        RECT 107.230 -294.880 107.460 -293.380 ;
        RECT 108.805 -294.380 109.035 -293.380 ;
        RECT 109.295 -294.380 109.525 -293.380 ;
        RECT 110.250 -295.325 110.550 -291.900 ;
        RECT 110.945 -292.105 111.245 -289.985 ;
        RECT 113.190 -291.380 113.420 -289.380 ;
        RECT 114.170 -291.380 114.400 -289.380 ;
        RECT 115.065 -291.645 115.350 -289.035 ;
        RECT 131.705 -289.090 132.480 -277.145 ;
        RECT 116.045 -289.440 132.480 -289.090 ;
        RECT 116.045 -290.335 116.395 -289.440 ;
        RECT 110.945 -292.110 112.650 -292.105 ;
        RECT 110.945 -292.400 112.655 -292.110 ;
        RECT 114.920 -292.315 115.350 -291.645 ;
        RECT 110.945 -292.405 112.650 -292.400 ;
        RECT 110.055 -295.625 110.710 -295.325 ;
        RECT 110.945 -296.175 111.245 -292.405 ;
        RECT 112.700 -293.650 112.930 -292.650 ;
        RECT 113.190 -293.650 113.420 -292.650 ;
        RECT 113.750 -293.650 113.980 -292.650 ;
        RECT 114.240 -293.650 114.470 -292.650 ;
        RECT 116.850 -293.105 117.080 -289.605 ;
        RECT 117.340 -293.105 117.570 -289.605 ;
        RECT 118.850 -293.105 119.080 -289.605 ;
        RECT 119.340 -293.105 119.570 -289.605 ;
        RECT 121.265 -293.090 121.615 -289.440 ;
        RECT 121.850 -293.105 122.080 -289.605 ;
        RECT 122.340 -293.105 122.570 -289.605 ;
        RECT 123.850 -293.105 124.080 -289.605 ;
        RECT 124.340 -293.105 124.570 -289.605 ;
        RECT 126.220 -293.095 126.570 -289.440 ;
        RECT 126.850 -293.105 127.080 -289.605 ;
        RECT 127.340 -293.105 127.570 -289.605 ;
        RECT 128.850 -293.105 129.080 -289.605 ;
        RECT 129.340 -293.105 129.570 -289.605 ;
        RECT 136.500 -291.460 137.345 -273.220 ;
        RECT 146.625 -274.545 148.820 -274.310 ;
        RECT 146.625 -274.730 146.860 -274.545 ;
        RECT 140.825 -277.095 141.475 -276.345 ;
        RECT 142.255 -276.615 142.485 -275.615 ;
        RECT 142.745 -276.755 142.975 -275.615 ;
        RECT 143.235 -276.615 143.465 -275.615 ;
        RECT 143.725 -276.755 143.955 -275.615 ;
        RECT 146.630 -276.225 146.860 -274.730 ;
        RECT 147.120 -276.225 147.350 -274.725 ;
        RECT 147.610 -276.225 147.840 -274.545 ;
        RECT 142.255 -276.985 145.440 -276.755 ;
        RECT 141.075 -284.115 141.345 -277.095 ;
        RECT 142.255 -278.265 142.485 -276.985 ;
        RECT 142.745 -276.995 143.955 -276.985 ;
        RECT 143.235 -278.265 143.465 -276.995 ;
        RECT 144.215 -278.265 144.445 -276.985 ;
        RECT 147.120 -278.910 147.350 -277.410 ;
        RECT 148.100 -278.910 148.330 -274.725 ;
        RECT 148.590 -276.225 148.820 -274.545 ;
        RECT 152.100 -277.085 155.640 -276.520 ;
        RECT 150.165 -277.760 150.395 -277.260 ;
        RECT 150.655 -277.905 150.885 -277.260 ;
        RECT 151.145 -277.760 151.375 -277.260 ;
        RECT 151.635 -277.905 151.865 -277.260 ;
        RECT 150.165 -278.135 153.350 -277.905 ;
        RECT 150.165 -278.915 150.395 -278.135 ;
        RECT 150.655 -278.145 151.865 -278.135 ;
        RECT 151.145 -278.915 151.375 -278.145 ;
        RECT 152.125 -278.915 152.355 -278.135 ;
        RECT 142.125 -283.410 142.355 -281.910 ;
        RECT 140.360 -284.385 141.345 -284.115 ;
        RECT 141.635 -286.090 141.865 -284.595 ;
        RECT 141.630 -286.275 141.865 -286.090 ;
        RECT 142.125 -286.095 142.355 -284.595 ;
        RECT 142.615 -286.275 142.845 -284.595 ;
        RECT 143.105 -286.095 143.335 -281.910 ;
        RECT 145.170 -282.685 145.400 -281.905 ;
        RECT 146.150 -282.675 146.380 -281.905 ;
        RECT 145.660 -282.685 146.870 -282.675 ;
        RECT 147.130 -282.685 147.360 -281.905 ;
        RECT 145.170 -282.915 148.355 -282.685 ;
        RECT 145.170 -283.560 145.400 -283.060 ;
        RECT 145.660 -283.560 145.890 -282.915 ;
        RECT 146.150 -283.560 146.380 -283.060 ;
        RECT 146.640 -283.560 146.870 -282.915 ;
        RECT 149.360 -284.465 149.590 -281.465 ;
        RECT 150.415 -284.465 150.645 -281.465 ;
        RECT 150.905 -284.465 151.135 -281.465 ;
        RECT 151.395 -284.465 151.625 -281.465 ;
        RECT 152.455 -284.465 152.685 -281.465 ;
        RECT 143.595 -286.275 143.825 -284.595 ;
        RECT 153.610 -285.120 154.135 -284.760 ;
        RECT 153.640 -285.535 153.965 -285.120 ;
        RECT 148.865 -285.860 153.965 -285.535 ;
        RECT 141.630 -286.510 143.825 -286.275 ;
        RECT 149.360 -287.525 149.590 -286.025 ;
        RECT 149.850 -287.525 150.080 -286.025 ;
        RECT 150.340 -287.525 150.570 -286.025 ;
        RECT 151.550 -287.525 151.780 -286.025 ;
        RECT 152.040 -287.525 152.270 -286.025 ;
        RECT 153.205 -288.065 153.770 -288.060 ;
        RECT 155.075 -288.065 155.640 -277.085 ;
        RECT 159.320 -283.255 159.550 -280.755 ;
        RECT 160.665 -283.255 160.895 -280.755 ;
        RECT 161.155 -283.255 161.385 -280.755 ;
        RECT 161.645 -283.255 161.875 -280.755 ;
        RECT 162.295 -283.255 162.525 -280.755 ;
        RECT 163.925 -283.255 164.155 -280.755 ;
        RECT 165.065 -282.255 165.295 -280.755 ;
        RECT 158.165 -284.055 158.855 -284.035 ;
        RECT 162.195 -284.055 162.885 -284.035 ;
        RECT 164.120 -284.055 164.390 -283.690 ;
        RECT 158.165 -284.275 164.390 -284.055 ;
        RECT 158.165 -284.305 158.855 -284.275 ;
        RECT 162.195 -284.305 162.885 -284.275 ;
        RECT 164.120 -284.380 164.390 -284.275 ;
        RECT 164.980 -284.455 165.310 -284.395 ;
        RECT 167.980 -284.455 168.825 -273.220 ;
        RECT 174.360 -273.830 175.605 -267.660 ;
        RECT 176.415 -272.960 211.825 -272.005 ;
        RECT 173.905 -274.510 175.690 -273.830 ;
        RECT 173.905 -274.780 175.720 -274.510 ;
        RECT 173.905 -275.165 175.690 -274.780 ;
        RECT 157.360 -285.990 157.875 -285.535 ;
        RECT 152.255 -288.630 155.640 -288.065 ;
        RECT 136.500 -291.890 138.250 -291.460 ;
        RECT 146.585 -291.810 148.780 -291.575 ;
        RECT 136.500 -292.160 145.140 -291.890 ;
        RECT 146.585 -291.995 146.820 -291.810 ;
        RECT 136.500 -292.305 138.250 -292.160 ;
        RECT 119.910 -293.355 120.500 -293.295 ;
        RECT 119.910 -293.525 120.945 -293.355 ;
        RECT 129.775 -293.390 130.365 -293.370 ;
        RECT 132.530 -293.390 133.135 -293.275 ;
        RECT 119.910 -293.585 120.500 -293.525 ;
        RECT 112.450 -295.985 112.680 -295.485 ;
        RECT 112.940 -295.985 113.170 -295.485 ;
        RECT 113.430 -295.985 113.660 -295.485 ;
        RECT 113.920 -295.985 114.150 -295.485 ;
        RECT 114.410 -295.985 114.640 -295.485 ;
        RECT 114.900 -295.985 115.130 -295.485 ;
        RECT 110.945 -296.475 112.580 -296.175 ;
        RECT 102.140 -297.140 102.440 -296.480 ;
        RECT 103.645 -297.920 103.875 -296.920 ;
        RECT 104.625 -297.920 104.855 -296.920 ;
        RECT 105.605 -297.920 105.835 -296.920 ;
        RECT 109.295 -297.920 109.525 -296.920 ;
        RECT 112.940 -297.885 113.170 -296.885 ;
        RECT 113.920 -297.885 114.150 -296.885 ;
        RECT 114.900 -297.885 115.130 -296.885 ;
        RECT 117.340 -297.530 117.570 -294.030 ;
        RECT 119.340 -297.530 119.570 -294.030 ;
        RECT 120.775 -298.030 120.945 -293.525 ;
        RECT 125.295 -293.720 125.885 -293.430 ;
        RECT 129.775 -293.615 133.135 -293.390 ;
        RECT 129.775 -293.660 130.365 -293.615 ;
        RECT 122.340 -297.530 122.570 -294.030 ;
        RECT 124.340 -297.530 124.570 -294.030 ;
        RECT 125.325 -297.705 125.495 -293.720 ;
        RECT 127.340 -297.530 127.570 -294.030 ;
        RECT 129.340 -297.530 129.570 -294.030 ;
        RECT 125.325 -297.875 131.865 -297.705 ;
        RECT 120.775 -298.200 131.425 -298.030 ;
        RECT 60.325 -302.810 60.555 -301.810 ;
        RECT 61.305 -302.810 61.535 -301.810 ;
        RECT 62.285 -302.810 62.515 -301.810 ;
        RECT 63.660 -303.075 63.945 -301.900 ;
        RECT 64.735 -302.810 64.965 -301.810 ;
        RECT 65.715 -302.810 65.945 -301.810 ;
        RECT 66.695 -302.810 66.925 -301.810 ;
        RECT 67.790 -302.385 68.020 -301.885 ;
        RECT 68.280 -302.385 68.510 -301.885 ;
        RECT 68.770 -302.385 69.000 -301.885 ;
        RECT 69.260 -302.385 69.490 -301.885 ;
        RECT 69.750 -302.385 69.980 -301.885 ;
        RECT 70.240 -302.385 70.470 -301.885 ;
        RECT 70.730 -302.385 70.960 -301.885 ;
        RECT 71.220 -302.385 71.450 -301.885 ;
        RECT 73.450 -302.810 73.680 -301.810 ;
        RECT 74.430 -302.810 74.660 -301.810 ;
        RECT 75.410 -302.810 75.640 -301.810 ;
        RECT 67.805 -303.075 68.650 -303.025 ;
        RECT 59.835 -304.210 60.065 -303.710 ;
        RECT 60.325 -304.210 60.555 -303.710 ;
        RECT 60.815 -304.210 61.045 -303.710 ;
        RECT 61.305 -304.210 61.535 -303.710 ;
        RECT 61.795 -304.210 62.025 -303.710 ;
        RECT 62.285 -304.210 62.515 -303.710 ;
        RECT 62.955 -303.865 63.255 -303.205 ;
        RECT 63.660 -303.360 68.650 -303.075 ;
        RECT 77.160 -303.075 77.445 -301.900 ;
        RECT 78.235 -302.810 78.465 -301.810 ;
        RECT 79.215 -302.810 79.445 -301.810 ;
        RECT 80.195 -302.810 80.425 -301.810 ;
        RECT 81.290 -302.385 81.520 -301.885 ;
        RECT 81.780 -302.385 82.010 -301.885 ;
        RECT 82.270 -302.385 82.500 -301.885 ;
        RECT 82.760 -302.385 82.990 -301.885 ;
        RECT 83.250 -302.385 83.480 -301.885 ;
        RECT 83.740 -302.385 83.970 -301.885 ;
        RECT 84.230 -302.385 84.460 -301.885 ;
        RECT 84.720 -302.385 84.950 -301.885 ;
        RECT 86.950 -302.810 87.180 -301.810 ;
        RECT 87.930 -302.810 88.160 -301.810 ;
        RECT 88.910 -302.810 89.140 -301.810 ;
        RECT 81.305 -303.075 82.150 -303.025 ;
        RECT 61.200 -304.810 61.885 -304.510 ;
        RECT 61.235 -305.855 61.710 -304.810 ;
        RECT 62.955 -305.005 63.245 -303.865 ;
        RECT 62.750 -305.305 63.410 -305.005 ;
        RECT 63.660 -305.545 63.945 -303.360 ;
        RECT 67.805 -303.395 68.650 -303.360 ;
        RECT 64.245 -304.210 64.475 -303.710 ;
        RECT 64.735 -304.210 64.965 -303.710 ;
        RECT 65.225 -304.210 65.455 -303.710 ;
        RECT 65.715 -304.210 65.945 -303.710 ;
        RECT 66.205 -304.210 66.435 -303.710 ;
        RECT 66.695 -304.210 66.925 -303.710 ;
        RECT 67.790 -304.460 68.020 -303.960 ;
        RECT 68.280 -304.460 68.510 -303.960 ;
        RECT 68.770 -304.460 69.000 -303.960 ;
        RECT 69.260 -304.460 69.490 -303.960 ;
        RECT 69.750 -304.460 69.980 -303.960 ;
        RECT 70.240 -304.460 70.470 -303.960 ;
        RECT 70.730 -304.460 70.960 -303.960 ;
        RECT 71.205 -304.460 71.450 -303.960 ;
        RECT 72.960 -304.210 73.190 -303.710 ;
        RECT 73.450 -304.210 73.680 -303.710 ;
        RECT 73.940 -304.210 74.170 -303.710 ;
        RECT 74.430 -304.210 74.660 -303.710 ;
        RECT 74.920 -304.210 75.150 -303.710 ;
        RECT 75.410 -304.210 75.640 -303.710 ;
        RECT 76.040 -303.760 76.340 -303.325 ;
        RECT 77.160 -303.360 82.150 -303.075 ;
        RECT 81.305 -303.395 82.150 -303.360 ;
        RECT 76.035 -303.985 76.340 -303.760 ;
        RECT 68.295 -304.945 68.505 -304.460 ;
        RECT 69.275 -304.945 69.485 -304.460 ;
        RECT 70.250 -304.945 70.460 -304.460 ;
        RECT 71.205 -304.945 71.435 -304.460 ;
        RECT 74.335 -304.815 75.020 -304.515 ;
        RECT 62.615 -305.830 63.945 -305.545 ;
        RECT 67.635 -305.175 71.435 -304.945 ;
        RECT 61.135 -306.155 61.795 -305.855 ;
        RECT 62.615 -306.435 62.900 -305.830 ;
        RECT 67.635 -306.005 67.865 -305.175 ;
        RECT 74.455 -305.855 74.930 -304.815 ;
        RECT 63.810 -306.010 67.865 -306.005 ;
        RECT 58.060 -306.720 62.900 -306.435 ;
        RECT 63.770 -306.235 67.865 -306.010 ;
        RECT 74.300 -306.155 74.985 -305.855 ;
        RECT -24.435 -308.665 -23.740 -308.575 ;
        RECT -21.360 -308.635 -20.665 -308.575 ;
        RECT -11.935 -308.665 -11.240 -308.575 ;
        RECT -8.860 -308.635 -8.165 -308.575 ;
        RECT 0.565 -308.665 1.260 -308.575 ;
        RECT 3.640 -308.635 4.335 -308.575 ;
        RECT 13.065 -308.665 13.760 -308.575 ;
        RECT 16.140 -308.635 16.835 -308.575 ;
        RECT 25.565 -308.665 26.260 -308.575 ;
        RECT 28.640 -308.635 29.335 -308.575 ;
        RECT 40.565 -308.665 41.260 -308.575 ;
        RECT 43.640 -308.635 44.335 -308.575 ;
        RECT -30.250 -310.215 -30.020 -309.215 ;
        RECT -29.760 -310.215 -29.530 -309.215 ;
        RECT -29.270 -310.215 -29.040 -309.215 ;
        RECT -28.670 -310.215 -28.440 -309.215 ;
        RECT -28.180 -310.215 -27.950 -309.215 ;
        RECT -27.690 -310.215 -27.460 -309.215 ;
        RECT -25.880 -310.215 -25.650 -309.215 ;
        RECT -24.900 -310.215 -24.670 -309.215 ;
        RECT -23.350 -310.215 -23.120 -309.215 ;
        RECT -21.805 -310.215 -21.575 -309.215 ;
        RECT -17.750 -310.215 -17.520 -309.215 ;
        RECT -17.260 -310.215 -17.030 -309.215 ;
        RECT -16.770 -310.215 -16.540 -309.215 ;
        RECT -16.170 -310.215 -15.940 -309.215 ;
        RECT -15.680 -310.215 -15.450 -309.215 ;
        RECT -15.190 -310.215 -14.960 -309.215 ;
        RECT -13.380 -310.215 -13.150 -309.215 ;
        RECT -12.400 -310.215 -12.170 -309.215 ;
        RECT -10.850 -310.215 -10.620 -309.215 ;
        RECT -9.305 -310.215 -9.075 -309.215 ;
        RECT -5.250 -310.215 -5.020 -309.215 ;
        RECT -4.760 -310.215 -4.530 -309.215 ;
        RECT -4.270 -310.215 -4.040 -309.215 ;
        RECT -3.670 -310.215 -3.440 -309.215 ;
        RECT -3.180 -310.215 -2.950 -309.215 ;
        RECT -2.690 -310.215 -2.460 -309.215 ;
        RECT -0.880 -310.215 -0.650 -309.215 ;
        RECT 0.100 -310.215 0.330 -309.215 ;
        RECT 1.650 -310.215 1.880 -309.215 ;
        RECT 3.195 -310.215 3.425 -309.215 ;
        RECT 7.250 -310.215 7.480 -309.215 ;
        RECT 7.740 -310.215 7.970 -309.215 ;
        RECT 8.230 -310.215 8.460 -309.215 ;
        RECT 8.830 -310.215 9.060 -309.215 ;
        RECT 9.320 -310.215 9.550 -309.215 ;
        RECT 9.810 -310.215 10.040 -309.215 ;
        RECT 11.620 -310.215 11.850 -309.215 ;
        RECT 12.600 -310.215 12.830 -309.215 ;
        RECT 14.150 -310.215 14.380 -309.215 ;
        RECT 15.695 -310.215 15.925 -309.215 ;
        RECT 19.750 -310.215 19.980 -309.215 ;
        RECT 20.240 -310.215 20.470 -309.215 ;
        RECT 20.730 -310.215 20.960 -309.215 ;
        RECT 21.330 -310.215 21.560 -309.215 ;
        RECT 21.820 -310.215 22.050 -309.215 ;
        RECT 22.310 -310.215 22.540 -309.215 ;
        RECT 24.120 -310.215 24.350 -309.215 ;
        RECT 25.100 -310.215 25.330 -309.215 ;
        RECT 26.650 -310.215 26.880 -309.215 ;
        RECT 28.195 -310.215 28.425 -309.215 ;
        RECT 34.750 -310.215 34.980 -309.215 ;
        RECT 35.240 -310.215 35.470 -309.215 ;
        RECT 35.730 -310.215 35.960 -309.215 ;
        RECT 36.330 -310.215 36.560 -309.215 ;
        RECT 36.820 -310.215 37.050 -309.215 ;
        RECT 37.310 -310.215 37.540 -309.215 ;
        RECT 39.120 -310.215 39.350 -309.215 ;
        RECT 40.100 -310.215 40.330 -309.215 ;
        RECT 41.650 -310.215 41.880 -309.215 ;
        RECT 43.195 -310.215 43.425 -309.215 ;
        RECT -91.515 -311.940 -90.825 -311.255 ;
        RECT -33.040 -312.030 -32.225 -311.155 ;
        RECT -92.205 -312.430 -91.520 -312.140 ;
        RECT -108.645 -321.950 -108.030 -321.335 ;
        RECT -32.985 -323.805 -32.325 -312.030 ;
        RECT 48.340 -317.970 48.645 -311.085 ;
        RECT 47.995 -317.975 48.645 -317.970 ;
        RECT 47.995 -318.140 48.650 -317.975 ;
        RECT 48.000 -318.565 48.650 -318.140 ;
        RECT 48.910 -318.610 49.230 -311.065 ;
        RECT 48.900 -319.470 49.230 -318.610 ;
        RECT 48.795 -319.475 49.230 -319.470 ;
        RECT 48.795 -320.090 49.410 -319.475 ;
        RECT 49.635 -321.310 49.935 -310.885 ;
        RECT 49.550 -321.925 50.165 -321.310 ;
        RECT -32.985 -324.485 -32.305 -323.805 ;
        RECT 58.060 -325.670 59.060 -306.720 ;
        RECT 63.770 -307.610 64.000 -306.235 ;
        RECT 64.250 -307.250 64.480 -306.750 ;
        RECT 64.740 -307.250 64.970 -306.750 ;
        RECT 65.230 -307.250 65.460 -306.750 ;
        RECT 65.720 -307.250 65.950 -306.750 ;
        RECT 66.210 -307.250 66.440 -306.750 ;
        RECT 66.700 -307.250 66.930 -306.750 ;
        RECT 67.190 -307.250 67.420 -306.750 ;
        RECT 67.680 -307.250 67.910 -306.750 ;
        RECT 68.775 -307.500 69.005 -307.000 ;
        RECT 69.265 -307.500 69.495 -307.000 ;
        RECT 69.755 -307.500 69.985 -307.000 ;
        RECT 70.245 -307.500 70.475 -307.000 ;
        RECT 70.735 -307.500 70.965 -307.000 ;
        RECT 71.225 -307.500 71.455 -307.000 ;
        RECT 72.960 -307.500 73.190 -307.000 ;
        RECT 73.450 -307.500 73.680 -307.000 ;
        RECT 73.940 -307.500 74.170 -307.000 ;
        RECT 74.430 -307.500 74.660 -307.000 ;
        RECT 74.920 -307.500 75.150 -307.000 ;
        RECT 75.410 -307.500 75.640 -307.000 ;
        RECT 63.770 -307.910 64.540 -307.610 ;
        RECT 76.035 -307.725 76.335 -303.985 ;
        RECT 77.745 -304.210 77.975 -303.710 ;
        RECT 78.235 -304.210 78.465 -303.710 ;
        RECT 78.725 -304.210 78.955 -303.710 ;
        RECT 79.215 -304.210 79.445 -303.710 ;
        RECT 79.705 -304.210 79.935 -303.710 ;
        RECT 80.195 -304.210 80.425 -303.710 ;
        RECT 81.290 -304.460 81.520 -303.960 ;
        RECT 81.780 -304.365 82.010 -303.960 ;
        RECT 81.760 -304.955 82.065 -304.365 ;
        RECT 82.270 -304.460 82.500 -303.960 ;
        RECT 82.760 -304.355 82.990 -303.960 ;
        RECT 82.715 -304.955 83.020 -304.355 ;
        RECT 83.250 -304.460 83.480 -303.960 ;
        RECT 83.740 -304.365 83.970 -303.960 ;
        RECT 83.695 -304.955 84.000 -304.365 ;
        RECT 84.230 -304.460 84.460 -303.960 ;
        RECT 84.720 -304.185 84.950 -303.960 ;
        RECT 84.720 -304.955 84.960 -304.185 ;
        RECT 86.460 -304.210 86.690 -303.710 ;
        RECT 86.950 -304.210 87.180 -303.710 ;
        RECT 87.440 -304.210 87.670 -303.710 ;
        RECT 87.930 -304.210 88.160 -303.710 ;
        RECT 88.420 -304.210 88.650 -303.710 ;
        RECT 88.910 -304.210 89.140 -303.710 ;
        RECT 87.355 -304.795 88.015 -304.495 ;
        RECT 77.305 -305.195 84.960 -304.955 ;
        RECT 77.305 -307.620 77.510 -305.195 ;
        RECT 85.365 -305.295 86.025 -304.995 ;
        RECT 77.750 -307.250 77.980 -306.750 ;
        RECT 78.240 -307.250 78.470 -306.750 ;
        RECT 78.730 -307.250 78.960 -306.750 ;
        RECT 79.220 -307.250 79.450 -306.750 ;
        RECT 79.710 -307.250 79.940 -306.750 ;
        RECT 80.200 -307.250 80.430 -306.750 ;
        RECT 80.690 -307.250 80.920 -306.750 ;
        RECT 81.180 -307.250 81.410 -306.750 ;
        RECT 82.275 -307.500 82.505 -307.000 ;
        RECT 82.765 -307.500 82.995 -307.000 ;
        RECT 83.255 -307.500 83.485 -307.000 ;
        RECT 83.745 -307.500 83.975 -307.000 ;
        RECT 84.235 -307.500 84.465 -307.000 ;
        RECT 84.725 -307.500 84.955 -307.000 ;
        RECT 67.050 -307.850 67.895 -307.815 ;
        RECT 67.050 -308.135 72.040 -307.850 ;
        RECT 75.620 -308.025 76.335 -307.725 ;
        RECT 77.300 -307.920 77.985 -307.620 ;
        RECT 85.545 -307.630 85.845 -305.295 ;
        RECT 87.420 -305.885 87.895 -304.795 ;
        RECT 89.410 -305.275 89.710 -305.145 ;
        RECT 89.410 -305.595 91.690 -305.275 ;
        RECT 89.410 -305.830 89.710 -305.595 ;
        RECT 87.285 -306.185 87.970 -305.885 ;
        RECT 86.460 -307.500 86.690 -307.000 ;
        RECT 86.950 -307.500 87.180 -307.000 ;
        RECT 87.440 -307.500 87.670 -307.000 ;
        RECT 87.930 -307.500 88.160 -307.000 ;
        RECT 88.420 -307.500 88.650 -307.000 ;
        RECT 88.910 -307.500 89.140 -307.000 ;
        RECT 80.550 -307.850 81.395 -307.815 ;
        RECT 77.305 -307.925 77.510 -307.920 ;
        RECT 76.035 -308.055 76.335 -308.025 ;
        RECT 67.050 -308.185 67.895 -308.135 ;
        RECT 64.250 -309.325 64.480 -308.825 ;
        RECT 64.740 -309.325 64.970 -308.825 ;
        RECT 65.230 -309.325 65.460 -308.825 ;
        RECT 65.720 -309.325 65.950 -308.825 ;
        RECT 66.210 -309.325 66.440 -308.825 ;
        RECT 66.700 -309.325 66.930 -308.825 ;
        RECT 67.190 -309.325 67.420 -308.825 ;
        RECT 67.680 -309.325 67.910 -308.825 ;
        RECT 68.775 -309.400 69.005 -308.400 ;
        RECT 69.755 -309.400 69.985 -308.400 ;
        RECT 70.735 -309.400 70.965 -308.400 ;
        RECT 71.755 -309.310 72.040 -308.135 ;
        RECT 80.550 -308.135 85.540 -307.850 ;
        RECT 80.550 -308.185 81.395 -308.135 ;
        RECT 72.960 -309.400 73.190 -308.400 ;
        RECT 73.940 -309.400 74.170 -308.400 ;
        RECT 74.920 -309.400 75.150 -308.400 ;
        RECT 77.750 -309.325 77.980 -308.825 ;
        RECT 78.240 -309.325 78.470 -308.825 ;
        RECT 78.730 -309.325 78.960 -308.825 ;
        RECT 79.220 -309.325 79.450 -308.825 ;
        RECT 79.710 -309.325 79.940 -308.825 ;
        RECT 80.200 -309.325 80.430 -308.825 ;
        RECT 80.690 -309.325 80.920 -308.825 ;
        RECT 81.180 -309.325 81.410 -308.825 ;
        RECT 82.275 -309.400 82.505 -308.400 ;
        RECT 83.255 -309.400 83.485 -308.400 ;
        RECT 84.235 -309.400 84.465 -308.400 ;
        RECT 85.255 -309.310 85.540 -308.135 ;
        RECT 86.460 -309.400 86.690 -308.400 ;
        RECT 87.440 -309.400 87.670 -308.400 ;
        RECT 88.420 -309.400 88.650 -308.400 ;
        RECT 91.050 -323.805 91.690 -305.595 ;
        RECT 128.560 -309.055 128.910 -298.200 ;
        RECT 131.695 -298.515 131.865 -297.875 ;
        RECT 127.965 -310.155 129.820 -309.055 ;
        RECT 131.390 -311.800 131.995 -298.515 ;
        RECT 91.025 -324.485 91.690 -323.805 ;
        RECT 124.990 -312.405 131.995 -311.800 ;
        RECT 124.990 -326.620 125.595 -312.405 ;
        RECT 132.530 -323.610 133.135 -293.615 ;
        RECT 140.785 -294.360 141.435 -293.610 ;
        RECT 142.215 -293.880 142.445 -292.880 ;
        RECT 142.705 -294.020 142.935 -292.880 ;
        RECT 143.195 -293.880 143.425 -292.880 ;
        RECT 143.685 -294.020 143.915 -292.880 ;
        RECT 144.870 -293.610 145.140 -292.160 ;
        RECT 146.590 -293.490 146.820 -291.995 ;
        RECT 147.080 -293.490 147.310 -291.990 ;
        RECT 147.570 -293.490 147.800 -291.810 ;
        RECT 144.870 -293.880 146.510 -293.610 ;
        RECT 142.215 -294.250 145.400 -294.020 ;
        RECT 146.240 -294.155 146.510 -293.880 ;
        RECT 141.035 -301.380 141.305 -294.360 ;
        RECT 142.215 -295.530 142.445 -294.250 ;
        RECT 142.705 -294.260 143.915 -294.250 ;
        RECT 143.195 -295.530 143.425 -294.260 ;
        RECT 144.175 -295.530 144.405 -294.250 ;
        RECT 146.110 -294.445 146.905 -294.155 ;
        RECT 147.080 -296.175 147.310 -294.675 ;
        RECT 148.060 -296.175 148.290 -291.990 ;
        RECT 148.550 -293.490 148.780 -291.810 ;
        RECT 153.205 -293.785 153.770 -288.630 ;
        RECT 157.420 -289.155 157.815 -285.990 ;
        RECT 158.830 -287.235 159.060 -285.735 ;
        RECT 159.320 -287.235 159.550 -285.735 ;
        RECT 161.180 -287.235 161.410 -284.735 ;
        RECT 161.670 -287.235 161.900 -284.735 ;
        RECT 162.295 -287.235 162.525 -284.735 ;
        RECT 162.785 -287.235 163.015 -284.735 ;
        RECT 163.435 -287.235 163.665 -284.735 ;
        RECT 163.925 -287.235 164.155 -284.735 ;
        RECT 164.415 -287.235 164.645 -284.735 ;
        RECT 164.980 -284.765 173.090 -284.455 ;
        RECT 164.980 -284.810 165.310 -284.765 ;
        RECT 165.065 -287.235 165.295 -285.735 ;
        RECT 165.555 -287.235 165.785 -285.735 ;
        RECT 154.920 -289.550 157.815 -289.155 ;
        RECT 154.920 -291.325 155.315 -289.550 ;
        RECT 154.790 -291.810 155.370 -291.325 ;
        RECT 164.925 -291.965 167.120 -291.730 ;
        RECT 157.935 -292.045 158.420 -292.015 ;
        RECT 157.935 -292.315 163.480 -292.045 ;
        RECT 164.925 -292.150 165.160 -291.965 ;
        RECT 157.935 -292.345 158.420 -292.315 ;
        RECT 152.060 -294.350 155.600 -293.785 ;
        RECT 150.125 -295.025 150.355 -294.525 ;
        RECT 150.615 -295.170 150.845 -294.525 ;
        RECT 151.105 -295.025 151.335 -294.525 ;
        RECT 151.595 -295.170 151.825 -294.525 ;
        RECT 150.125 -295.400 153.310 -295.170 ;
        RECT 150.125 -296.180 150.355 -295.400 ;
        RECT 150.615 -295.410 151.825 -295.400 ;
        RECT 151.105 -296.180 151.335 -295.410 ;
        RECT 152.085 -296.180 152.315 -295.400 ;
        RECT 142.085 -300.675 142.315 -299.175 ;
        RECT 140.320 -301.650 141.305 -301.380 ;
        RECT 141.595 -303.355 141.825 -301.860 ;
        RECT 141.590 -303.540 141.825 -303.355 ;
        RECT 142.085 -303.360 142.315 -301.860 ;
        RECT 142.575 -303.540 142.805 -301.860 ;
        RECT 143.065 -303.360 143.295 -299.175 ;
        RECT 145.130 -299.950 145.360 -299.170 ;
        RECT 146.110 -299.940 146.340 -299.170 ;
        RECT 145.620 -299.950 146.830 -299.940 ;
        RECT 147.090 -299.950 147.320 -299.170 ;
        RECT 145.130 -300.180 148.315 -299.950 ;
        RECT 145.130 -300.825 145.360 -300.325 ;
        RECT 145.620 -300.825 145.850 -300.180 ;
        RECT 146.110 -300.825 146.340 -300.325 ;
        RECT 146.600 -300.825 146.830 -300.180 ;
        RECT 149.320 -301.730 149.550 -298.730 ;
        RECT 150.375 -301.730 150.605 -298.730 ;
        RECT 150.865 -301.730 151.095 -298.730 ;
        RECT 151.355 -301.730 151.585 -298.730 ;
        RECT 152.415 -301.730 152.645 -298.730 ;
        RECT 143.555 -303.540 143.785 -301.860 ;
        RECT 153.570 -302.385 154.095 -302.025 ;
        RECT 153.600 -302.800 153.925 -302.385 ;
        RECT 148.825 -303.125 153.925 -302.800 ;
        RECT 141.590 -303.775 143.785 -303.540 ;
        RECT 149.320 -304.790 149.550 -303.290 ;
        RECT 149.810 -304.790 150.040 -303.290 ;
        RECT 150.300 -304.790 150.530 -303.290 ;
        RECT 151.510 -304.790 151.740 -303.290 ;
        RECT 152.000 -304.790 152.230 -303.290 ;
        RECT 155.035 -305.330 155.600 -294.350 ;
        RECT 159.125 -294.515 159.775 -293.765 ;
        RECT 160.555 -294.035 160.785 -293.035 ;
        RECT 161.045 -294.175 161.275 -293.035 ;
        RECT 161.535 -294.035 161.765 -293.035 ;
        RECT 162.025 -294.175 162.255 -293.035 ;
        RECT 163.210 -293.765 163.480 -292.315 ;
        RECT 164.930 -293.645 165.160 -292.150 ;
        RECT 165.420 -293.645 165.650 -292.145 ;
        RECT 165.910 -293.645 166.140 -291.965 ;
        RECT 163.210 -294.035 164.850 -293.765 ;
        RECT 160.555 -294.405 163.740 -294.175 ;
        RECT 164.580 -294.310 164.850 -294.035 ;
        RECT 159.375 -301.535 159.645 -294.515 ;
        RECT 160.555 -295.685 160.785 -294.405 ;
        RECT 161.045 -294.415 162.255 -294.405 ;
        RECT 161.535 -295.685 161.765 -294.415 ;
        RECT 162.515 -295.685 162.745 -294.405 ;
        RECT 164.450 -294.600 165.245 -294.310 ;
        RECT 165.420 -296.330 165.650 -294.830 ;
        RECT 166.400 -296.330 166.630 -292.145 ;
        RECT 166.890 -293.645 167.120 -291.965 ;
        RECT 170.400 -294.505 173.940 -293.940 ;
        RECT 168.465 -295.180 168.695 -294.680 ;
        RECT 168.955 -295.325 169.185 -294.680 ;
        RECT 169.445 -295.180 169.675 -294.680 ;
        RECT 169.935 -295.325 170.165 -294.680 ;
        RECT 168.465 -295.555 171.650 -295.325 ;
        RECT 168.465 -296.335 168.695 -295.555 ;
        RECT 168.955 -295.565 170.165 -295.555 ;
        RECT 169.445 -296.335 169.675 -295.565 ;
        RECT 170.425 -296.335 170.655 -295.555 ;
        RECT 160.425 -300.830 160.655 -299.330 ;
        RECT 158.660 -301.805 159.645 -301.535 ;
        RECT 159.935 -303.510 160.165 -302.015 ;
        RECT 159.930 -303.695 160.165 -303.510 ;
        RECT 160.425 -303.515 160.655 -302.015 ;
        RECT 160.915 -303.695 161.145 -302.015 ;
        RECT 161.405 -303.515 161.635 -299.330 ;
        RECT 163.470 -300.105 163.700 -299.325 ;
        RECT 164.450 -300.095 164.680 -299.325 ;
        RECT 163.960 -300.105 165.170 -300.095 ;
        RECT 165.430 -300.105 165.660 -299.325 ;
        RECT 163.470 -300.335 166.655 -300.105 ;
        RECT 163.470 -300.980 163.700 -300.480 ;
        RECT 163.960 -300.980 164.190 -300.335 ;
        RECT 164.450 -300.980 164.680 -300.480 ;
        RECT 164.940 -300.980 165.170 -300.335 ;
        RECT 167.660 -301.885 167.890 -298.885 ;
        RECT 168.715 -301.885 168.945 -298.885 ;
        RECT 169.205 -301.885 169.435 -298.885 ;
        RECT 169.695 -301.885 169.925 -298.885 ;
        RECT 170.755 -301.885 170.985 -298.885 ;
        RECT 161.895 -303.695 162.125 -302.015 ;
        RECT 171.910 -302.540 172.435 -302.180 ;
        RECT 171.940 -302.955 172.265 -302.540 ;
        RECT 167.165 -303.280 172.265 -302.955 ;
        RECT 159.930 -303.930 162.125 -303.695 ;
        RECT 167.660 -304.945 167.890 -303.445 ;
        RECT 168.150 -304.945 168.380 -303.445 ;
        RECT 168.640 -304.945 168.870 -303.445 ;
        RECT 169.850 -304.945 170.080 -303.445 ;
        RECT 170.340 -304.945 170.570 -303.445 ;
        RECT 152.215 -305.485 155.600 -305.330 ;
        RECT 173.375 -305.485 173.940 -294.505 ;
        RECT 174.360 -302.610 175.605 -275.165 ;
        RECT 176.415 -291.530 177.370 -272.960 ;
        RECT 179.795 -274.680 181.580 -274.000 ;
        RECT 188.825 -274.600 191.020 -274.365 ;
        RECT 179.795 -274.950 187.380 -274.680 ;
        RECT 188.825 -274.785 189.060 -274.600 ;
        RECT 179.795 -275.335 181.580 -274.950 ;
        RECT 183.025 -277.150 183.675 -276.400 ;
        RECT 184.455 -276.670 184.685 -275.670 ;
        RECT 184.945 -276.810 185.175 -275.670 ;
        RECT 185.435 -276.670 185.665 -275.670 ;
        RECT 185.925 -276.810 186.155 -275.670 ;
        RECT 187.110 -276.400 187.380 -274.950 ;
        RECT 188.830 -276.280 189.060 -274.785 ;
        RECT 189.320 -276.280 189.550 -274.780 ;
        RECT 189.810 -276.280 190.040 -274.600 ;
        RECT 187.110 -276.670 188.750 -276.400 ;
        RECT 184.455 -277.040 187.640 -276.810 ;
        RECT 188.480 -276.945 188.750 -276.670 ;
        RECT 183.275 -284.170 183.545 -277.150 ;
        RECT 184.455 -278.320 184.685 -277.040 ;
        RECT 184.945 -277.050 186.155 -277.040 ;
        RECT 185.435 -278.320 185.665 -277.050 ;
        RECT 186.415 -278.320 186.645 -277.040 ;
        RECT 188.350 -277.235 189.145 -276.945 ;
        RECT 189.320 -278.965 189.550 -277.465 ;
        RECT 190.300 -278.965 190.530 -274.780 ;
        RECT 190.790 -276.280 191.020 -274.600 ;
        RECT 194.300 -277.140 197.840 -276.575 ;
        RECT 192.365 -277.815 192.595 -277.315 ;
        RECT 192.855 -277.960 193.085 -277.315 ;
        RECT 193.345 -277.815 193.575 -277.315 ;
        RECT 193.835 -277.960 194.065 -277.315 ;
        RECT 192.365 -278.190 195.550 -277.960 ;
        RECT 192.365 -278.970 192.595 -278.190 ;
        RECT 192.855 -278.200 194.065 -278.190 ;
        RECT 193.345 -278.970 193.575 -278.200 ;
        RECT 194.325 -278.970 194.555 -278.190 ;
        RECT 184.325 -283.465 184.555 -281.965 ;
        RECT 182.560 -284.440 183.545 -284.170 ;
        RECT 183.835 -286.145 184.065 -284.650 ;
        RECT 183.830 -286.330 184.065 -286.145 ;
        RECT 184.325 -286.150 184.555 -284.650 ;
        RECT 184.815 -286.330 185.045 -284.650 ;
        RECT 185.305 -286.150 185.535 -281.965 ;
        RECT 187.370 -282.740 187.600 -281.960 ;
        RECT 188.350 -282.730 188.580 -281.960 ;
        RECT 187.860 -282.740 189.070 -282.730 ;
        RECT 189.330 -282.740 189.560 -281.960 ;
        RECT 187.370 -282.970 190.555 -282.740 ;
        RECT 187.370 -283.615 187.600 -283.115 ;
        RECT 187.860 -283.615 188.090 -282.970 ;
        RECT 188.350 -283.615 188.580 -283.115 ;
        RECT 188.840 -283.615 189.070 -282.970 ;
        RECT 191.560 -284.520 191.790 -281.520 ;
        RECT 192.615 -284.520 192.845 -281.520 ;
        RECT 193.105 -284.520 193.335 -281.520 ;
        RECT 193.595 -284.520 193.825 -281.520 ;
        RECT 194.655 -284.520 194.885 -281.520 ;
        RECT 185.795 -286.330 186.025 -284.650 ;
        RECT 195.810 -285.175 196.335 -284.815 ;
        RECT 195.840 -285.590 196.165 -285.175 ;
        RECT 191.065 -285.915 196.165 -285.590 ;
        RECT 183.830 -286.565 186.025 -286.330 ;
        RECT 191.560 -287.580 191.790 -286.080 ;
        RECT 192.050 -287.580 192.280 -286.080 ;
        RECT 192.540 -287.580 192.770 -286.080 ;
        RECT 193.750 -287.580 193.980 -286.080 ;
        RECT 194.240 -287.580 194.470 -286.080 ;
        RECT 195.405 -288.120 195.970 -288.115 ;
        RECT 197.275 -288.120 197.840 -277.140 ;
        RECT 201.520 -283.310 201.750 -280.810 ;
        RECT 202.865 -283.310 203.095 -280.810 ;
        RECT 203.355 -283.310 203.585 -280.810 ;
        RECT 203.845 -283.310 204.075 -280.810 ;
        RECT 204.495 -283.310 204.725 -280.810 ;
        RECT 206.125 -283.310 206.355 -280.810 ;
        RECT 207.265 -282.310 207.495 -280.810 ;
        RECT 200.365 -284.110 201.055 -284.090 ;
        RECT 204.395 -284.110 205.085 -284.090 ;
        RECT 206.320 -284.110 206.590 -283.745 ;
        RECT 200.365 -284.330 206.590 -284.110 ;
        RECT 200.365 -284.360 201.055 -284.330 ;
        RECT 204.395 -284.360 205.085 -284.330 ;
        RECT 206.320 -284.435 206.590 -284.330 ;
        RECT 207.180 -284.510 207.510 -284.450 ;
        RECT 210.745 -284.510 211.825 -272.960 ;
        RECT 199.560 -286.045 200.075 -285.590 ;
        RECT 194.455 -288.685 197.840 -288.120 ;
        RECT 176.415 -291.945 180.665 -291.530 ;
        RECT 188.785 -291.865 190.980 -291.630 ;
        RECT 176.415 -292.215 187.340 -291.945 ;
        RECT 188.785 -292.050 189.020 -291.865 ;
        RECT 176.415 -292.485 180.665 -292.215 ;
        RECT 182.985 -294.415 183.635 -293.665 ;
        RECT 184.415 -293.935 184.645 -292.935 ;
        RECT 184.905 -294.075 185.135 -292.935 ;
        RECT 185.395 -293.935 185.625 -292.935 ;
        RECT 185.885 -294.075 186.115 -292.935 ;
        RECT 187.070 -293.665 187.340 -292.215 ;
        RECT 188.790 -293.545 189.020 -292.050 ;
        RECT 189.280 -293.545 189.510 -292.045 ;
        RECT 189.770 -293.545 190.000 -291.865 ;
        RECT 187.070 -293.935 188.710 -293.665 ;
        RECT 184.415 -294.305 187.600 -294.075 ;
        RECT 188.440 -294.210 188.710 -293.935 ;
        RECT 183.235 -301.435 183.505 -294.415 ;
        RECT 184.415 -295.585 184.645 -294.305 ;
        RECT 184.905 -294.315 186.115 -294.305 ;
        RECT 185.395 -295.585 185.625 -294.315 ;
        RECT 186.375 -295.585 186.605 -294.305 ;
        RECT 188.310 -294.500 189.105 -294.210 ;
        RECT 189.280 -296.230 189.510 -294.730 ;
        RECT 190.260 -296.230 190.490 -292.045 ;
        RECT 190.750 -293.545 190.980 -291.865 ;
        RECT 195.405 -293.840 195.970 -288.685 ;
        RECT 199.620 -289.210 200.015 -286.045 ;
        RECT 201.030 -287.290 201.260 -285.790 ;
        RECT 201.520 -287.290 201.750 -285.790 ;
        RECT 203.380 -287.290 203.610 -284.790 ;
        RECT 203.870 -287.290 204.100 -284.790 ;
        RECT 204.495 -287.290 204.725 -284.790 ;
        RECT 204.985 -287.290 205.215 -284.790 ;
        RECT 205.635 -287.290 205.865 -284.790 ;
        RECT 206.125 -287.290 206.355 -284.790 ;
        RECT 206.615 -287.290 206.845 -284.790 ;
        RECT 207.180 -284.820 215.290 -284.510 ;
        RECT 207.180 -284.865 207.510 -284.820 ;
        RECT 207.265 -287.290 207.495 -285.790 ;
        RECT 207.755 -287.290 207.985 -285.790 ;
        RECT 197.120 -289.605 200.015 -289.210 ;
        RECT 197.120 -291.380 197.515 -289.605 ;
        RECT 196.990 -291.865 197.570 -291.380 ;
        RECT 207.125 -292.020 209.320 -291.785 ;
        RECT 200.135 -292.100 200.620 -292.070 ;
        RECT 200.135 -292.370 205.680 -292.100 ;
        RECT 207.125 -292.205 207.360 -292.020 ;
        RECT 200.135 -292.400 200.620 -292.370 ;
        RECT 194.260 -294.405 197.800 -293.840 ;
        RECT 192.325 -295.080 192.555 -294.580 ;
        RECT 192.815 -295.225 193.045 -294.580 ;
        RECT 193.305 -295.080 193.535 -294.580 ;
        RECT 193.795 -295.225 194.025 -294.580 ;
        RECT 192.325 -295.455 195.510 -295.225 ;
        RECT 192.325 -296.235 192.555 -295.455 ;
        RECT 192.815 -295.465 194.025 -295.455 ;
        RECT 193.305 -296.235 193.535 -295.465 ;
        RECT 194.285 -296.235 194.515 -295.455 ;
        RECT 184.285 -300.730 184.515 -299.230 ;
        RECT 182.520 -301.705 183.505 -301.435 ;
        RECT 174.440 -303.455 175.555 -302.610 ;
        RECT 183.795 -303.410 184.025 -301.915 ;
        RECT 183.790 -303.595 184.025 -303.410 ;
        RECT 184.285 -303.415 184.515 -301.915 ;
        RECT 184.775 -303.595 185.005 -301.915 ;
        RECT 185.265 -303.415 185.495 -299.230 ;
        RECT 187.330 -300.005 187.560 -299.225 ;
        RECT 188.310 -299.995 188.540 -299.225 ;
        RECT 187.820 -300.005 189.030 -299.995 ;
        RECT 189.290 -300.005 189.520 -299.225 ;
        RECT 187.330 -300.235 190.515 -300.005 ;
        RECT 187.330 -300.880 187.560 -300.380 ;
        RECT 187.820 -300.880 188.050 -300.235 ;
        RECT 188.310 -300.880 188.540 -300.380 ;
        RECT 188.800 -300.880 189.030 -300.235 ;
        RECT 191.520 -301.785 191.750 -298.785 ;
        RECT 192.575 -301.785 192.805 -298.785 ;
        RECT 193.065 -301.785 193.295 -298.785 ;
        RECT 193.555 -301.785 193.785 -298.785 ;
        RECT 194.615 -301.785 194.845 -298.785 ;
        RECT 185.755 -303.595 185.985 -301.915 ;
        RECT 195.770 -302.440 196.295 -302.080 ;
        RECT 195.800 -302.855 196.125 -302.440 ;
        RECT 191.025 -303.180 196.125 -302.855 ;
        RECT 183.790 -303.830 185.985 -303.595 ;
        RECT 191.520 -304.845 191.750 -303.345 ;
        RECT 192.010 -304.845 192.240 -303.345 ;
        RECT 192.500 -304.845 192.730 -303.345 ;
        RECT 193.710 -304.845 193.940 -303.345 ;
        RECT 194.200 -304.845 194.430 -303.345 ;
        RECT 197.235 -305.385 197.800 -294.405 ;
        RECT 201.325 -294.570 201.975 -293.820 ;
        RECT 202.755 -294.090 202.985 -293.090 ;
        RECT 203.245 -294.230 203.475 -293.090 ;
        RECT 203.735 -294.090 203.965 -293.090 ;
        RECT 204.225 -294.230 204.455 -293.090 ;
        RECT 205.410 -293.820 205.680 -292.370 ;
        RECT 207.130 -293.700 207.360 -292.205 ;
        RECT 207.620 -293.700 207.850 -292.200 ;
        RECT 208.110 -293.700 208.340 -292.020 ;
        RECT 205.410 -294.090 207.050 -293.820 ;
        RECT 202.755 -294.460 205.940 -294.230 ;
        RECT 206.780 -294.365 207.050 -294.090 ;
        RECT 201.575 -301.590 201.845 -294.570 ;
        RECT 202.755 -295.740 202.985 -294.460 ;
        RECT 203.245 -294.470 204.455 -294.460 ;
        RECT 203.735 -295.740 203.965 -294.470 ;
        RECT 204.715 -295.740 204.945 -294.460 ;
        RECT 206.650 -294.655 207.445 -294.365 ;
        RECT 207.620 -296.385 207.850 -294.885 ;
        RECT 208.600 -296.385 208.830 -292.200 ;
        RECT 209.090 -293.700 209.320 -292.020 ;
        RECT 212.600 -294.560 216.140 -293.995 ;
        RECT 210.665 -295.235 210.895 -294.735 ;
        RECT 211.155 -295.380 211.385 -294.735 ;
        RECT 211.645 -295.235 211.875 -294.735 ;
        RECT 212.135 -295.380 212.365 -294.735 ;
        RECT 210.665 -295.610 213.850 -295.380 ;
        RECT 210.665 -296.390 210.895 -295.610 ;
        RECT 211.155 -295.620 212.365 -295.610 ;
        RECT 211.645 -296.390 211.875 -295.620 ;
        RECT 212.625 -296.390 212.855 -295.610 ;
        RECT 202.625 -300.885 202.855 -299.385 ;
        RECT 200.860 -301.860 201.845 -301.590 ;
        RECT 202.135 -303.565 202.365 -302.070 ;
        RECT 202.130 -303.750 202.365 -303.565 ;
        RECT 202.625 -303.570 202.855 -302.070 ;
        RECT 203.115 -303.750 203.345 -302.070 ;
        RECT 203.605 -303.570 203.835 -299.385 ;
        RECT 205.670 -300.160 205.900 -299.380 ;
        RECT 206.650 -300.150 206.880 -299.380 ;
        RECT 206.160 -300.160 207.370 -300.150 ;
        RECT 207.630 -300.160 207.860 -299.380 ;
        RECT 205.670 -300.390 208.855 -300.160 ;
        RECT 205.670 -301.035 205.900 -300.535 ;
        RECT 206.160 -301.035 206.390 -300.390 ;
        RECT 206.650 -301.035 206.880 -300.535 ;
        RECT 207.140 -301.035 207.370 -300.390 ;
        RECT 209.860 -301.940 210.090 -298.940 ;
        RECT 210.915 -301.940 211.145 -298.940 ;
        RECT 211.405 -301.940 211.635 -298.940 ;
        RECT 211.895 -301.940 212.125 -298.940 ;
        RECT 212.955 -301.940 213.185 -298.940 ;
        RECT 204.095 -303.750 204.325 -302.070 ;
        RECT 214.110 -302.595 214.635 -302.235 ;
        RECT 214.140 -303.010 214.465 -302.595 ;
        RECT 209.365 -303.335 214.465 -303.010 ;
        RECT 202.130 -303.985 204.325 -303.750 ;
        RECT 209.860 -305.000 210.090 -303.500 ;
        RECT 210.350 -305.000 210.580 -303.500 ;
        RECT 210.840 -305.000 211.070 -303.500 ;
        RECT 212.050 -305.000 212.280 -303.500 ;
        RECT 212.540 -305.000 212.770 -303.500 ;
        RECT 152.215 -305.895 173.940 -305.485 ;
        RECT 152.235 -306.050 173.940 -305.895 ;
        RECT 194.415 -305.540 197.800 -305.385 ;
        RECT 215.575 -305.540 216.140 -294.560 ;
        RECT 216.685 -302.295 218.010 -265.630 ;
        RECT 218.895 -272.925 258.700 -271.915 ;
        RECT 218.895 -291.875 219.905 -272.925 ;
        RECT 224.315 -274.875 225.800 -274.445 ;
        RECT 233.140 -274.795 235.335 -274.560 ;
        RECT 224.315 -275.145 231.695 -274.875 ;
        RECT 233.140 -274.980 233.375 -274.795 ;
        RECT 224.315 -275.555 225.800 -275.145 ;
        RECT 227.340 -277.345 227.990 -276.595 ;
        RECT 228.770 -276.865 229.000 -275.865 ;
        RECT 229.260 -277.005 229.490 -275.865 ;
        RECT 229.750 -276.865 229.980 -275.865 ;
        RECT 230.240 -277.005 230.470 -275.865 ;
        RECT 231.425 -276.595 231.695 -275.145 ;
        RECT 233.145 -276.475 233.375 -274.980 ;
        RECT 233.635 -276.475 233.865 -274.975 ;
        RECT 234.125 -276.475 234.355 -274.795 ;
        RECT 231.425 -276.865 233.065 -276.595 ;
        RECT 228.770 -277.235 231.955 -277.005 ;
        RECT 232.795 -277.140 233.065 -276.865 ;
        RECT 227.590 -284.365 227.860 -277.345 ;
        RECT 228.770 -278.515 229.000 -277.235 ;
        RECT 229.260 -277.245 230.470 -277.235 ;
        RECT 229.750 -278.515 229.980 -277.245 ;
        RECT 230.730 -278.515 230.960 -277.235 ;
        RECT 232.665 -277.430 233.460 -277.140 ;
        RECT 233.635 -279.160 233.865 -277.660 ;
        RECT 234.615 -279.160 234.845 -274.975 ;
        RECT 235.105 -276.475 235.335 -274.795 ;
        RECT 238.615 -277.335 242.155 -276.770 ;
        RECT 236.680 -278.010 236.910 -277.510 ;
        RECT 237.170 -278.155 237.400 -277.510 ;
        RECT 237.660 -278.010 237.890 -277.510 ;
        RECT 238.150 -278.155 238.380 -277.510 ;
        RECT 236.680 -278.385 239.865 -278.155 ;
        RECT 236.680 -279.165 236.910 -278.385 ;
        RECT 237.170 -278.395 238.380 -278.385 ;
        RECT 237.660 -279.165 237.890 -278.395 ;
        RECT 238.640 -279.165 238.870 -278.385 ;
        RECT 228.640 -283.660 228.870 -282.160 ;
        RECT 226.875 -284.635 227.860 -284.365 ;
        RECT 228.150 -286.340 228.380 -284.845 ;
        RECT 228.145 -286.525 228.380 -286.340 ;
        RECT 228.640 -286.345 228.870 -284.845 ;
        RECT 229.130 -286.525 229.360 -284.845 ;
        RECT 229.620 -286.345 229.850 -282.160 ;
        RECT 231.685 -282.935 231.915 -282.155 ;
        RECT 232.665 -282.925 232.895 -282.155 ;
        RECT 232.175 -282.935 233.385 -282.925 ;
        RECT 233.645 -282.935 233.875 -282.155 ;
        RECT 231.685 -283.165 234.870 -282.935 ;
        RECT 231.685 -283.810 231.915 -283.310 ;
        RECT 232.175 -283.810 232.405 -283.165 ;
        RECT 232.665 -283.810 232.895 -283.310 ;
        RECT 233.155 -283.810 233.385 -283.165 ;
        RECT 235.875 -284.715 236.105 -281.715 ;
        RECT 236.930 -284.715 237.160 -281.715 ;
        RECT 237.420 -284.715 237.650 -281.715 ;
        RECT 237.910 -284.715 238.140 -281.715 ;
        RECT 238.970 -284.715 239.200 -281.715 ;
        RECT 230.110 -286.525 230.340 -284.845 ;
        RECT 240.125 -285.370 240.650 -285.010 ;
        RECT 240.155 -285.785 240.480 -285.370 ;
        RECT 235.380 -286.110 240.480 -285.785 ;
        RECT 228.145 -286.760 230.340 -286.525 ;
        RECT 235.875 -287.775 236.105 -286.275 ;
        RECT 236.365 -287.775 236.595 -286.275 ;
        RECT 236.855 -287.775 237.085 -286.275 ;
        RECT 238.065 -287.775 238.295 -286.275 ;
        RECT 238.555 -287.775 238.785 -286.275 ;
        RECT 239.720 -288.315 240.285 -288.310 ;
        RECT 241.590 -288.315 242.155 -277.335 ;
        RECT 245.835 -283.505 246.065 -281.005 ;
        RECT 247.180 -283.505 247.410 -281.005 ;
        RECT 247.670 -283.505 247.900 -281.005 ;
        RECT 248.160 -283.505 248.390 -281.005 ;
        RECT 248.810 -283.505 249.040 -281.005 ;
        RECT 250.440 -283.505 250.670 -281.005 ;
        RECT 251.580 -282.505 251.810 -281.005 ;
        RECT 244.680 -284.305 245.370 -284.285 ;
        RECT 248.710 -284.305 249.400 -284.285 ;
        RECT 250.635 -284.305 250.905 -283.940 ;
        RECT 244.680 -284.525 250.905 -284.305 ;
        RECT 244.680 -284.555 245.370 -284.525 ;
        RECT 248.710 -284.555 249.400 -284.525 ;
        RECT 250.635 -284.630 250.905 -284.525 ;
        RECT 251.495 -284.705 251.825 -284.645 ;
        RECT 257.690 -284.705 258.700 -272.925 ;
        RECT 243.875 -286.240 244.390 -285.785 ;
        RECT 238.770 -288.880 242.155 -288.315 ;
        RECT 218.895 -292.140 225.545 -291.875 ;
        RECT 233.100 -292.060 235.295 -291.825 ;
        RECT 218.895 -292.410 231.655 -292.140 ;
        RECT 233.100 -292.245 233.335 -292.060 ;
        RECT 218.895 -292.885 225.545 -292.410 ;
        RECT 227.300 -294.610 227.950 -293.860 ;
        RECT 228.730 -294.130 228.960 -293.130 ;
        RECT 229.220 -294.270 229.450 -293.130 ;
        RECT 229.710 -294.130 229.940 -293.130 ;
        RECT 230.200 -294.270 230.430 -293.130 ;
        RECT 231.385 -293.860 231.655 -292.410 ;
        RECT 233.105 -293.740 233.335 -292.245 ;
        RECT 233.595 -293.740 233.825 -292.240 ;
        RECT 234.085 -293.740 234.315 -292.060 ;
        RECT 231.385 -294.130 233.025 -293.860 ;
        RECT 228.730 -294.500 231.915 -294.270 ;
        RECT 232.755 -294.405 233.025 -294.130 ;
        RECT 227.550 -301.630 227.820 -294.610 ;
        RECT 228.730 -295.780 228.960 -294.500 ;
        RECT 229.220 -294.510 230.430 -294.500 ;
        RECT 229.710 -295.780 229.940 -294.510 ;
        RECT 230.690 -295.780 230.920 -294.500 ;
        RECT 232.625 -294.695 233.420 -294.405 ;
        RECT 233.595 -296.425 233.825 -294.925 ;
        RECT 234.575 -296.425 234.805 -292.240 ;
        RECT 235.065 -293.740 235.295 -292.060 ;
        RECT 239.720 -294.035 240.285 -288.880 ;
        RECT 243.935 -289.405 244.330 -286.240 ;
        RECT 245.345 -287.485 245.575 -285.985 ;
        RECT 245.835 -287.485 246.065 -285.985 ;
        RECT 247.695 -287.485 247.925 -284.985 ;
        RECT 248.185 -287.485 248.415 -284.985 ;
        RECT 248.810 -287.485 249.040 -284.985 ;
        RECT 249.300 -287.485 249.530 -284.985 ;
        RECT 249.950 -287.485 250.180 -284.985 ;
        RECT 250.440 -287.485 250.670 -284.985 ;
        RECT 250.930 -287.485 251.160 -284.985 ;
        RECT 251.495 -285.015 259.605 -284.705 ;
        RECT 251.495 -285.060 251.825 -285.015 ;
        RECT 251.580 -287.485 251.810 -285.985 ;
        RECT 252.070 -287.485 252.300 -285.985 ;
        RECT 241.435 -289.800 244.330 -289.405 ;
        RECT 241.435 -291.575 241.830 -289.800 ;
        RECT 241.305 -292.060 241.885 -291.575 ;
        RECT 251.440 -292.215 253.635 -291.980 ;
        RECT 244.450 -292.295 244.935 -292.265 ;
        RECT 244.450 -292.565 249.995 -292.295 ;
        RECT 251.440 -292.400 251.675 -292.215 ;
        RECT 244.450 -292.595 244.935 -292.565 ;
        RECT 238.575 -294.600 242.115 -294.035 ;
        RECT 236.640 -295.275 236.870 -294.775 ;
        RECT 237.130 -295.420 237.360 -294.775 ;
        RECT 237.620 -295.275 237.850 -294.775 ;
        RECT 238.110 -295.420 238.340 -294.775 ;
        RECT 236.640 -295.650 239.825 -295.420 ;
        RECT 236.640 -296.430 236.870 -295.650 ;
        RECT 237.130 -295.660 238.340 -295.650 ;
        RECT 237.620 -296.430 237.850 -295.660 ;
        RECT 238.600 -296.430 238.830 -295.650 ;
        RECT 228.600 -300.925 228.830 -299.425 ;
        RECT 226.835 -301.900 227.820 -301.630 ;
        RECT 216.685 -303.950 218.370 -302.295 ;
        RECT 228.110 -303.605 228.340 -302.110 ;
        RECT 228.105 -303.790 228.340 -303.605 ;
        RECT 228.600 -303.610 228.830 -302.110 ;
        RECT 229.090 -303.790 229.320 -302.110 ;
        RECT 229.580 -303.610 229.810 -299.425 ;
        RECT 231.645 -300.200 231.875 -299.420 ;
        RECT 232.625 -300.190 232.855 -299.420 ;
        RECT 232.135 -300.200 233.345 -300.190 ;
        RECT 233.605 -300.200 233.835 -299.420 ;
        RECT 231.645 -300.430 234.830 -300.200 ;
        RECT 231.645 -301.075 231.875 -300.575 ;
        RECT 232.135 -301.075 232.365 -300.430 ;
        RECT 232.625 -301.075 232.855 -300.575 ;
        RECT 233.115 -301.075 233.345 -300.430 ;
        RECT 235.835 -301.980 236.065 -298.980 ;
        RECT 236.890 -301.980 237.120 -298.980 ;
        RECT 237.380 -301.980 237.610 -298.980 ;
        RECT 237.870 -301.980 238.100 -298.980 ;
        RECT 238.930 -301.980 239.160 -298.980 ;
        RECT 230.070 -303.790 230.300 -302.110 ;
        RECT 240.085 -302.635 240.610 -302.275 ;
        RECT 240.115 -303.050 240.440 -302.635 ;
        RECT 235.340 -303.375 240.440 -303.050 ;
        RECT 228.105 -304.025 230.300 -303.790 ;
        RECT 235.835 -305.040 236.065 -303.540 ;
        RECT 236.325 -305.040 236.555 -303.540 ;
        RECT 236.815 -305.040 237.045 -303.540 ;
        RECT 238.025 -305.040 238.255 -303.540 ;
        RECT 238.515 -305.040 238.745 -303.540 ;
        RECT 194.415 -305.950 216.140 -305.540 ;
        RECT 241.550 -305.580 242.115 -294.600 ;
        RECT 245.640 -294.765 246.290 -294.015 ;
        RECT 247.070 -294.285 247.300 -293.285 ;
        RECT 247.560 -294.425 247.790 -293.285 ;
        RECT 248.050 -294.285 248.280 -293.285 ;
        RECT 248.540 -294.425 248.770 -293.285 ;
        RECT 249.725 -294.015 249.995 -292.565 ;
        RECT 251.445 -293.895 251.675 -292.400 ;
        RECT 251.935 -293.895 252.165 -292.395 ;
        RECT 252.425 -293.895 252.655 -292.215 ;
        RECT 249.725 -294.285 251.365 -294.015 ;
        RECT 247.070 -294.655 250.255 -294.425 ;
        RECT 251.095 -294.560 251.365 -294.285 ;
        RECT 245.890 -301.785 246.160 -294.765 ;
        RECT 247.070 -295.935 247.300 -294.655 ;
        RECT 247.560 -294.665 248.770 -294.655 ;
        RECT 248.050 -295.935 248.280 -294.665 ;
        RECT 249.030 -295.935 249.260 -294.655 ;
        RECT 250.965 -294.850 251.760 -294.560 ;
        RECT 251.935 -296.580 252.165 -295.080 ;
        RECT 252.915 -296.580 253.145 -292.395 ;
        RECT 253.405 -293.895 253.635 -292.215 ;
        RECT 256.915 -294.755 260.455 -294.190 ;
        RECT 254.980 -295.430 255.210 -294.930 ;
        RECT 255.470 -295.575 255.700 -294.930 ;
        RECT 255.960 -295.430 256.190 -294.930 ;
        RECT 256.450 -295.575 256.680 -294.930 ;
        RECT 254.980 -295.805 258.165 -295.575 ;
        RECT 254.980 -296.585 255.210 -295.805 ;
        RECT 255.470 -295.815 256.680 -295.805 ;
        RECT 255.960 -296.585 256.190 -295.815 ;
        RECT 256.940 -296.585 257.170 -295.805 ;
        RECT 246.940 -301.080 247.170 -299.580 ;
        RECT 245.175 -302.055 246.160 -301.785 ;
        RECT 246.450 -303.760 246.680 -302.265 ;
        RECT 246.445 -303.945 246.680 -303.760 ;
        RECT 246.940 -303.765 247.170 -302.265 ;
        RECT 247.430 -303.945 247.660 -302.265 ;
        RECT 247.920 -303.765 248.150 -299.580 ;
        RECT 249.985 -300.355 250.215 -299.575 ;
        RECT 250.965 -300.345 251.195 -299.575 ;
        RECT 250.475 -300.355 251.685 -300.345 ;
        RECT 251.945 -300.355 252.175 -299.575 ;
        RECT 249.985 -300.585 253.170 -300.355 ;
        RECT 249.985 -301.230 250.215 -300.730 ;
        RECT 250.475 -301.230 250.705 -300.585 ;
        RECT 250.965 -301.230 251.195 -300.730 ;
        RECT 251.455 -301.230 251.685 -300.585 ;
        RECT 254.175 -302.135 254.405 -299.135 ;
        RECT 255.230 -302.135 255.460 -299.135 ;
        RECT 255.720 -302.135 255.950 -299.135 ;
        RECT 256.210 -302.135 256.440 -299.135 ;
        RECT 257.270 -302.135 257.500 -299.135 ;
        RECT 248.410 -303.945 248.640 -302.265 ;
        RECT 258.425 -302.790 258.950 -302.430 ;
        RECT 258.455 -303.205 258.780 -302.790 ;
        RECT 253.680 -303.530 258.780 -303.205 ;
        RECT 246.445 -304.180 248.640 -303.945 ;
        RECT 254.175 -305.195 254.405 -303.695 ;
        RECT 254.665 -305.195 254.895 -303.695 ;
        RECT 255.155 -305.195 255.385 -303.695 ;
        RECT 256.365 -305.195 256.595 -303.695 ;
        RECT 256.855 -305.195 257.085 -303.695 ;
        RECT 194.435 -306.105 216.140 -305.950 ;
        RECT 238.730 -305.735 242.115 -305.580 ;
        RECT 259.890 -305.735 260.455 -294.755 ;
        RECT 261.005 -301.600 262.135 -263.230 ;
        RECT 265.290 -273.250 305.220 -271.955 ;
        RECT 265.290 -291.270 266.585 -273.250 ;
        RECT 269.270 -274.705 270.500 -274.225 ;
        RECT 279.130 -274.625 281.325 -274.390 ;
        RECT 269.270 -274.975 277.685 -274.705 ;
        RECT 279.130 -274.810 279.365 -274.625 ;
        RECT 269.270 -275.325 270.500 -274.975 ;
        RECT 273.330 -277.175 273.980 -276.425 ;
        RECT 274.760 -276.695 274.990 -275.695 ;
        RECT 275.250 -276.835 275.480 -275.695 ;
        RECT 275.740 -276.695 275.970 -275.695 ;
        RECT 276.230 -276.835 276.460 -275.695 ;
        RECT 277.415 -276.425 277.685 -274.975 ;
        RECT 279.135 -276.305 279.365 -274.810 ;
        RECT 279.625 -276.305 279.855 -274.805 ;
        RECT 280.115 -276.305 280.345 -274.625 ;
        RECT 277.415 -276.695 279.055 -276.425 ;
        RECT 274.760 -277.065 277.945 -276.835 ;
        RECT 278.785 -276.970 279.055 -276.695 ;
        RECT 273.580 -284.195 273.850 -277.175 ;
        RECT 274.760 -278.345 274.990 -277.065 ;
        RECT 275.250 -277.075 276.460 -277.065 ;
        RECT 275.740 -278.345 275.970 -277.075 ;
        RECT 276.720 -278.345 276.950 -277.065 ;
        RECT 278.655 -277.260 279.450 -276.970 ;
        RECT 279.625 -278.990 279.855 -277.490 ;
        RECT 280.605 -278.990 280.835 -274.805 ;
        RECT 281.095 -276.305 281.325 -274.625 ;
        RECT 284.605 -277.165 288.145 -276.600 ;
        RECT 282.670 -277.840 282.900 -277.340 ;
        RECT 283.160 -277.985 283.390 -277.340 ;
        RECT 283.650 -277.840 283.880 -277.340 ;
        RECT 284.140 -277.985 284.370 -277.340 ;
        RECT 282.670 -278.215 285.855 -277.985 ;
        RECT 282.670 -278.995 282.900 -278.215 ;
        RECT 283.160 -278.225 284.370 -278.215 ;
        RECT 283.650 -278.995 283.880 -278.225 ;
        RECT 284.630 -278.995 284.860 -278.215 ;
        RECT 274.630 -283.490 274.860 -281.990 ;
        RECT 272.865 -284.465 273.850 -284.195 ;
        RECT 274.140 -286.170 274.370 -284.675 ;
        RECT 274.135 -286.355 274.370 -286.170 ;
        RECT 274.630 -286.175 274.860 -284.675 ;
        RECT 275.120 -286.355 275.350 -284.675 ;
        RECT 275.610 -286.175 275.840 -281.990 ;
        RECT 277.675 -282.765 277.905 -281.985 ;
        RECT 278.655 -282.755 278.885 -281.985 ;
        RECT 278.165 -282.765 279.375 -282.755 ;
        RECT 279.635 -282.765 279.865 -281.985 ;
        RECT 277.675 -282.995 280.860 -282.765 ;
        RECT 277.675 -283.640 277.905 -283.140 ;
        RECT 278.165 -283.640 278.395 -282.995 ;
        RECT 278.655 -283.640 278.885 -283.140 ;
        RECT 279.145 -283.640 279.375 -282.995 ;
        RECT 281.865 -284.545 282.095 -281.545 ;
        RECT 282.920 -284.545 283.150 -281.545 ;
        RECT 283.410 -284.545 283.640 -281.545 ;
        RECT 283.900 -284.545 284.130 -281.545 ;
        RECT 284.960 -284.545 285.190 -281.545 ;
        RECT 276.100 -286.355 276.330 -284.675 ;
        RECT 286.115 -285.200 286.640 -284.840 ;
        RECT 286.145 -285.615 286.470 -285.200 ;
        RECT 281.370 -285.940 286.470 -285.615 ;
        RECT 274.135 -286.590 276.330 -286.355 ;
        RECT 281.865 -287.605 282.095 -286.105 ;
        RECT 282.355 -287.605 282.585 -286.105 ;
        RECT 282.845 -287.605 283.075 -286.105 ;
        RECT 284.055 -287.605 284.285 -286.105 ;
        RECT 284.545 -287.605 284.775 -286.105 ;
        RECT 285.710 -288.145 286.275 -288.140 ;
        RECT 287.580 -288.145 288.145 -277.165 ;
        RECT 291.825 -283.335 292.055 -280.835 ;
        RECT 293.170 -283.335 293.400 -280.835 ;
        RECT 293.660 -283.335 293.890 -280.835 ;
        RECT 294.150 -283.335 294.380 -280.835 ;
        RECT 294.800 -283.335 295.030 -280.835 ;
        RECT 296.430 -283.335 296.660 -280.835 ;
        RECT 297.570 -282.335 297.800 -280.835 ;
        RECT 290.670 -284.135 291.360 -284.115 ;
        RECT 294.700 -284.135 295.390 -284.115 ;
        RECT 296.625 -284.135 296.895 -283.770 ;
        RECT 290.670 -284.355 296.895 -284.135 ;
        RECT 290.670 -284.385 291.360 -284.355 ;
        RECT 294.700 -284.385 295.390 -284.355 ;
        RECT 296.625 -284.460 296.895 -284.355 ;
        RECT 297.485 -284.535 297.815 -284.475 ;
        RECT 303.925 -284.535 305.220 -273.250 ;
        RECT 306.975 -273.535 308.080 -260.445 ;
        RECT 309.235 -273.350 349.155 -272.160 ;
        RECT 306.460 -275.105 308.340 -273.535 ;
        RECT 289.865 -286.070 290.380 -285.615 ;
        RECT 284.760 -288.710 288.145 -288.145 ;
        RECT 265.290 -291.970 271.330 -291.270 ;
        RECT 279.090 -291.890 281.285 -291.655 ;
        RECT 265.290 -292.240 277.645 -291.970 ;
        RECT 279.090 -292.075 279.325 -291.890 ;
        RECT 265.290 -292.565 271.330 -292.240 ;
        RECT 273.290 -294.440 273.940 -293.690 ;
        RECT 274.720 -293.960 274.950 -292.960 ;
        RECT 275.210 -294.100 275.440 -292.960 ;
        RECT 275.700 -293.960 275.930 -292.960 ;
        RECT 276.190 -294.100 276.420 -292.960 ;
        RECT 277.375 -293.690 277.645 -292.240 ;
        RECT 279.095 -293.570 279.325 -292.075 ;
        RECT 279.585 -293.570 279.815 -292.070 ;
        RECT 280.075 -293.570 280.305 -291.890 ;
        RECT 277.375 -293.960 279.015 -293.690 ;
        RECT 274.720 -294.330 277.905 -294.100 ;
        RECT 278.745 -294.235 279.015 -293.960 ;
        RECT 273.540 -301.460 273.810 -294.440 ;
        RECT 274.720 -295.610 274.950 -294.330 ;
        RECT 275.210 -294.340 276.420 -294.330 ;
        RECT 275.700 -295.610 275.930 -294.340 ;
        RECT 276.680 -295.610 276.910 -294.330 ;
        RECT 278.615 -294.525 279.410 -294.235 ;
        RECT 279.585 -296.255 279.815 -294.755 ;
        RECT 280.565 -296.255 280.795 -292.070 ;
        RECT 281.055 -293.570 281.285 -291.890 ;
        RECT 285.710 -293.865 286.275 -288.710 ;
        RECT 289.925 -289.235 290.320 -286.070 ;
        RECT 291.335 -287.315 291.565 -285.815 ;
        RECT 291.825 -287.315 292.055 -285.815 ;
        RECT 293.685 -287.315 293.915 -284.815 ;
        RECT 294.175 -287.315 294.405 -284.815 ;
        RECT 294.800 -287.315 295.030 -284.815 ;
        RECT 295.290 -287.315 295.520 -284.815 ;
        RECT 295.940 -287.315 296.170 -284.815 ;
        RECT 296.430 -287.315 296.660 -284.815 ;
        RECT 296.920 -287.315 297.150 -284.815 ;
        RECT 297.485 -284.845 305.595 -284.535 ;
        RECT 297.485 -284.890 297.815 -284.845 ;
        RECT 297.570 -287.315 297.800 -285.815 ;
        RECT 298.060 -287.315 298.290 -285.815 ;
        RECT 287.425 -289.630 290.320 -289.235 ;
        RECT 287.425 -291.405 287.820 -289.630 ;
        RECT 287.295 -291.890 287.875 -291.405 ;
        RECT 297.430 -292.045 299.625 -291.810 ;
        RECT 290.440 -292.125 290.925 -292.095 ;
        RECT 290.440 -292.395 295.985 -292.125 ;
        RECT 297.430 -292.230 297.665 -292.045 ;
        RECT 290.440 -292.425 290.925 -292.395 ;
        RECT 284.565 -294.430 288.105 -293.865 ;
        RECT 282.630 -295.105 282.860 -294.605 ;
        RECT 283.120 -295.250 283.350 -294.605 ;
        RECT 283.610 -295.105 283.840 -294.605 ;
        RECT 284.100 -295.250 284.330 -294.605 ;
        RECT 282.630 -295.480 285.815 -295.250 ;
        RECT 282.630 -296.260 282.860 -295.480 ;
        RECT 283.120 -295.490 284.330 -295.480 ;
        RECT 283.610 -296.260 283.840 -295.490 ;
        RECT 284.590 -296.260 284.820 -295.480 ;
        RECT 274.590 -300.755 274.820 -299.255 ;
        RECT 260.895 -304.100 262.385 -301.600 ;
        RECT 272.825 -301.730 273.810 -301.460 ;
        RECT 274.100 -303.435 274.330 -301.940 ;
        RECT 274.095 -303.620 274.330 -303.435 ;
        RECT 274.590 -303.440 274.820 -301.940 ;
        RECT 275.080 -303.620 275.310 -301.940 ;
        RECT 275.570 -303.440 275.800 -299.255 ;
        RECT 277.635 -300.030 277.865 -299.250 ;
        RECT 278.615 -300.020 278.845 -299.250 ;
        RECT 278.125 -300.030 279.335 -300.020 ;
        RECT 279.595 -300.030 279.825 -299.250 ;
        RECT 277.635 -300.260 280.820 -300.030 ;
        RECT 277.635 -300.905 277.865 -300.405 ;
        RECT 278.125 -300.905 278.355 -300.260 ;
        RECT 278.615 -300.905 278.845 -300.405 ;
        RECT 279.105 -300.905 279.335 -300.260 ;
        RECT 281.825 -301.810 282.055 -298.810 ;
        RECT 282.880 -301.810 283.110 -298.810 ;
        RECT 283.370 -301.810 283.600 -298.810 ;
        RECT 283.860 -301.810 284.090 -298.810 ;
        RECT 284.920 -301.810 285.150 -298.810 ;
        RECT 276.060 -303.620 276.290 -301.940 ;
        RECT 286.075 -302.465 286.600 -302.105 ;
        RECT 286.105 -302.880 286.430 -302.465 ;
        RECT 281.330 -303.205 286.430 -302.880 ;
        RECT 274.095 -303.855 276.290 -303.620 ;
        RECT 281.825 -304.870 282.055 -303.370 ;
        RECT 282.315 -304.870 282.545 -303.370 ;
        RECT 282.805 -304.870 283.035 -303.370 ;
        RECT 284.015 -304.870 284.245 -303.370 ;
        RECT 284.505 -304.870 284.735 -303.370 ;
        RECT 287.540 -305.410 288.105 -294.430 ;
        RECT 291.630 -294.595 292.280 -293.845 ;
        RECT 293.060 -294.115 293.290 -293.115 ;
        RECT 293.550 -294.255 293.780 -293.115 ;
        RECT 294.040 -294.115 294.270 -293.115 ;
        RECT 294.530 -294.255 294.760 -293.115 ;
        RECT 295.715 -293.845 295.985 -292.395 ;
        RECT 297.435 -293.725 297.665 -292.230 ;
        RECT 297.925 -293.725 298.155 -292.225 ;
        RECT 298.415 -293.725 298.645 -292.045 ;
        RECT 295.715 -294.115 297.355 -293.845 ;
        RECT 293.060 -294.485 296.245 -294.255 ;
        RECT 297.085 -294.390 297.355 -294.115 ;
        RECT 291.880 -301.615 292.150 -294.595 ;
        RECT 293.060 -295.765 293.290 -294.485 ;
        RECT 293.550 -294.495 294.760 -294.485 ;
        RECT 294.040 -295.765 294.270 -294.495 ;
        RECT 295.020 -295.765 295.250 -294.485 ;
        RECT 296.955 -294.680 297.750 -294.390 ;
        RECT 297.925 -296.410 298.155 -294.910 ;
        RECT 298.905 -296.410 299.135 -292.225 ;
        RECT 299.395 -293.725 299.625 -292.045 ;
        RECT 302.905 -294.585 306.445 -294.020 ;
        RECT 300.970 -295.260 301.200 -294.760 ;
        RECT 301.460 -295.405 301.690 -294.760 ;
        RECT 301.950 -295.260 302.180 -294.760 ;
        RECT 302.440 -295.405 302.670 -294.760 ;
        RECT 300.970 -295.635 304.155 -295.405 ;
        RECT 300.970 -296.415 301.200 -295.635 ;
        RECT 301.460 -295.645 302.670 -295.635 ;
        RECT 301.950 -296.415 302.180 -295.645 ;
        RECT 302.930 -296.415 303.160 -295.635 ;
        RECT 292.930 -300.910 293.160 -299.410 ;
        RECT 291.165 -301.885 292.150 -301.615 ;
        RECT 292.440 -303.590 292.670 -302.095 ;
        RECT 292.435 -303.775 292.670 -303.590 ;
        RECT 292.930 -303.595 293.160 -302.095 ;
        RECT 293.420 -303.775 293.650 -302.095 ;
        RECT 293.910 -303.595 294.140 -299.410 ;
        RECT 295.975 -300.185 296.205 -299.405 ;
        RECT 296.955 -300.175 297.185 -299.405 ;
        RECT 296.465 -300.185 297.675 -300.175 ;
        RECT 297.935 -300.185 298.165 -299.405 ;
        RECT 295.975 -300.415 299.160 -300.185 ;
        RECT 295.975 -301.060 296.205 -300.560 ;
        RECT 296.465 -301.060 296.695 -300.415 ;
        RECT 296.955 -301.060 297.185 -300.560 ;
        RECT 297.445 -301.060 297.675 -300.415 ;
        RECT 300.165 -301.965 300.395 -298.965 ;
        RECT 301.220 -301.965 301.450 -298.965 ;
        RECT 301.710 -301.965 301.940 -298.965 ;
        RECT 302.200 -301.965 302.430 -298.965 ;
        RECT 303.260 -301.965 303.490 -298.965 ;
        RECT 294.400 -303.775 294.630 -302.095 ;
        RECT 304.415 -302.620 304.940 -302.260 ;
        RECT 304.445 -303.035 304.770 -302.620 ;
        RECT 299.670 -303.360 304.770 -303.035 ;
        RECT 292.435 -304.010 294.630 -303.775 ;
        RECT 300.165 -305.025 300.395 -303.525 ;
        RECT 300.655 -305.025 300.885 -303.525 ;
        RECT 301.145 -305.025 301.375 -303.525 ;
        RECT 302.355 -305.025 302.585 -303.525 ;
        RECT 302.845 -305.025 303.075 -303.525 ;
        RECT 238.730 -306.145 260.455 -305.735 ;
        RECT 284.720 -305.565 288.105 -305.410 ;
        RECT 305.880 -305.565 306.445 -294.585 ;
        RECT 306.975 -302.290 308.080 -275.105 ;
        RECT 309.235 -290.970 310.425 -273.350 ;
        RECT 314.465 -274.375 315.715 -273.875 ;
        RECT 322.900 -274.295 325.095 -274.060 ;
        RECT 314.465 -274.645 321.455 -274.375 ;
        RECT 322.900 -274.480 323.135 -274.295 ;
        RECT 314.465 -275.020 315.715 -274.645 ;
        RECT 317.100 -276.845 317.750 -276.095 ;
        RECT 318.530 -276.365 318.760 -275.365 ;
        RECT 319.020 -276.505 319.250 -275.365 ;
        RECT 319.510 -276.365 319.740 -275.365 ;
        RECT 320.000 -276.505 320.230 -275.365 ;
        RECT 321.185 -276.095 321.455 -274.645 ;
        RECT 322.905 -275.975 323.135 -274.480 ;
        RECT 323.395 -275.975 323.625 -274.475 ;
        RECT 323.885 -275.975 324.115 -274.295 ;
        RECT 321.185 -276.365 322.825 -276.095 ;
        RECT 318.530 -276.735 321.715 -276.505 ;
        RECT 322.555 -276.640 322.825 -276.365 ;
        RECT 317.350 -283.865 317.620 -276.845 ;
        RECT 318.530 -278.015 318.760 -276.735 ;
        RECT 319.020 -276.745 320.230 -276.735 ;
        RECT 319.510 -278.015 319.740 -276.745 ;
        RECT 320.490 -278.015 320.720 -276.735 ;
        RECT 322.425 -276.930 323.220 -276.640 ;
        RECT 323.395 -278.660 323.625 -277.160 ;
        RECT 324.375 -278.660 324.605 -274.475 ;
        RECT 324.865 -275.975 325.095 -274.295 ;
        RECT 328.375 -276.835 331.915 -276.270 ;
        RECT 326.440 -277.510 326.670 -277.010 ;
        RECT 326.930 -277.655 327.160 -277.010 ;
        RECT 327.420 -277.510 327.650 -277.010 ;
        RECT 327.910 -277.655 328.140 -277.010 ;
        RECT 326.440 -277.885 329.625 -277.655 ;
        RECT 326.440 -278.665 326.670 -277.885 ;
        RECT 326.930 -277.895 328.140 -277.885 ;
        RECT 327.420 -278.665 327.650 -277.895 ;
        RECT 328.400 -278.665 328.630 -277.885 ;
        RECT 318.400 -283.160 318.630 -281.660 ;
        RECT 316.635 -284.135 317.620 -283.865 ;
        RECT 317.910 -285.840 318.140 -284.345 ;
        RECT 317.905 -286.025 318.140 -285.840 ;
        RECT 318.400 -285.845 318.630 -284.345 ;
        RECT 318.890 -286.025 319.120 -284.345 ;
        RECT 319.380 -285.845 319.610 -281.660 ;
        RECT 321.445 -282.435 321.675 -281.655 ;
        RECT 322.425 -282.425 322.655 -281.655 ;
        RECT 321.935 -282.435 323.145 -282.425 ;
        RECT 323.405 -282.435 323.635 -281.655 ;
        RECT 321.445 -282.665 324.630 -282.435 ;
        RECT 321.445 -283.310 321.675 -282.810 ;
        RECT 321.935 -283.310 322.165 -282.665 ;
        RECT 322.425 -283.310 322.655 -282.810 ;
        RECT 322.915 -283.310 323.145 -282.665 ;
        RECT 325.635 -284.215 325.865 -281.215 ;
        RECT 326.690 -284.215 326.920 -281.215 ;
        RECT 327.180 -284.215 327.410 -281.215 ;
        RECT 327.670 -284.215 327.900 -281.215 ;
        RECT 328.730 -284.215 328.960 -281.215 ;
        RECT 319.870 -286.025 320.100 -284.345 ;
        RECT 329.885 -284.870 330.410 -284.510 ;
        RECT 329.915 -285.285 330.240 -284.870 ;
        RECT 325.140 -285.610 330.240 -285.285 ;
        RECT 317.905 -286.260 320.100 -286.025 ;
        RECT 325.635 -287.275 325.865 -285.775 ;
        RECT 326.125 -287.275 326.355 -285.775 ;
        RECT 326.615 -287.275 326.845 -285.775 ;
        RECT 327.825 -287.275 328.055 -285.775 ;
        RECT 328.315 -287.275 328.545 -285.775 ;
        RECT 329.480 -287.815 330.045 -287.810 ;
        RECT 331.350 -287.815 331.915 -276.835 ;
        RECT 335.595 -283.005 335.825 -280.505 ;
        RECT 336.940 -283.005 337.170 -280.505 ;
        RECT 337.430 -283.005 337.660 -280.505 ;
        RECT 337.920 -283.005 338.150 -280.505 ;
        RECT 338.570 -283.005 338.800 -280.505 ;
        RECT 340.200 -283.005 340.430 -280.505 ;
        RECT 341.340 -282.005 341.570 -280.505 ;
        RECT 334.440 -283.805 335.130 -283.785 ;
        RECT 338.470 -283.805 339.160 -283.785 ;
        RECT 340.395 -283.805 340.665 -283.440 ;
        RECT 334.440 -284.025 340.665 -283.805 ;
        RECT 334.440 -284.055 335.130 -284.025 ;
        RECT 338.470 -284.055 339.160 -284.025 ;
        RECT 340.395 -284.130 340.665 -284.025 ;
        RECT 341.255 -284.205 341.585 -284.145 ;
        RECT 347.965 -284.205 349.155 -273.350 ;
        RECT 350.740 -273.560 351.625 -257.650 ;
        RECT 353.165 -273.390 395.105 -271.890 ;
        RECT 350.340 -275.015 352.030 -273.560 ;
        RECT 333.635 -285.740 334.150 -285.285 ;
        RECT 328.530 -288.380 331.915 -287.815 ;
        RECT 309.235 -291.640 314.915 -290.970 ;
        RECT 322.860 -291.560 325.055 -291.325 ;
        RECT 309.235 -291.910 321.415 -291.640 ;
        RECT 322.860 -291.745 323.095 -291.560 ;
        RECT 309.235 -292.160 314.915 -291.910 ;
        RECT 317.060 -294.110 317.710 -293.360 ;
        RECT 318.490 -293.630 318.720 -292.630 ;
        RECT 318.980 -293.770 319.210 -292.630 ;
        RECT 319.470 -293.630 319.700 -292.630 ;
        RECT 319.960 -293.770 320.190 -292.630 ;
        RECT 321.145 -293.360 321.415 -291.910 ;
        RECT 322.865 -293.240 323.095 -291.745 ;
        RECT 323.355 -293.240 323.585 -291.740 ;
        RECT 323.845 -293.240 324.075 -291.560 ;
        RECT 321.145 -293.630 322.785 -293.360 ;
        RECT 318.490 -294.000 321.675 -293.770 ;
        RECT 322.515 -293.905 322.785 -293.630 ;
        RECT 317.310 -301.130 317.580 -294.110 ;
        RECT 318.490 -295.280 318.720 -294.000 ;
        RECT 318.980 -294.010 320.190 -294.000 ;
        RECT 319.470 -295.280 319.700 -294.010 ;
        RECT 320.450 -295.280 320.680 -294.000 ;
        RECT 322.385 -294.195 323.180 -293.905 ;
        RECT 323.355 -295.925 323.585 -294.425 ;
        RECT 324.335 -295.925 324.565 -291.740 ;
        RECT 324.825 -293.240 325.055 -291.560 ;
        RECT 329.480 -293.535 330.045 -288.380 ;
        RECT 333.695 -288.905 334.090 -285.740 ;
        RECT 335.105 -286.985 335.335 -285.485 ;
        RECT 335.595 -286.985 335.825 -285.485 ;
        RECT 337.455 -286.985 337.685 -284.485 ;
        RECT 337.945 -286.985 338.175 -284.485 ;
        RECT 338.570 -286.985 338.800 -284.485 ;
        RECT 339.060 -286.985 339.290 -284.485 ;
        RECT 339.710 -286.985 339.940 -284.485 ;
        RECT 340.200 -286.985 340.430 -284.485 ;
        RECT 340.690 -286.985 340.920 -284.485 ;
        RECT 341.255 -284.515 349.365 -284.205 ;
        RECT 341.255 -284.560 341.585 -284.515 ;
        RECT 341.340 -286.985 341.570 -285.485 ;
        RECT 341.830 -286.985 342.060 -285.485 ;
        RECT 331.195 -289.300 334.090 -288.905 ;
        RECT 331.195 -291.075 331.590 -289.300 ;
        RECT 331.065 -291.560 331.645 -291.075 ;
        RECT 341.200 -291.715 343.395 -291.480 ;
        RECT 334.210 -291.795 334.695 -291.765 ;
        RECT 334.210 -292.065 339.755 -291.795 ;
        RECT 341.200 -291.900 341.435 -291.715 ;
        RECT 334.210 -292.095 334.695 -292.065 ;
        RECT 328.335 -294.100 331.875 -293.535 ;
        RECT 326.400 -294.775 326.630 -294.275 ;
        RECT 326.890 -294.920 327.120 -294.275 ;
        RECT 327.380 -294.775 327.610 -294.275 ;
        RECT 327.870 -294.920 328.100 -294.275 ;
        RECT 326.400 -295.150 329.585 -294.920 ;
        RECT 326.400 -295.930 326.630 -295.150 ;
        RECT 326.890 -295.160 328.100 -295.150 ;
        RECT 327.380 -295.930 327.610 -295.160 ;
        RECT 328.360 -295.930 328.590 -295.150 ;
        RECT 318.360 -300.425 318.590 -298.925 ;
        RECT 316.595 -301.400 317.580 -301.130 ;
        RECT 306.705 -303.785 308.165 -302.290 ;
        RECT 317.870 -303.105 318.100 -301.610 ;
        RECT 317.865 -303.290 318.100 -303.105 ;
        RECT 318.360 -303.110 318.590 -301.610 ;
        RECT 318.850 -303.290 319.080 -301.610 ;
        RECT 319.340 -303.110 319.570 -298.925 ;
        RECT 321.405 -299.700 321.635 -298.920 ;
        RECT 322.385 -299.690 322.615 -298.920 ;
        RECT 321.895 -299.700 323.105 -299.690 ;
        RECT 323.365 -299.700 323.595 -298.920 ;
        RECT 321.405 -299.930 324.590 -299.700 ;
        RECT 321.405 -300.575 321.635 -300.075 ;
        RECT 321.895 -300.575 322.125 -299.930 ;
        RECT 322.385 -300.575 322.615 -300.075 ;
        RECT 322.875 -300.575 323.105 -299.930 ;
        RECT 325.595 -301.480 325.825 -298.480 ;
        RECT 326.650 -301.480 326.880 -298.480 ;
        RECT 327.140 -301.480 327.370 -298.480 ;
        RECT 327.630 -301.480 327.860 -298.480 ;
        RECT 328.690 -301.480 328.920 -298.480 ;
        RECT 319.830 -303.290 320.060 -301.610 ;
        RECT 329.845 -302.135 330.370 -301.775 ;
        RECT 329.875 -302.550 330.200 -302.135 ;
        RECT 325.100 -302.875 330.200 -302.550 ;
        RECT 317.865 -303.525 320.060 -303.290 ;
        RECT 325.595 -304.540 325.825 -303.040 ;
        RECT 326.085 -304.540 326.315 -303.040 ;
        RECT 326.575 -304.540 326.805 -303.040 ;
        RECT 327.785 -304.540 328.015 -303.040 ;
        RECT 328.275 -304.540 328.505 -303.040 ;
        RECT 331.310 -305.080 331.875 -294.100 ;
        RECT 335.400 -294.265 336.050 -293.515 ;
        RECT 336.830 -293.785 337.060 -292.785 ;
        RECT 337.320 -293.925 337.550 -292.785 ;
        RECT 337.810 -293.785 338.040 -292.785 ;
        RECT 338.300 -293.925 338.530 -292.785 ;
        RECT 339.485 -293.515 339.755 -292.065 ;
        RECT 341.205 -293.395 341.435 -291.900 ;
        RECT 341.695 -293.395 341.925 -291.895 ;
        RECT 342.185 -293.395 342.415 -291.715 ;
        RECT 339.485 -293.785 341.125 -293.515 ;
        RECT 336.830 -294.155 340.015 -293.925 ;
        RECT 340.855 -294.060 341.125 -293.785 ;
        RECT 335.650 -301.285 335.920 -294.265 ;
        RECT 336.830 -295.435 337.060 -294.155 ;
        RECT 337.320 -294.165 338.530 -294.155 ;
        RECT 337.810 -295.435 338.040 -294.165 ;
        RECT 338.790 -295.435 339.020 -294.155 ;
        RECT 340.725 -294.350 341.520 -294.060 ;
        RECT 341.695 -296.080 341.925 -294.580 ;
        RECT 342.675 -296.080 342.905 -291.895 ;
        RECT 343.165 -293.395 343.395 -291.715 ;
        RECT 346.675 -294.255 350.215 -293.690 ;
        RECT 344.740 -294.930 344.970 -294.430 ;
        RECT 345.230 -295.075 345.460 -294.430 ;
        RECT 345.720 -294.930 345.950 -294.430 ;
        RECT 346.210 -295.075 346.440 -294.430 ;
        RECT 344.740 -295.305 347.925 -295.075 ;
        RECT 344.740 -296.085 344.970 -295.305 ;
        RECT 345.230 -295.315 346.440 -295.305 ;
        RECT 345.720 -296.085 345.950 -295.315 ;
        RECT 346.700 -296.085 346.930 -295.305 ;
        RECT 336.700 -300.580 336.930 -299.080 ;
        RECT 334.935 -301.555 335.920 -301.285 ;
        RECT 336.210 -303.260 336.440 -301.765 ;
        RECT 336.205 -303.445 336.440 -303.260 ;
        RECT 336.700 -303.265 336.930 -301.765 ;
        RECT 337.190 -303.445 337.420 -301.765 ;
        RECT 337.680 -303.265 337.910 -299.080 ;
        RECT 339.745 -299.855 339.975 -299.075 ;
        RECT 340.725 -299.845 340.955 -299.075 ;
        RECT 340.235 -299.855 341.445 -299.845 ;
        RECT 341.705 -299.855 341.935 -299.075 ;
        RECT 339.745 -300.085 342.930 -299.855 ;
        RECT 339.745 -300.730 339.975 -300.230 ;
        RECT 340.235 -300.730 340.465 -300.085 ;
        RECT 340.725 -300.730 340.955 -300.230 ;
        RECT 341.215 -300.730 341.445 -300.085 ;
        RECT 343.935 -301.635 344.165 -298.635 ;
        RECT 344.990 -301.635 345.220 -298.635 ;
        RECT 345.480 -301.635 345.710 -298.635 ;
        RECT 345.970 -301.635 346.200 -298.635 ;
        RECT 347.030 -301.635 347.260 -298.635 ;
        RECT 338.170 -303.445 338.400 -301.765 ;
        RECT 348.185 -302.290 348.710 -301.930 ;
        RECT 348.215 -302.705 348.540 -302.290 ;
        RECT 343.440 -303.030 348.540 -302.705 ;
        RECT 336.205 -303.680 338.400 -303.445 ;
        RECT 343.935 -304.695 344.165 -303.195 ;
        RECT 344.425 -304.695 344.655 -303.195 ;
        RECT 344.915 -304.695 345.145 -303.195 ;
        RECT 346.125 -304.695 346.355 -303.195 ;
        RECT 346.615 -304.695 346.845 -303.195 ;
        RECT 284.720 -305.975 306.445 -305.565 ;
        RECT 328.490 -305.235 331.875 -305.080 ;
        RECT 349.650 -305.235 350.215 -294.255 ;
        RECT 350.740 -302.000 351.625 -275.015 ;
        RECT 353.165 -290.640 354.665 -273.390 ;
        RECT 360.280 -274.290 361.620 -273.835 ;
        RECT 368.665 -274.210 370.860 -273.975 ;
        RECT 360.280 -274.560 367.220 -274.290 ;
        RECT 368.665 -274.395 368.900 -274.210 ;
        RECT 360.280 -275.035 361.620 -274.560 ;
        RECT 362.865 -276.760 363.515 -276.010 ;
        RECT 364.295 -276.280 364.525 -275.280 ;
        RECT 364.785 -276.420 365.015 -275.280 ;
        RECT 365.275 -276.280 365.505 -275.280 ;
        RECT 365.765 -276.420 365.995 -275.280 ;
        RECT 366.950 -276.010 367.220 -274.560 ;
        RECT 368.670 -275.890 368.900 -274.395 ;
        RECT 369.160 -275.890 369.390 -274.390 ;
        RECT 369.650 -275.890 369.880 -274.210 ;
        RECT 366.950 -276.280 368.590 -276.010 ;
        RECT 364.295 -276.650 367.480 -276.420 ;
        RECT 368.320 -276.555 368.590 -276.280 ;
        RECT 363.115 -283.780 363.385 -276.760 ;
        RECT 364.295 -277.930 364.525 -276.650 ;
        RECT 364.785 -276.660 365.995 -276.650 ;
        RECT 365.275 -277.930 365.505 -276.660 ;
        RECT 366.255 -277.930 366.485 -276.650 ;
        RECT 368.190 -276.845 368.985 -276.555 ;
        RECT 369.160 -278.575 369.390 -277.075 ;
        RECT 370.140 -278.575 370.370 -274.390 ;
        RECT 370.630 -275.890 370.860 -274.210 ;
        RECT 374.140 -276.750 377.680 -276.185 ;
        RECT 372.205 -277.425 372.435 -276.925 ;
        RECT 372.695 -277.570 372.925 -276.925 ;
        RECT 373.185 -277.425 373.415 -276.925 ;
        RECT 373.675 -277.570 373.905 -276.925 ;
        RECT 372.205 -277.800 375.390 -277.570 ;
        RECT 372.205 -278.580 372.435 -277.800 ;
        RECT 372.695 -277.810 373.905 -277.800 ;
        RECT 373.185 -278.580 373.415 -277.810 ;
        RECT 374.165 -278.580 374.395 -277.800 ;
        RECT 364.165 -283.075 364.395 -281.575 ;
        RECT 362.400 -284.050 363.385 -283.780 ;
        RECT 363.675 -285.755 363.905 -284.260 ;
        RECT 363.670 -285.940 363.905 -285.755 ;
        RECT 364.165 -285.760 364.395 -284.260 ;
        RECT 364.655 -285.940 364.885 -284.260 ;
        RECT 365.145 -285.760 365.375 -281.575 ;
        RECT 367.210 -282.350 367.440 -281.570 ;
        RECT 368.190 -282.340 368.420 -281.570 ;
        RECT 367.700 -282.350 368.910 -282.340 ;
        RECT 369.170 -282.350 369.400 -281.570 ;
        RECT 367.210 -282.580 370.395 -282.350 ;
        RECT 367.210 -283.225 367.440 -282.725 ;
        RECT 367.700 -283.225 367.930 -282.580 ;
        RECT 368.190 -283.225 368.420 -282.725 ;
        RECT 368.680 -283.225 368.910 -282.580 ;
        RECT 371.400 -284.130 371.630 -281.130 ;
        RECT 372.455 -284.130 372.685 -281.130 ;
        RECT 372.945 -284.130 373.175 -281.130 ;
        RECT 373.435 -284.130 373.665 -281.130 ;
        RECT 374.495 -284.130 374.725 -281.130 ;
        RECT 365.635 -285.940 365.865 -284.260 ;
        RECT 375.650 -284.785 376.175 -284.425 ;
        RECT 375.680 -285.200 376.005 -284.785 ;
        RECT 370.905 -285.525 376.005 -285.200 ;
        RECT 363.670 -286.175 365.865 -285.940 ;
        RECT 371.400 -287.190 371.630 -285.690 ;
        RECT 371.890 -287.190 372.120 -285.690 ;
        RECT 372.380 -287.190 372.610 -285.690 ;
        RECT 373.590 -287.190 373.820 -285.690 ;
        RECT 374.080 -287.190 374.310 -285.690 ;
        RECT 375.245 -287.730 375.810 -287.725 ;
        RECT 377.115 -287.730 377.680 -276.750 ;
        RECT 381.360 -282.920 381.590 -280.420 ;
        RECT 382.705 -282.920 382.935 -280.420 ;
        RECT 383.195 -282.920 383.425 -280.420 ;
        RECT 383.685 -282.920 383.915 -280.420 ;
        RECT 384.335 -282.920 384.565 -280.420 ;
        RECT 385.965 -282.920 386.195 -280.420 ;
        RECT 387.105 -281.920 387.335 -280.420 ;
        RECT 380.205 -283.720 380.895 -283.700 ;
        RECT 384.235 -283.720 384.925 -283.700 ;
        RECT 386.160 -283.720 386.430 -283.355 ;
        RECT 380.205 -283.940 386.430 -283.720 ;
        RECT 380.205 -283.970 380.895 -283.940 ;
        RECT 384.235 -283.970 384.925 -283.940 ;
        RECT 386.160 -284.045 386.430 -283.940 ;
        RECT 387.020 -284.120 387.350 -284.060 ;
        RECT 393.570 -284.120 395.105 -273.390 ;
        RECT 379.400 -285.655 379.915 -285.200 ;
        RECT 374.295 -288.295 377.680 -287.730 ;
        RECT 353.165 -291.555 360.615 -290.640 ;
        RECT 368.625 -291.475 370.820 -291.240 ;
        RECT 353.165 -291.825 367.180 -291.555 ;
        RECT 368.625 -291.660 368.860 -291.475 ;
        RECT 353.165 -292.140 360.615 -291.825 ;
        RECT 362.825 -294.025 363.475 -293.275 ;
        RECT 364.255 -293.545 364.485 -292.545 ;
        RECT 364.745 -293.685 364.975 -292.545 ;
        RECT 365.235 -293.545 365.465 -292.545 ;
        RECT 365.725 -293.685 365.955 -292.545 ;
        RECT 366.910 -293.275 367.180 -291.825 ;
        RECT 368.630 -293.155 368.860 -291.660 ;
        RECT 369.120 -293.155 369.350 -291.655 ;
        RECT 369.610 -293.155 369.840 -291.475 ;
        RECT 366.910 -293.545 368.550 -293.275 ;
        RECT 364.255 -293.915 367.440 -293.685 ;
        RECT 368.280 -293.820 368.550 -293.545 ;
        RECT 363.075 -301.045 363.345 -294.025 ;
        RECT 364.255 -295.195 364.485 -293.915 ;
        RECT 364.745 -293.925 365.955 -293.915 ;
        RECT 365.235 -295.195 365.465 -293.925 ;
        RECT 366.215 -295.195 366.445 -293.915 ;
        RECT 368.150 -294.110 368.945 -293.820 ;
        RECT 369.120 -295.840 369.350 -294.340 ;
        RECT 370.100 -295.840 370.330 -291.655 ;
        RECT 370.590 -293.155 370.820 -291.475 ;
        RECT 375.245 -293.450 375.810 -288.295 ;
        RECT 379.460 -288.820 379.855 -285.655 ;
        RECT 380.870 -286.900 381.100 -285.400 ;
        RECT 381.360 -286.900 381.590 -285.400 ;
        RECT 383.220 -286.900 383.450 -284.400 ;
        RECT 383.710 -286.900 383.940 -284.400 ;
        RECT 384.335 -286.900 384.565 -284.400 ;
        RECT 384.825 -286.900 385.055 -284.400 ;
        RECT 385.475 -286.900 385.705 -284.400 ;
        RECT 385.965 -286.900 386.195 -284.400 ;
        RECT 386.455 -286.900 386.685 -284.400 ;
        RECT 387.020 -284.430 395.130 -284.120 ;
        RECT 387.020 -284.475 387.350 -284.430 ;
        RECT 387.105 -286.900 387.335 -285.400 ;
        RECT 387.595 -286.900 387.825 -285.400 ;
        RECT 376.960 -289.215 379.855 -288.820 ;
        RECT 376.960 -290.990 377.355 -289.215 ;
        RECT 376.830 -291.475 377.410 -290.990 ;
        RECT 386.965 -291.630 389.160 -291.395 ;
        RECT 379.975 -291.710 380.460 -291.680 ;
        RECT 379.975 -291.980 385.520 -291.710 ;
        RECT 386.965 -291.815 387.200 -291.630 ;
        RECT 379.975 -292.010 380.460 -291.980 ;
        RECT 374.100 -294.015 377.640 -293.450 ;
        RECT 372.165 -294.690 372.395 -294.190 ;
        RECT 372.655 -294.835 372.885 -294.190 ;
        RECT 373.145 -294.690 373.375 -294.190 ;
        RECT 373.635 -294.835 373.865 -294.190 ;
        RECT 372.165 -295.065 375.350 -294.835 ;
        RECT 372.165 -295.845 372.395 -295.065 ;
        RECT 372.655 -295.075 373.865 -295.065 ;
        RECT 373.145 -295.845 373.375 -295.075 ;
        RECT 374.125 -295.845 374.355 -295.065 ;
        RECT 364.125 -300.340 364.355 -298.840 ;
        RECT 362.360 -301.315 363.345 -301.045 ;
        RECT 350.530 -303.520 351.835 -302.000 ;
        RECT 363.635 -303.020 363.865 -301.525 ;
        RECT 363.630 -303.205 363.865 -303.020 ;
        RECT 364.125 -303.025 364.355 -301.525 ;
        RECT 364.615 -303.205 364.845 -301.525 ;
        RECT 365.105 -303.025 365.335 -298.840 ;
        RECT 367.170 -299.615 367.400 -298.835 ;
        RECT 368.150 -299.605 368.380 -298.835 ;
        RECT 367.660 -299.615 368.870 -299.605 ;
        RECT 369.130 -299.615 369.360 -298.835 ;
        RECT 367.170 -299.845 370.355 -299.615 ;
        RECT 367.170 -300.490 367.400 -299.990 ;
        RECT 367.660 -300.490 367.890 -299.845 ;
        RECT 368.150 -300.490 368.380 -299.990 ;
        RECT 368.640 -300.490 368.870 -299.845 ;
        RECT 371.360 -301.395 371.590 -298.395 ;
        RECT 372.415 -301.395 372.645 -298.395 ;
        RECT 372.905 -301.395 373.135 -298.395 ;
        RECT 373.395 -301.395 373.625 -298.395 ;
        RECT 374.455 -301.395 374.685 -298.395 ;
        RECT 365.595 -303.205 365.825 -301.525 ;
        RECT 375.610 -302.050 376.135 -301.690 ;
        RECT 375.640 -302.465 375.965 -302.050 ;
        RECT 370.865 -302.790 375.965 -302.465 ;
        RECT 363.630 -303.440 365.825 -303.205 ;
        RECT 371.360 -304.455 371.590 -302.955 ;
        RECT 371.850 -304.455 372.080 -302.955 ;
        RECT 372.340 -304.455 372.570 -302.955 ;
        RECT 373.550 -304.455 373.780 -302.955 ;
        RECT 374.040 -304.455 374.270 -302.955 ;
        RECT 377.075 -304.995 377.640 -294.015 ;
        RECT 381.165 -294.180 381.815 -293.430 ;
        RECT 382.595 -293.700 382.825 -292.700 ;
        RECT 383.085 -293.840 383.315 -292.700 ;
        RECT 383.575 -293.700 383.805 -292.700 ;
        RECT 384.065 -293.840 384.295 -292.700 ;
        RECT 385.250 -293.430 385.520 -291.980 ;
        RECT 386.970 -293.310 387.200 -291.815 ;
        RECT 387.460 -293.310 387.690 -291.810 ;
        RECT 387.950 -293.310 388.180 -291.630 ;
        RECT 385.250 -293.700 386.890 -293.430 ;
        RECT 382.595 -294.070 385.780 -293.840 ;
        RECT 386.620 -293.975 386.890 -293.700 ;
        RECT 381.415 -301.200 381.685 -294.180 ;
        RECT 382.595 -295.350 382.825 -294.070 ;
        RECT 383.085 -294.080 384.295 -294.070 ;
        RECT 383.575 -295.350 383.805 -294.080 ;
        RECT 384.555 -295.350 384.785 -294.070 ;
        RECT 386.490 -294.265 387.285 -293.975 ;
        RECT 387.460 -295.995 387.690 -294.495 ;
        RECT 388.440 -295.995 388.670 -291.810 ;
        RECT 388.930 -293.310 389.160 -291.630 ;
        RECT 392.440 -294.170 395.980 -293.605 ;
        RECT 390.505 -294.845 390.735 -294.345 ;
        RECT 390.995 -294.990 391.225 -294.345 ;
        RECT 391.485 -294.845 391.715 -294.345 ;
        RECT 391.975 -294.990 392.205 -294.345 ;
        RECT 390.505 -295.220 393.690 -294.990 ;
        RECT 390.505 -296.000 390.735 -295.220 ;
        RECT 390.995 -295.230 392.205 -295.220 ;
        RECT 391.485 -296.000 391.715 -295.230 ;
        RECT 392.465 -296.000 392.695 -295.220 ;
        RECT 382.465 -300.495 382.695 -298.995 ;
        RECT 380.700 -301.470 381.685 -301.200 ;
        RECT 381.975 -303.175 382.205 -301.680 ;
        RECT 381.970 -303.360 382.205 -303.175 ;
        RECT 382.465 -303.180 382.695 -301.680 ;
        RECT 382.955 -303.360 383.185 -301.680 ;
        RECT 383.445 -303.180 383.675 -298.995 ;
        RECT 385.510 -299.770 385.740 -298.990 ;
        RECT 386.490 -299.760 386.720 -298.990 ;
        RECT 386.000 -299.770 387.210 -299.760 ;
        RECT 387.470 -299.770 387.700 -298.990 ;
        RECT 385.510 -300.000 388.695 -299.770 ;
        RECT 385.510 -300.645 385.740 -300.145 ;
        RECT 386.000 -300.645 386.230 -300.000 ;
        RECT 386.490 -300.645 386.720 -300.145 ;
        RECT 386.980 -300.645 387.210 -300.000 ;
        RECT 389.700 -301.550 389.930 -298.550 ;
        RECT 390.755 -301.550 390.985 -298.550 ;
        RECT 391.245 -301.550 391.475 -298.550 ;
        RECT 391.735 -301.550 391.965 -298.550 ;
        RECT 392.795 -301.550 393.025 -298.550 ;
        RECT 383.935 -303.360 384.165 -301.680 ;
        RECT 393.950 -302.205 394.475 -301.845 ;
        RECT 393.980 -302.620 394.305 -302.205 ;
        RECT 389.205 -302.945 394.305 -302.620 ;
        RECT 381.970 -303.595 384.165 -303.360 ;
        RECT 389.700 -304.610 389.930 -303.110 ;
        RECT 390.190 -304.610 390.420 -303.110 ;
        RECT 390.680 -304.610 390.910 -303.110 ;
        RECT 391.890 -304.610 392.120 -303.110 ;
        RECT 392.380 -304.610 392.610 -303.110 ;
        RECT 328.490 -305.645 350.215 -305.235 ;
        RECT 374.255 -305.150 377.640 -304.995 ;
        RECT 395.415 -305.150 395.980 -294.170 ;
        RECT 396.410 -303.620 397.965 -255.400 ;
        RECT 399.290 -272.980 441.885 -271.885 ;
        RECT 399.290 -291.170 400.385 -272.980 ;
        RECT 406.555 -274.100 408.030 -273.525 ;
        RECT 415.485 -274.020 417.680 -273.785 ;
        RECT 406.555 -274.370 414.040 -274.100 ;
        RECT 415.485 -274.205 415.720 -274.020 ;
        RECT 406.555 -274.890 408.030 -274.370 ;
        RECT 409.685 -276.570 410.335 -275.820 ;
        RECT 411.115 -276.090 411.345 -275.090 ;
        RECT 411.605 -276.230 411.835 -275.090 ;
        RECT 412.095 -276.090 412.325 -275.090 ;
        RECT 412.585 -276.230 412.815 -275.090 ;
        RECT 413.770 -275.820 414.040 -274.370 ;
        RECT 415.490 -275.700 415.720 -274.205 ;
        RECT 415.980 -275.700 416.210 -274.200 ;
        RECT 416.470 -275.700 416.700 -274.020 ;
        RECT 413.770 -276.090 415.410 -275.820 ;
        RECT 411.115 -276.460 414.300 -276.230 ;
        RECT 415.140 -276.365 415.410 -276.090 ;
        RECT 409.935 -283.590 410.205 -276.570 ;
        RECT 411.115 -277.740 411.345 -276.460 ;
        RECT 411.605 -276.470 412.815 -276.460 ;
        RECT 412.095 -277.740 412.325 -276.470 ;
        RECT 413.075 -277.740 413.305 -276.460 ;
        RECT 415.010 -276.655 415.805 -276.365 ;
        RECT 415.980 -278.385 416.210 -276.885 ;
        RECT 416.960 -278.385 417.190 -274.200 ;
        RECT 417.450 -275.700 417.680 -274.020 ;
        RECT 420.960 -276.560 424.500 -275.995 ;
        RECT 419.025 -277.235 419.255 -276.735 ;
        RECT 419.515 -277.380 419.745 -276.735 ;
        RECT 420.005 -277.235 420.235 -276.735 ;
        RECT 420.495 -277.380 420.725 -276.735 ;
        RECT 419.025 -277.610 422.210 -277.380 ;
        RECT 419.025 -278.390 419.255 -277.610 ;
        RECT 419.515 -277.620 420.725 -277.610 ;
        RECT 420.005 -278.390 420.235 -277.620 ;
        RECT 420.985 -278.390 421.215 -277.610 ;
        RECT 410.985 -282.885 411.215 -281.385 ;
        RECT 409.220 -283.860 410.205 -283.590 ;
        RECT 410.495 -285.565 410.725 -284.070 ;
        RECT 410.490 -285.750 410.725 -285.565 ;
        RECT 410.985 -285.570 411.215 -284.070 ;
        RECT 411.475 -285.750 411.705 -284.070 ;
        RECT 411.965 -285.570 412.195 -281.385 ;
        RECT 414.030 -282.160 414.260 -281.380 ;
        RECT 415.010 -282.150 415.240 -281.380 ;
        RECT 414.520 -282.160 415.730 -282.150 ;
        RECT 415.990 -282.160 416.220 -281.380 ;
        RECT 414.030 -282.390 417.215 -282.160 ;
        RECT 414.030 -283.035 414.260 -282.535 ;
        RECT 414.520 -283.035 414.750 -282.390 ;
        RECT 415.010 -283.035 415.240 -282.535 ;
        RECT 415.500 -283.035 415.730 -282.390 ;
        RECT 418.220 -283.940 418.450 -280.940 ;
        RECT 419.275 -283.940 419.505 -280.940 ;
        RECT 419.765 -283.940 419.995 -280.940 ;
        RECT 420.255 -283.940 420.485 -280.940 ;
        RECT 421.315 -283.940 421.545 -280.940 ;
        RECT 412.455 -285.750 412.685 -284.070 ;
        RECT 422.470 -284.595 422.995 -284.235 ;
        RECT 422.500 -285.010 422.825 -284.595 ;
        RECT 417.725 -285.335 422.825 -285.010 ;
        RECT 410.490 -285.985 412.685 -285.750 ;
        RECT 418.220 -287.000 418.450 -285.500 ;
        RECT 418.710 -287.000 418.940 -285.500 ;
        RECT 419.200 -287.000 419.430 -285.500 ;
        RECT 420.410 -287.000 420.640 -285.500 ;
        RECT 420.900 -287.000 421.130 -285.500 ;
        RECT 422.065 -287.540 422.630 -287.535 ;
        RECT 423.935 -287.540 424.500 -276.560 ;
        RECT 428.180 -282.730 428.410 -280.230 ;
        RECT 429.525 -282.730 429.755 -280.230 ;
        RECT 430.015 -282.730 430.245 -280.230 ;
        RECT 430.505 -282.730 430.735 -280.230 ;
        RECT 431.155 -282.730 431.385 -280.230 ;
        RECT 432.785 -282.730 433.015 -280.230 ;
        RECT 433.925 -281.730 434.155 -280.230 ;
        RECT 427.025 -283.530 427.715 -283.510 ;
        RECT 431.055 -283.530 431.745 -283.510 ;
        RECT 432.980 -283.530 433.250 -283.165 ;
        RECT 427.025 -283.750 433.250 -283.530 ;
        RECT 427.025 -283.780 427.715 -283.750 ;
        RECT 431.055 -283.780 431.745 -283.750 ;
        RECT 432.980 -283.855 433.250 -283.750 ;
        RECT 433.840 -283.930 434.170 -283.870 ;
        RECT 440.790 -283.930 441.885 -272.980 ;
        RECT 426.220 -285.465 426.735 -285.010 ;
        RECT 421.115 -288.105 424.500 -287.540 ;
        RECT 399.290 -291.365 408.185 -291.170 ;
        RECT 415.445 -291.285 417.640 -291.050 ;
        RECT 399.290 -291.635 414.000 -291.365 ;
        RECT 415.445 -291.470 415.680 -291.285 ;
        RECT 399.290 -292.265 408.185 -291.635 ;
        RECT 409.645 -293.835 410.295 -293.085 ;
        RECT 411.075 -293.355 411.305 -292.355 ;
        RECT 411.565 -293.495 411.795 -292.355 ;
        RECT 412.055 -293.355 412.285 -292.355 ;
        RECT 412.545 -293.495 412.775 -292.355 ;
        RECT 413.730 -293.085 414.000 -291.635 ;
        RECT 415.450 -292.965 415.680 -291.470 ;
        RECT 415.940 -292.965 416.170 -291.465 ;
        RECT 416.430 -292.965 416.660 -291.285 ;
        RECT 413.730 -293.355 415.370 -293.085 ;
        RECT 411.075 -293.725 414.260 -293.495 ;
        RECT 415.100 -293.630 415.370 -293.355 ;
        RECT 409.895 -300.855 410.165 -293.835 ;
        RECT 411.075 -295.005 411.305 -293.725 ;
        RECT 411.565 -293.735 412.775 -293.725 ;
        RECT 412.055 -295.005 412.285 -293.735 ;
        RECT 413.035 -295.005 413.265 -293.725 ;
        RECT 414.970 -293.920 415.765 -293.630 ;
        RECT 415.940 -295.650 416.170 -294.150 ;
        RECT 416.920 -295.650 417.150 -291.465 ;
        RECT 417.410 -292.965 417.640 -291.285 ;
        RECT 422.065 -293.260 422.630 -288.105 ;
        RECT 426.280 -288.630 426.675 -285.465 ;
        RECT 427.690 -286.710 427.920 -285.210 ;
        RECT 428.180 -286.710 428.410 -285.210 ;
        RECT 430.040 -286.710 430.270 -284.210 ;
        RECT 430.530 -286.710 430.760 -284.210 ;
        RECT 431.155 -286.710 431.385 -284.210 ;
        RECT 431.645 -286.710 431.875 -284.210 ;
        RECT 432.295 -286.710 432.525 -284.210 ;
        RECT 432.785 -286.710 433.015 -284.210 ;
        RECT 433.275 -286.710 433.505 -284.210 ;
        RECT 433.840 -284.240 441.950 -283.930 ;
        RECT 433.840 -284.285 434.170 -284.240 ;
        RECT 433.925 -286.710 434.155 -285.210 ;
        RECT 434.415 -286.710 434.645 -285.210 ;
        RECT 423.780 -289.025 426.675 -288.630 ;
        RECT 423.780 -290.800 424.175 -289.025 ;
        RECT 423.650 -291.285 424.230 -290.800 ;
        RECT 433.785 -291.440 435.980 -291.205 ;
        RECT 426.795 -291.520 427.280 -291.490 ;
        RECT 426.795 -291.790 432.340 -291.520 ;
        RECT 433.785 -291.625 434.020 -291.440 ;
        RECT 426.795 -291.820 427.280 -291.790 ;
        RECT 420.920 -293.825 424.460 -293.260 ;
        RECT 418.985 -294.500 419.215 -294.000 ;
        RECT 419.475 -294.645 419.705 -294.000 ;
        RECT 419.965 -294.500 420.195 -294.000 ;
        RECT 420.455 -294.645 420.685 -294.000 ;
        RECT 418.985 -294.875 422.170 -294.645 ;
        RECT 418.985 -295.655 419.215 -294.875 ;
        RECT 419.475 -294.885 420.685 -294.875 ;
        RECT 419.965 -295.655 420.195 -294.885 ;
        RECT 420.945 -295.655 421.175 -294.875 ;
        RECT 410.945 -300.150 411.175 -298.650 ;
        RECT 409.180 -301.125 410.165 -300.855 ;
        RECT 410.455 -302.830 410.685 -301.335 ;
        RECT 410.450 -303.015 410.685 -302.830 ;
        RECT 410.945 -302.835 411.175 -301.335 ;
        RECT 411.435 -303.015 411.665 -301.335 ;
        RECT 411.925 -302.835 412.155 -298.650 ;
        RECT 413.990 -299.425 414.220 -298.645 ;
        RECT 414.970 -299.415 415.200 -298.645 ;
        RECT 414.480 -299.425 415.690 -299.415 ;
        RECT 415.950 -299.425 416.180 -298.645 ;
        RECT 413.990 -299.655 417.175 -299.425 ;
        RECT 413.990 -300.300 414.220 -299.800 ;
        RECT 414.480 -300.300 414.710 -299.655 ;
        RECT 414.970 -300.300 415.200 -299.800 ;
        RECT 415.460 -300.300 415.690 -299.655 ;
        RECT 418.180 -301.205 418.410 -298.205 ;
        RECT 419.235 -301.205 419.465 -298.205 ;
        RECT 419.725 -301.205 419.955 -298.205 ;
        RECT 420.215 -301.205 420.445 -298.205 ;
        RECT 421.275 -301.205 421.505 -298.205 ;
        RECT 412.415 -303.015 412.645 -301.335 ;
        RECT 422.430 -301.860 422.955 -301.500 ;
        RECT 422.460 -302.275 422.785 -301.860 ;
        RECT 417.685 -302.600 422.785 -302.275 ;
        RECT 410.450 -303.250 412.645 -303.015 ;
        RECT 418.180 -304.265 418.410 -302.765 ;
        RECT 418.670 -304.265 418.900 -302.765 ;
        RECT 419.160 -304.265 419.390 -302.765 ;
        RECT 420.370 -304.265 420.600 -302.765 ;
        RECT 420.860 -304.265 421.090 -302.765 ;
        RECT 423.895 -304.805 424.460 -293.825 ;
        RECT 427.985 -293.990 428.635 -293.240 ;
        RECT 429.415 -293.510 429.645 -292.510 ;
        RECT 429.905 -293.650 430.135 -292.510 ;
        RECT 430.395 -293.510 430.625 -292.510 ;
        RECT 430.885 -293.650 431.115 -292.510 ;
        RECT 432.070 -293.240 432.340 -291.790 ;
        RECT 433.790 -293.120 434.020 -291.625 ;
        RECT 434.280 -293.120 434.510 -291.620 ;
        RECT 434.770 -293.120 435.000 -291.440 ;
        RECT 432.070 -293.510 433.710 -293.240 ;
        RECT 429.415 -293.880 432.600 -293.650 ;
        RECT 433.440 -293.785 433.710 -293.510 ;
        RECT 428.235 -301.010 428.505 -293.990 ;
        RECT 429.415 -295.160 429.645 -293.880 ;
        RECT 429.905 -293.890 431.115 -293.880 ;
        RECT 430.395 -295.160 430.625 -293.890 ;
        RECT 431.375 -295.160 431.605 -293.880 ;
        RECT 433.310 -294.075 434.105 -293.785 ;
        RECT 434.280 -295.805 434.510 -294.305 ;
        RECT 435.260 -295.805 435.490 -291.620 ;
        RECT 435.750 -293.120 435.980 -291.440 ;
        RECT 439.260 -293.980 442.800 -293.415 ;
        RECT 437.325 -294.655 437.555 -294.155 ;
        RECT 437.815 -294.800 438.045 -294.155 ;
        RECT 438.305 -294.655 438.535 -294.155 ;
        RECT 438.795 -294.800 439.025 -294.155 ;
        RECT 437.325 -295.030 440.510 -294.800 ;
        RECT 437.325 -295.810 437.555 -295.030 ;
        RECT 437.815 -295.040 439.025 -295.030 ;
        RECT 438.305 -295.810 438.535 -295.040 ;
        RECT 439.285 -295.810 439.515 -295.030 ;
        RECT 429.285 -300.305 429.515 -298.805 ;
        RECT 427.520 -301.280 428.505 -301.010 ;
        RECT 428.795 -302.985 429.025 -301.490 ;
        RECT 428.790 -303.170 429.025 -302.985 ;
        RECT 429.285 -302.990 429.515 -301.490 ;
        RECT 429.775 -303.170 430.005 -301.490 ;
        RECT 430.265 -302.990 430.495 -298.805 ;
        RECT 432.330 -299.580 432.560 -298.800 ;
        RECT 433.310 -299.570 433.540 -298.800 ;
        RECT 432.820 -299.580 434.030 -299.570 ;
        RECT 434.290 -299.580 434.520 -298.800 ;
        RECT 432.330 -299.810 435.515 -299.580 ;
        RECT 432.330 -300.455 432.560 -299.955 ;
        RECT 432.820 -300.455 433.050 -299.810 ;
        RECT 433.310 -300.455 433.540 -299.955 ;
        RECT 433.800 -300.455 434.030 -299.810 ;
        RECT 436.520 -301.360 436.750 -298.360 ;
        RECT 437.575 -301.360 437.805 -298.360 ;
        RECT 438.065 -301.360 438.295 -298.360 ;
        RECT 438.555 -301.360 438.785 -298.360 ;
        RECT 439.615 -301.360 439.845 -298.360 ;
        RECT 430.755 -303.170 430.985 -301.490 ;
        RECT 440.770 -302.015 441.295 -301.655 ;
        RECT 440.800 -302.430 441.125 -302.015 ;
        RECT 436.025 -302.755 441.125 -302.430 ;
        RECT 428.790 -303.405 430.985 -303.170 ;
        RECT 436.520 -304.420 436.750 -302.920 ;
        RECT 437.010 -304.420 437.240 -302.920 ;
        RECT 437.500 -304.420 437.730 -302.920 ;
        RECT 438.710 -304.420 438.940 -302.920 ;
        RECT 439.200 -304.420 439.430 -302.920 ;
        RECT 374.255 -305.560 395.980 -305.150 ;
        RECT 421.075 -304.960 424.460 -304.805 ;
        RECT 442.235 -304.960 442.800 -293.980 ;
        RECT 444.065 -301.780 445.485 -250.735 ;
        RECT 443.915 -303.495 445.710 -301.780 ;
        RECT 421.075 -305.370 442.800 -304.960 ;
        RECT 421.095 -305.525 442.800 -305.370 ;
        RECT 328.510 -305.800 350.215 -305.645 ;
        RECT 374.275 -305.715 395.980 -305.560 ;
        RECT 284.740 -306.130 306.445 -305.975 ;
        RECT 238.750 -306.300 260.455 -306.145 ;
        RECT 214.890 -309.170 216.475 -308.755 ;
        RECT 136.390 -310.075 180.390 -309.170 ;
        RECT 214.890 -310.075 413.640 -309.170 ;
        RECT 214.890 -310.210 216.475 -310.075 ;
        RECT 214.675 -314.670 216.520 -312.785 ;
        RECT 221.275 -314.275 413.640 -312.850 ;
        RECT 214.720 -323.610 216.220 -314.670 ;
        RECT 127.330 -325.110 216.220 -323.610 ;
        RECT 221.275 -326.325 222.700 -314.275 ;
        RECT 126.305 -326.620 222.700 -326.325 ;
        RECT 124.990 -327.225 222.700 -326.620 ;
        RECT 126.305 -327.750 222.700 -327.225 ;
      LAYER met2 ;
        RECT 469.655 62.300 475.760 192.475 ;
        RECT -0.785 54.610 0.435 62.285 ;
        RECT 7.495 9.270 8.590 9.665 ;
        RECT 8.175 4.655 8.590 9.270 ;
      LAYER met3 ;
        RECT 469.655 62.300 475.760 192.475 ;
        RECT -0.785 54.610 0.435 62.285 ;
      LAYER met4 ;
        RECT 91.695 432.280 116.305 444.325 ;
        RECT 118.295 432.280 142.905 444.325 ;
        RECT 144.895 432.280 169.505 444.325 ;
        RECT 171.495 432.280 196.105 444.325 ;
        RECT 198.095 432.280 222.705 444.325 ;
        RECT 224.695 432.280 249.305 444.325 ;
        RECT 251.295 432.280 275.905 444.325 ;
        RECT 277.895 432.280 302.505 444.325 ;
        RECT 304.495 432.280 329.105 444.325 ;
        RECT 331.095 432.280 355.705 444.325 ;
        RECT 357.695 432.280 382.305 444.325 ;
        RECT 384.295 432.280 408.905 444.325 ;
        RECT 410.895 432.280 435.505 444.325 ;
        RECT 437.495 432.280 462.105 444.325 ;
        RECT 467.885 432.280 478.000 445.340 ;
        RECT 90.700 431.760 478.000 432.280 ;
        RECT 91.695 419.715 116.305 431.760 ;
        RECT 118.295 419.715 142.905 431.760 ;
        RECT 144.895 419.715 169.505 431.760 ;
        RECT 171.495 419.715 196.105 431.760 ;
        RECT 198.095 419.715 222.705 431.760 ;
        RECT 224.695 419.715 249.305 431.760 ;
        RECT 251.295 419.715 275.905 431.760 ;
        RECT 277.895 419.715 302.505 431.760 ;
        RECT 304.495 419.715 329.105 431.760 ;
        RECT 331.095 419.715 355.705 431.760 ;
        RECT 357.695 419.715 382.305 431.760 ;
        RECT 384.295 419.715 408.905 431.760 ;
        RECT 410.895 419.715 435.505 431.760 ;
        RECT 437.495 419.715 462.105 431.760 ;
        RECT 91.695 404.220 116.305 416.265 ;
        RECT 118.295 404.220 142.905 416.265 ;
        RECT 144.895 404.220 169.505 416.265 ;
        RECT 171.495 404.220 196.105 416.265 ;
        RECT 198.095 404.220 222.705 416.265 ;
        RECT 224.695 404.220 249.305 416.265 ;
        RECT 251.295 404.220 275.905 416.265 ;
        RECT 277.895 404.220 302.505 416.265 ;
        RECT 304.495 404.220 329.105 416.265 ;
        RECT 331.095 404.220 355.705 416.265 ;
        RECT 357.695 404.220 382.305 416.265 ;
        RECT 384.295 404.220 408.905 416.265 ;
        RECT 410.895 404.220 435.505 416.265 ;
        RECT 437.495 404.220 462.105 416.265 ;
        RECT 467.885 404.220 478.000 431.760 ;
        RECT 90.700 403.700 478.000 404.220 ;
        RECT 91.695 391.655 116.305 403.700 ;
        RECT 118.295 391.655 142.905 403.700 ;
        RECT 144.895 391.655 169.505 403.700 ;
        RECT 171.495 391.655 196.105 403.700 ;
        RECT 198.095 391.655 222.705 403.700 ;
        RECT 224.695 391.655 249.305 403.700 ;
        RECT 251.295 391.655 275.905 403.700 ;
        RECT 277.895 391.655 302.505 403.700 ;
        RECT 304.495 391.655 329.105 403.700 ;
        RECT 331.095 391.655 355.705 403.700 ;
        RECT 357.695 391.655 382.305 403.700 ;
        RECT 384.295 391.655 408.905 403.700 ;
        RECT 410.895 391.655 435.505 403.700 ;
        RECT 437.495 391.655 462.105 403.700 ;
        RECT 91.695 376.160 116.305 388.205 ;
        RECT 118.295 376.160 142.905 388.205 ;
        RECT 144.895 376.160 169.505 388.205 ;
        RECT 171.495 376.160 196.105 388.205 ;
        RECT 198.095 376.160 222.705 388.205 ;
        RECT 224.695 376.160 249.305 388.205 ;
        RECT 251.295 376.160 275.905 388.205 ;
        RECT 277.895 376.160 302.505 388.205 ;
        RECT 304.495 376.160 329.105 388.205 ;
        RECT 331.095 376.160 355.705 388.205 ;
        RECT 357.695 376.160 382.305 388.205 ;
        RECT 384.295 376.160 408.905 388.205 ;
        RECT 410.895 376.160 435.505 388.205 ;
        RECT 437.495 376.160 462.105 388.205 ;
        RECT 467.885 376.160 478.000 403.700 ;
        RECT 90.700 375.640 478.000 376.160 ;
        RECT 91.695 363.595 116.305 375.640 ;
        RECT 118.295 363.595 142.905 375.640 ;
        RECT 144.895 363.595 169.505 375.640 ;
        RECT 171.495 363.595 196.105 375.640 ;
        RECT 198.095 363.595 222.705 375.640 ;
        RECT 224.695 363.595 249.305 375.640 ;
        RECT 251.295 363.595 275.905 375.640 ;
        RECT 277.895 363.595 302.505 375.640 ;
        RECT 304.495 363.595 329.105 375.640 ;
        RECT 331.095 363.595 355.705 375.640 ;
        RECT 357.695 363.595 382.305 375.640 ;
        RECT 384.295 363.595 408.905 375.640 ;
        RECT 410.895 363.595 435.505 375.640 ;
        RECT 437.495 363.595 462.105 375.640 ;
        RECT 91.695 348.100 116.305 360.145 ;
        RECT 118.295 348.100 142.905 360.145 ;
        RECT 144.895 348.100 169.505 360.145 ;
        RECT 171.495 348.100 196.105 360.145 ;
        RECT 198.095 348.100 222.705 360.145 ;
        RECT 224.695 348.100 249.305 360.145 ;
        RECT 251.295 348.100 275.905 360.145 ;
        RECT 277.895 348.100 302.505 360.145 ;
        RECT 304.495 348.100 329.105 360.145 ;
        RECT 331.095 348.100 355.705 360.145 ;
        RECT 357.695 348.100 382.305 360.145 ;
        RECT 384.295 348.100 408.905 360.145 ;
        RECT 410.895 348.100 435.505 360.145 ;
        RECT 437.495 348.100 462.105 360.145 ;
        RECT 467.885 348.100 478.000 375.640 ;
        RECT 90.700 347.580 478.000 348.100 ;
        RECT 91.695 335.535 116.305 347.580 ;
        RECT 118.295 335.535 142.905 347.580 ;
        RECT 144.895 335.535 169.505 347.580 ;
        RECT 171.495 335.535 196.105 347.580 ;
        RECT 198.095 335.535 222.705 347.580 ;
        RECT 224.695 335.535 249.305 347.580 ;
        RECT 251.295 335.535 275.905 347.580 ;
        RECT 277.895 335.535 302.505 347.580 ;
        RECT 304.495 335.535 329.105 347.580 ;
        RECT 331.095 335.535 355.705 347.580 ;
        RECT 357.695 335.535 382.305 347.580 ;
        RECT 384.295 335.535 408.905 347.580 ;
        RECT 410.895 335.535 435.505 347.580 ;
        RECT 437.495 335.535 462.105 347.580 ;
        RECT 91.695 320.040 116.305 332.085 ;
        RECT 118.295 320.040 142.905 332.085 ;
        RECT 144.895 320.040 169.505 332.085 ;
        RECT 171.495 320.040 196.105 332.085 ;
        RECT 198.095 320.040 222.705 332.085 ;
        RECT 224.695 320.040 249.305 332.085 ;
        RECT 251.295 320.040 275.905 332.085 ;
        RECT 277.895 320.040 302.505 332.085 ;
        RECT 304.495 320.040 329.105 332.085 ;
        RECT 331.095 320.040 355.705 332.085 ;
        RECT 357.695 320.040 382.305 332.085 ;
        RECT 384.295 320.040 408.905 332.085 ;
        RECT 410.895 320.040 435.505 332.085 ;
        RECT 437.495 320.040 462.105 332.085 ;
        RECT 467.885 320.040 478.000 347.580 ;
        RECT 90.700 319.520 478.000 320.040 ;
        RECT 91.695 307.475 116.305 319.520 ;
        RECT 118.295 307.475 142.905 319.520 ;
        RECT 144.895 307.475 169.505 319.520 ;
        RECT 171.495 307.475 196.105 319.520 ;
        RECT 198.095 307.475 222.705 319.520 ;
        RECT 224.695 307.475 249.305 319.520 ;
        RECT 251.295 307.475 275.905 319.520 ;
        RECT 277.895 307.475 302.505 319.520 ;
        RECT 304.495 307.475 329.105 319.520 ;
        RECT 331.095 307.475 355.705 319.520 ;
        RECT 357.695 307.475 382.305 319.520 ;
        RECT 384.295 307.475 408.905 319.520 ;
        RECT 410.895 307.475 435.505 319.520 ;
        RECT 437.495 307.475 462.105 319.520 ;
        RECT 91.695 291.980 116.305 304.025 ;
        RECT 118.295 291.980 142.905 304.025 ;
        RECT 144.895 291.980 169.505 304.025 ;
        RECT 171.495 291.980 196.105 304.025 ;
        RECT 198.095 291.980 222.705 304.025 ;
        RECT 224.695 291.980 249.305 304.025 ;
        RECT 251.295 291.980 275.905 304.025 ;
        RECT 277.895 291.980 302.505 304.025 ;
        RECT 304.495 291.980 329.105 304.025 ;
        RECT 331.095 291.980 355.705 304.025 ;
        RECT 357.695 291.980 382.305 304.025 ;
        RECT 384.295 291.980 408.905 304.025 ;
        RECT 410.895 291.980 435.505 304.025 ;
        RECT 437.495 291.980 462.105 304.025 ;
        RECT 467.885 291.980 478.000 319.520 ;
        RECT 90.700 291.460 478.000 291.980 ;
        RECT 91.695 279.415 116.305 291.460 ;
        RECT 118.295 279.415 142.905 291.460 ;
        RECT 144.895 279.415 169.505 291.460 ;
        RECT 171.495 279.415 196.105 291.460 ;
        RECT 198.095 279.415 222.705 291.460 ;
        RECT 224.695 279.415 249.305 291.460 ;
        RECT 251.295 279.415 275.905 291.460 ;
        RECT 277.895 279.415 302.505 291.460 ;
        RECT 304.495 279.415 329.105 291.460 ;
        RECT 331.095 279.415 355.705 291.460 ;
        RECT 357.695 279.415 382.305 291.460 ;
        RECT 384.295 279.415 408.905 291.460 ;
        RECT 410.895 279.415 435.505 291.460 ;
        RECT 437.495 279.415 462.105 291.460 ;
        RECT 91.695 263.920 116.305 275.965 ;
        RECT 118.295 263.920 142.905 275.965 ;
        RECT 144.895 263.920 169.505 275.965 ;
        RECT 171.495 263.920 196.105 275.965 ;
        RECT 198.095 263.920 222.705 275.965 ;
        RECT 224.695 263.920 249.305 275.965 ;
        RECT 251.295 263.920 275.905 275.965 ;
        RECT 277.895 263.920 302.505 275.965 ;
        RECT 304.495 263.920 329.105 275.965 ;
        RECT 331.095 263.920 355.705 275.965 ;
        RECT 357.695 263.920 382.305 275.965 ;
        RECT 384.295 263.920 408.905 275.965 ;
        RECT 410.895 263.920 435.505 275.965 ;
        RECT 437.495 263.920 462.105 275.965 ;
        RECT 467.885 263.920 478.000 291.460 ;
        RECT 90.700 263.400 478.000 263.920 ;
        RECT 91.695 251.355 116.305 263.400 ;
        RECT 118.295 251.355 142.905 263.400 ;
        RECT 144.895 251.355 169.505 263.400 ;
        RECT 171.495 251.355 196.105 263.400 ;
        RECT 198.095 251.355 222.705 263.400 ;
        RECT 224.695 251.355 249.305 263.400 ;
        RECT 251.295 251.355 275.905 263.400 ;
        RECT 277.895 251.355 302.505 263.400 ;
        RECT 304.495 251.355 329.105 263.400 ;
        RECT 331.095 251.355 355.705 263.400 ;
        RECT 357.695 251.355 382.305 263.400 ;
        RECT 384.295 251.355 408.905 263.400 ;
        RECT 410.895 251.355 435.505 263.400 ;
        RECT 437.495 251.355 462.105 263.400 ;
        RECT 91.695 235.860 116.305 247.905 ;
        RECT 118.295 235.860 142.905 247.905 ;
        RECT 144.895 235.860 169.505 247.905 ;
        RECT 171.495 235.860 196.105 247.905 ;
        RECT 198.095 235.860 222.705 247.905 ;
        RECT 224.695 235.860 249.305 247.905 ;
        RECT 251.295 235.860 275.905 247.905 ;
        RECT 277.895 235.860 302.505 247.905 ;
        RECT 304.495 235.860 329.105 247.905 ;
        RECT 331.095 235.860 355.705 247.905 ;
        RECT 357.695 235.860 382.305 247.905 ;
        RECT 384.295 235.860 408.905 247.905 ;
        RECT 410.895 235.860 435.505 247.905 ;
        RECT 437.495 235.860 462.105 247.905 ;
        RECT 467.885 235.860 478.000 263.400 ;
        RECT 90.700 235.340 478.000 235.860 ;
        RECT 91.695 223.295 116.305 235.340 ;
        RECT 118.295 223.295 142.905 235.340 ;
        RECT 144.895 223.295 169.505 235.340 ;
        RECT 171.495 223.295 196.105 235.340 ;
        RECT 198.095 223.295 222.705 235.340 ;
        RECT 224.695 223.295 249.305 235.340 ;
        RECT 251.295 223.295 275.905 235.340 ;
        RECT 277.895 223.295 302.505 235.340 ;
        RECT 304.495 223.295 329.105 235.340 ;
        RECT 331.095 223.295 355.705 235.340 ;
        RECT 357.695 223.295 382.305 235.340 ;
        RECT 384.295 223.295 408.905 235.340 ;
        RECT 410.895 223.295 435.505 235.340 ;
        RECT 437.495 223.295 462.105 235.340 ;
        RECT 91.695 207.800 116.305 219.845 ;
        RECT 118.295 207.800 142.905 219.845 ;
        RECT 144.895 207.800 169.505 219.845 ;
        RECT 171.495 207.800 196.105 219.845 ;
        RECT 198.095 207.800 222.705 219.845 ;
        RECT 224.695 207.800 249.305 219.845 ;
        RECT 251.295 207.800 275.905 219.845 ;
        RECT 277.895 207.800 302.505 219.845 ;
        RECT 304.495 207.800 329.105 219.845 ;
        RECT 331.095 207.800 355.705 219.845 ;
        RECT 357.695 207.800 382.305 219.845 ;
        RECT 384.295 207.800 408.905 219.845 ;
        RECT 410.895 207.800 435.505 219.845 ;
        RECT 437.495 207.800 462.105 219.845 ;
        RECT 467.885 207.800 478.000 235.340 ;
        RECT 90.700 207.280 478.000 207.800 ;
        RECT 91.695 195.235 116.305 207.280 ;
        RECT 118.295 195.235 142.905 207.280 ;
        RECT 144.895 195.235 169.505 207.280 ;
        RECT 171.495 195.235 196.105 207.280 ;
        RECT 198.095 195.235 222.705 207.280 ;
        RECT 224.695 195.235 249.305 207.280 ;
        RECT 251.295 195.235 275.905 207.280 ;
        RECT 277.895 195.235 302.505 207.280 ;
        RECT 304.495 195.235 329.105 207.280 ;
        RECT 331.095 195.235 355.705 207.280 ;
        RECT 357.695 195.235 382.305 207.280 ;
        RECT 384.295 195.235 408.905 207.280 ;
        RECT 410.895 195.235 435.505 207.280 ;
        RECT 437.495 195.235 462.105 207.280 ;
        RECT 91.695 179.740 116.305 191.785 ;
        RECT 118.295 179.740 142.905 191.785 ;
        RECT 144.895 179.740 169.505 191.785 ;
        RECT 171.495 179.740 196.105 191.785 ;
        RECT 198.095 179.740 222.705 191.785 ;
        RECT 224.695 179.740 249.305 191.785 ;
        RECT 251.295 179.740 275.905 191.785 ;
        RECT 277.895 179.740 302.505 191.785 ;
        RECT 304.495 179.740 329.105 191.785 ;
        RECT 331.095 179.740 355.705 191.785 ;
        RECT 357.695 179.740 382.305 191.785 ;
        RECT 384.295 179.740 408.905 191.785 ;
        RECT 410.895 179.740 435.505 191.785 ;
        RECT 437.495 179.740 462.105 191.785 ;
        RECT 467.885 179.740 478.000 207.280 ;
        RECT 90.700 179.220 478.000 179.740 ;
        RECT 91.695 167.175 116.305 179.220 ;
        RECT 118.295 167.175 142.905 179.220 ;
        RECT 144.895 167.175 169.505 179.220 ;
        RECT 171.495 167.175 196.105 179.220 ;
        RECT 198.095 167.175 222.705 179.220 ;
        RECT 224.695 167.175 249.305 179.220 ;
        RECT 251.295 167.175 275.905 179.220 ;
        RECT 277.895 167.175 302.505 179.220 ;
        RECT 304.495 167.175 329.105 179.220 ;
        RECT 331.095 167.175 355.705 179.220 ;
        RECT 357.695 167.175 382.305 179.220 ;
        RECT 384.295 167.175 408.905 179.220 ;
        RECT 410.895 167.175 435.505 179.220 ;
        RECT 437.495 167.175 462.105 179.220 ;
        RECT 91.695 151.680 116.305 163.725 ;
        RECT 118.295 151.680 142.905 163.725 ;
        RECT 144.895 151.680 169.505 163.725 ;
        RECT 171.495 151.680 196.105 163.725 ;
        RECT 198.095 151.680 222.705 163.725 ;
        RECT 224.695 151.680 249.305 163.725 ;
        RECT 251.295 151.680 275.905 163.725 ;
        RECT 277.895 151.680 302.505 163.725 ;
        RECT 304.495 151.680 329.105 163.725 ;
        RECT 331.095 151.680 355.705 163.725 ;
        RECT 357.695 151.680 382.305 163.725 ;
        RECT 384.295 151.680 408.905 163.725 ;
        RECT 410.895 151.680 435.505 163.725 ;
        RECT 437.495 151.680 462.105 163.725 ;
        RECT 467.885 151.680 478.000 179.220 ;
        RECT 90.700 151.160 478.000 151.680 ;
        RECT -0.970 137.895 0.485 144.570 ;
        RECT 1.980 137.895 11.590 142.440 ;
        RECT 13.580 137.895 23.190 142.440 ;
        RECT 25.180 137.895 34.790 142.440 ;
        RECT 36.780 137.895 46.390 142.440 ;
        RECT 48.380 137.895 57.990 142.440 ;
        RECT 59.980 137.895 69.590 142.440 ;
        RECT 71.580 137.895 81.190 142.440 ;
        RECT 91.695 139.115 116.305 151.160 ;
        RECT 118.295 139.115 142.905 151.160 ;
        RECT 144.895 139.115 169.505 151.160 ;
        RECT 171.495 139.115 196.105 151.160 ;
        RECT 198.095 139.115 222.705 151.160 ;
        RECT 224.695 139.115 249.305 151.160 ;
        RECT 251.295 139.115 275.905 151.160 ;
        RECT 277.895 139.115 302.505 151.160 ;
        RECT 304.495 139.115 329.105 151.160 ;
        RECT 331.095 139.115 355.705 151.160 ;
        RECT 357.695 139.115 382.305 151.160 ;
        RECT 384.295 139.115 408.905 151.160 ;
        RECT 410.895 139.115 435.505 151.160 ;
        RECT 437.495 139.115 462.105 151.160 ;
        RECT -0.970 137.375 82.185 137.895 ;
        RECT -0.970 124.835 0.485 137.375 ;
        RECT 1.980 132.830 11.590 137.375 ;
        RECT 13.580 132.830 23.190 137.375 ;
        RECT 25.180 132.830 34.790 137.375 ;
        RECT 36.780 132.830 46.390 137.375 ;
        RECT 48.380 132.830 57.990 137.375 ;
        RECT 59.980 132.830 69.590 137.375 ;
        RECT 71.580 132.830 81.190 137.375 ;
        RECT 1.980 124.835 11.590 129.380 ;
        RECT 13.580 124.835 23.190 129.380 ;
        RECT 25.180 124.835 34.790 129.380 ;
        RECT 36.780 124.835 46.390 129.380 ;
        RECT 48.380 124.835 57.990 129.380 ;
        RECT 59.980 124.835 69.590 129.380 ;
        RECT 71.580 124.835 81.190 129.380 ;
        RECT -0.970 124.315 82.185 124.835 ;
        RECT -0.970 111.775 0.485 124.315 ;
        RECT 1.980 119.770 11.590 124.315 ;
        RECT 13.580 119.770 23.190 124.315 ;
        RECT 25.180 119.770 34.790 124.315 ;
        RECT 36.780 119.770 46.390 124.315 ;
        RECT 48.380 119.770 57.990 124.315 ;
        RECT 59.980 119.770 69.590 124.315 ;
        RECT 71.580 119.770 81.190 124.315 ;
        RECT 91.695 123.620 116.305 135.665 ;
        RECT 118.295 123.620 142.905 135.665 ;
        RECT 144.895 123.620 169.505 135.665 ;
        RECT 171.495 123.620 196.105 135.665 ;
        RECT 198.095 123.620 222.705 135.665 ;
        RECT 224.695 123.620 249.305 135.665 ;
        RECT 251.295 123.620 275.905 135.665 ;
        RECT 277.895 123.620 302.505 135.665 ;
        RECT 304.495 123.620 329.105 135.665 ;
        RECT 331.095 123.620 355.705 135.665 ;
        RECT 357.695 123.620 382.305 135.665 ;
        RECT 384.295 123.620 408.905 135.665 ;
        RECT 410.895 123.620 435.505 135.665 ;
        RECT 437.495 123.620 462.105 135.665 ;
        RECT 467.885 123.620 478.000 151.160 ;
        RECT 90.700 123.100 478.000 123.620 ;
        RECT 1.980 111.775 11.590 116.320 ;
        RECT 13.580 111.775 23.190 116.320 ;
        RECT 25.180 111.775 34.790 116.320 ;
        RECT 36.780 111.775 46.390 116.320 ;
        RECT 48.380 111.775 57.990 116.320 ;
        RECT 59.980 111.775 69.590 116.320 ;
        RECT 71.580 111.775 81.190 116.320 ;
        RECT -0.970 111.255 82.185 111.775 ;
        RECT -0.970 98.715 0.485 111.255 ;
        RECT 1.980 106.710 11.590 111.255 ;
        RECT 13.580 106.710 23.190 111.255 ;
        RECT 25.180 106.710 34.790 111.255 ;
        RECT 36.780 106.710 46.390 111.255 ;
        RECT 48.380 106.710 57.990 111.255 ;
        RECT 59.980 106.710 69.590 111.255 ;
        RECT 71.580 106.710 81.190 111.255 ;
        RECT 91.695 111.055 116.305 123.100 ;
        RECT 118.295 111.055 142.905 123.100 ;
        RECT 144.895 111.055 169.505 123.100 ;
        RECT 171.495 111.055 196.105 123.100 ;
        RECT 198.095 111.055 222.705 123.100 ;
        RECT 224.695 111.055 249.305 123.100 ;
        RECT 251.295 111.055 275.905 123.100 ;
        RECT 277.895 111.055 302.505 123.100 ;
        RECT 304.495 111.055 329.105 123.100 ;
        RECT 331.095 111.055 355.705 123.100 ;
        RECT 357.695 111.055 382.305 123.100 ;
        RECT 384.295 111.055 408.905 123.100 ;
        RECT 410.895 111.055 435.505 123.100 ;
        RECT 437.495 111.055 462.105 123.100 ;
        RECT 1.980 98.715 11.590 103.260 ;
        RECT 13.580 98.715 23.190 103.260 ;
        RECT 25.180 98.715 34.790 103.260 ;
        RECT 36.780 98.715 46.390 103.260 ;
        RECT 48.380 98.715 57.990 103.260 ;
        RECT 59.980 98.715 69.590 103.260 ;
        RECT 71.580 98.715 81.190 103.260 ;
        RECT -0.970 98.195 82.185 98.715 ;
        RECT -0.970 85.655 0.485 98.195 ;
        RECT 1.980 93.650 11.590 98.195 ;
        RECT 13.580 93.650 23.190 98.195 ;
        RECT 25.180 93.650 34.790 98.195 ;
        RECT 36.780 93.650 46.390 98.195 ;
        RECT 48.380 93.650 57.990 98.195 ;
        RECT 59.980 93.650 69.590 98.195 ;
        RECT 71.580 93.650 81.190 98.195 ;
        RECT 91.695 95.560 116.305 107.605 ;
        RECT 118.295 95.560 142.905 107.605 ;
        RECT 144.895 95.560 169.505 107.605 ;
        RECT 171.495 95.560 196.105 107.605 ;
        RECT 198.095 95.560 222.705 107.605 ;
        RECT 224.695 95.560 249.305 107.605 ;
        RECT 251.295 95.560 275.905 107.605 ;
        RECT 277.895 95.560 302.505 107.605 ;
        RECT 304.495 95.560 329.105 107.605 ;
        RECT 331.095 95.560 355.705 107.605 ;
        RECT 357.695 95.560 382.305 107.605 ;
        RECT 384.295 95.560 408.905 107.605 ;
        RECT 410.895 95.560 435.505 107.605 ;
        RECT 437.495 95.560 462.105 107.605 ;
        RECT 467.885 95.560 478.000 123.100 ;
        RECT 90.700 95.040 478.000 95.560 ;
        RECT 1.980 85.655 11.590 90.200 ;
        RECT 13.580 85.655 23.190 90.200 ;
        RECT 25.180 85.655 34.790 90.200 ;
        RECT 36.780 85.655 46.390 90.200 ;
        RECT 48.380 85.655 57.990 90.200 ;
        RECT 59.980 85.655 69.590 90.200 ;
        RECT 71.580 85.655 81.190 90.200 ;
        RECT -0.970 85.135 82.185 85.655 ;
        RECT -0.970 72.595 0.485 85.135 ;
        RECT 1.980 80.590 11.590 85.135 ;
        RECT 13.580 80.590 23.190 85.135 ;
        RECT 25.180 80.590 34.790 85.135 ;
        RECT 36.780 80.590 46.390 85.135 ;
        RECT 48.380 80.590 57.990 85.135 ;
        RECT 59.980 80.590 69.590 85.135 ;
        RECT 71.580 80.590 81.190 85.135 ;
        RECT 91.695 82.995 116.305 95.040 ;
        RECT 118.295 82.995 142.905 95.040 ;
        RECT 144.895 82.995 169.505 95.040 ;
        RECT 171.495 82.995 196.105 95.040 ;
        RECT 198.095 82.995 222.705 95.040 ;
        RECT 224.695 82.995 249.305 95.040 ;
        RECT 251.295 82.995 275.905 95.040 ;
        RECT 277.895 82.995 302.505 95.040 ;
        RECT 304.495 82.995 329.105 95.040 ;
        RECT 331.095 82.995 355.705 95.040 ;
        RECT 357.695 82.995 382.305 95.040 ;
        RECT 384.295 82.995 408.905 95.040 ;
        RECT 410.895 82.995 435.505 95.040 ;
        RECT 437.495 82.995 462.105 95.040 ;
        RECT 1.980 72.595 11.590 77.140 ;
        RECT 13.580 72.595 23.190 77.140 ;
        RECT 25.180 72.595 34.790 77.140 ;
        RECT 36.780 72.595 46.390 77.140 ;
        RECT 48.380 72.595 57.990 77.140 ;
        RECT 59.980 72.595 69.590 77.140 ;
        RECT 71.580 72.595 81.190 77.140 ;
        RECT -0.970 72.075 82.185 72.595 ;
        RECT -0.970 59.535 0.485 72.075 ;
        RECT 1.980 67.530 11.590 72.075 ;
        RECT 13.580 67.530 23.190 72.075 ;
        RECT 25.180 67.530 34.790 72.075 ;
        RECT 36.780 67.530 46.390 72.075 ;
        RECT 48.380 67.530 57.990 72.075 ;
        RECT 59.980 67.530 69.590 72.075 ;
        RECT 71.580 67.530 81.190 72.075 ;
        RECT 91.695 67.500 116.305 79.545 ;
        RECT 118.295 67.500 142.905 79.545 ;
        RECT 144.895 67.500 169.505 79.545 ;
        RECT 171.495 67.500 196.105 79.545 ;
        RECT 198.095 67.500 222.705 79.545 ;
        RECT 224.695 67.500 249.305 79.545 ;
        RECT 251.295 67.500 275.905 79.545 ;
        RECT 277.895 67.500 302.505 79.545 ;
        RECT 304.495 67.500 329.105 79.545 ;
        RECT 331.095 67.500 355.705 79.545 ;
        RECT 357.695 67.500 382.305 79.545 ;
        RECT 384.295 67.500 408.905 79.545 ;
        RECT 410.895 67.500 435.505 79.545 ;
        RECT 437.495 67.500 462.105 79.545 ;
        RECT 467.885 67.500 478.000 95.040 ;
        RECT 90.700 66.980 478.000 67.500 ;
        RECT 1.980 59.535 11.590 64.080 ;
        RECT 13.580 59.535 23.190 64.080 ;
        RECT 25.180 59.535 34.790 64.080 ;
        RECT 36.780 59.535 46.390 64.080 ;
        RECT 48.380 59.535 57.990 64.080 ;
        RECT 59.980 59.535 69.590 64.080 ;
        RECT 71.580 59.535 81.190 64.080 ;
        RECT -0.970 59.015 82.185 59.535 ;
        RECT -0.970 54.325 0.485 59.015 ;
        RECT 1.980 54.470 11.590 59.015 ;
        RECT 13.580 54.470 23.190 59.015 ;
        RECT 25.180 54.470 34.790 59.015 ;
        RECT 36.780 54.470 46.390 59.015 ;
        RECT 48.380 54.470 57.990 59.015 ;
        RECT 59.980 54.470 69.590 59.015 ;
        RECT 71.580 54.470 81.190 59.015 ;
        RECT 91.695 54.935 116.305 66.980 ;
        RECT 118.295 54.935 142.905 66.980 ;
        RECT 144.895 54.935 169.505 66.980 ;
        RECT 171.495 54.935 196.105 66.980 ;
        RECT 198.095 54.935 222.705 66.980 ;
        RECT 224.695 54.935 249.305 66.980 ;
        RECT 251.295 54.935 275.905 66.980 ;
        RECT 277.895 54.935 302.505 66.980 ;
        RECT 304.495 54.935 329.105 66.980 ;
        RECT 331.095 54.935 355.705 66.980 ;
        RECT 357.695 54.935 382.305 66.980 ;
        RECT 384.295 54.935 408.905 66.980 ;
        RECT 410.895 54.935 435.505 66.980 ;
        RECT 437.495 54.935 462.105 66.980 ;
        RECT 467.885 53.885 478.000 66.980 ;
  END
END sky130_aa_ip__programmable_pll
END LIBRARY

