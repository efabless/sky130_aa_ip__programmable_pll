magic
tech sky130A
magscale 1 2
timestamp 1717691374
<< nwell >>
rect 1075 -1053 14393 -1041
rect 1075 -1057 5170 -1053
rect 1075 -1516 3578 -1057
rect 3586 -1076 5170 -1057
rect 5181 -1058 14393 -1053
rect 5181 -1067 5189 -1058
rect 4497 -1429 5170 -1076
rect 6104 -1427 6792 -1058
rect 7662 -1084 8753 -1058
rect 7353 -1163 8753 -1084
rect 7662 -1514 8753 -1163
<< locali >>
rect -361 1212 14601 1405
rect -316 1157 736 1212
rect 2866 1143 3459 1212
rect 5279 1155 5872 1212
rect 7118 757 7152 758
rect 1338 723 1830 757
rect 4543 723 4736 757
rect 6985 723 7152 757
rect 1796 356 1830 723
rect 4702 357 4736 723
rect 4701 356 4736 357
rect 7118 356 7152 723
rect 1790 344 1836 356
rect 1790 310 1796 344
rect 1830 310 1836 344
rect 1790 266 1836 310
rect 1790 232 1796 266
rect 1830 232 1836 266
rect 1790 220 1836 232
rect 4695 344 4741 356
rect 4695 310 4701 344
rect 4735 310 4741 344
rect 4695 266 4741 310
rect 4695 232 4701 266
rect 4735 232 4741 266
rect 4695 220 4741 232
rect 7112 344 7158 356
rect 7112 310 7118 344
rect 7152 310 7158 344
rect 7244 340 7359 1212
rect 7813 1143 8406 1212
rect 9493 723 9632 757
rect 9598 356 9632 723
rect 9592 344 9638 356
rect 7112 266 7158 310
rect 7112 232 7118 266
rect 7152 232 7158 266
rect 7112 220 7158 232
rect 7241 328 7364 340
rect 7241 294 7247 328
rect 7281 294 7324 328
rect 7358 294 7364 328
rect 7241 250 7364 294
rect 7241 216 7247 250
rect 7281 216 7324 250
rect 7358 216 7364 250
rect 9592 310 9598 344
rect 9632 310 9638 344
rect 9727 340 9841 1212
rect 10329 1136 10922 1212
rect 12058 723 12180 757
rect 12146 360 12180 723
rect 12294 375 12409 1212
rect 12684 1126 13736 1212
rect 14526 723 14623 757
rect 12291 363 12414 375
rect 12140 348 12186 360
rect 9592 266 9638 310
rect 9592 232 9598 266
rect 9632 232 9638 266
rect 9592 220 9638 232
rect 9724 328 9847 340
rect 9724 294 9730 328
rect 9764 294 9807 328
rect 9841 294 9847 328
rect 9724 250 9847 294
rect 7241 204 7364 216
rect 9724 216 9730 250
rect 9764 216 9807 250
rect 9841 216 9847 250
rect 12140 314 12146 348
rect 12180 314 12186 348
rect 12140 270 12186 314
rect 12140 236 12146 270
rect 12180 236 12186 270
rect 12291 329 12297 363
rect 12331 329 12374 363
rect 12408 329 12414 363
rect 12291 285 12414 329
rect 12291 251 12297 285
rect 12331 251 12374 285
rect 12408 251 12414 285
rect 12291 239 12414 251
rect 12140 224 12186 236
rect 9724 204 9847 216
rect -737 1 331 128
rect 1338 23 3121 76
rect 4419 23 5260 76
rect 6900 23 7814 76
rect 9419 23 10376 76
rect 11980 24 12804 111
rect -737 -2682 -476 1
rect 9337 -22 9473 -16
rect 6840 -32 6976 -29
rect 4838 -35 7009 -32
rect 4838 -66 6852 -35
rect 1752 -82 1888 -76
rect 1616 -116 1764 -82
rect 1798 -116 1842 -82
rect 1876 -116 1888 -82
rect 4657 -98 4793 -92
rect 4657 -101 4669 -98
rect 604 -1062 727 -1050
rect 604 -1096 610 -1062
rect 644 -1096 687 -1062
rect 721 -1096 727 -1062
rect 604 -1140 727 -1096
rect 604 -1174 610 -1140
rect 644 -1174 687 -1140
rect 721 -1174 727 -1140
rect 604 -1186 727 -1174
rect 1616 -1659 1650 -116
rect 1752 -122 1888 -116
rect 1992 -132 4669 -101
rect 4703 -132 4747 -98
rect 4781 -132 4793 -98
rect 1992 -135 4793 -132
rect 1992 -174 2026 -135
rect 4657 -138 4793 -135
rect 1686 -208 2026 -174
rect 4838 -190 4872 -66
rect 6840 -69 6852 -66
rect 6886 -69 6930 -35
rect 6964 -66 7009 -35
rect 9337 -56 9349 -22
rect 9383 -56 9427 -22
rect 9461 -56 9473 -22
rect 9337 -62 9473 -56
rect 6964 -69 6976 -66
rect 6840 -75 6976 -69
rect 9337 -110 9386 -62
rect 1686 -1577 1720 -208
rect 3370 -224 4872 -190
rect 4934 -146 9386 -110
rect 1820 -1061 1943 -1049
rect 1820 -1095 1826 -1061
rect 1860 -1095 1903 -1061
rect 1937 -1095 1943 -1061
rect 3176 -1056 3299 -1044
rect 3176 -1077 3182 -1056
rect 1820 -1139 1943 -1095
rect 1820 -1173 1826 -1139
rect 1860 -1173 1903 -1139
rect 1937 -1173 1943 -1139
rect 2403 -1090 3182 -1077
rect 3216 -1090 3259 -1056
rect 3293 -1090 3299 -1056
rect 2403 -1134 3299 -1090
rect 2403 -1150 3182 -1134
rect 1820 -1185 1943 -1173
rect 3176 -1168 3182 -1150
rect 3216 -1168 3259 -1134
rect 3293 -1168 3299 -1134
rect 3176 -1180 3299 -1168
rect 1776 -1500 1912 -1494
rect 1776 -1534 1788 -1500
rect 1822 -1534 1866 -1500
rect 1900 -1534 1912 -1500
rect 1776 -1540 1912 -1534
rect 1686 -1615 1795 -1577
rect 1616 -1693 1821 -1659
rect 3370 -1717 3410 -224
rect 4934 -258 4970 -146
rect 7242 -214 7365 -213
rect 3449 -294 4970 -258
rect 7059 -230 7365 -214
rect 7059 -264 7065 -230
rect 7099 -264 7142 -230
rect 7176 -264 7248 -230
rect 7282 -264 7325 -230
rect 7359 -264 7365 -230
rect 7059 -276 7365 -264
rect 9725 -260 9848 -248
rect 3449 -1621 3485 -294
rect 4998 -739 5134 -733
rect 4998 -773 5010 -739
rect 5044 -773 5088 -739
rect 5122 -773 5134 -739
rect 4998 -779 5134 -773
rect 3577 -1058 3700 -1046
rect 3577 -1092 3583 -1058
rect 3617 -1092 3660 -1058
rect 3694 -1092 3700 -1058
rect 3577 -1136 3700 -1092
rect 3577 -1170 3583 -1136
rect 3617 -1170 3660 -1136
rect 3694 -1170 3700 -1136
rect 3577 -1182 3700 -1170
rect 4805 -1081 4928 -1069
rect 4805 -1115 4811 -1081
rect 4845 -1115 4888 -1081
rect 4922 -1115 4928 -1081
rect 4805 -1159 4928 -1115
rect 4805 -1193 4811 -1159
rect 4845 -1193 4888 -1159
rect 4922 -1193 4928 -1159
rect 4805 -1205 4928 -1193
rect 3449 -1659 3541 -1621
rect 3469 -1661 3541 -1659
rect 3370 -1757 3530 -1717
rect 3081 -1897 3331 -1839
rect -278 -2682 -81 -2175
rect 225 -2682 422 -2190
rect 738 -2682 935 -2180
rect 1271 -2682 1468 -2195
rect 3266 -2352 3331 -1897
rect 1886 -2682 2032 -2356
rect 3265 -2358 3401 -2352
rect 2246 -2682 2392 -2364
rect 2512 -2682 2658 -2361
rect 2957 -2682 3103 -2359
rect 3265 -2392 3277 -2358
rect 3311 -2392 3355 -2358
rect 3389 -2392 3401 -2358
rect 3265 -2398 3401 -2392
rect 3592 -2682 3743 -2191
rect 3885 -2682 4036 -2186
rect 4327 -2682 4478 -2159
rect 4833 -2240 4903 -1435
rect 4998 -1715 5038 -779
rect 5083 -823 5238 -817
rect 5083 -857 5095 -823
rect 5129 -857 5173 -823
rect 5207 -857 5238 -823
rect 5083 -863 5238 -857
rect 5083 -1613 5119 -863
rect 5194 -1082 5317 -1070
rect 5194 -1116 5200 -1082
rect 5234 -1116 5277 -1082
rect 5311 -1084 5317 -1082
rect 7245 -1084 7360 -276
rect 9725 -294 9731 -260
rect 9765 -294 9808 -260
rect 9842 -294 9848 -260
rect 9725 -338 9848 -294
rect 9725 -372 9731 -338
rect 9765 -372 9808 -338
rect 9842 -372 9848 -338
rect 9725 -384 9848 -372
rect 12140 -358 12186 -346
rect 8293 -910 8430 -903
rect 8293 -944 8305 -910
rect 8339 -944 8383 -910
rect 8417 -944 8430 -910
rect 8293 -954 8430 -944
rect 8172 -1069 8295 -1057
rect 8172 -1084 8178 -1069
rect 5311 -1103 8178 -1084
rect 8212 -1103 8255 -1069
rect 8289 -1103 8295 -1069
rect 5311 -1116 8295 -1103
rect 5194 -1147 8295 -1116
rect 5194 -1160 8178 -1147
rect 5194 -1194 5200 -1160
rect 5234 -1194 5277 -1160
rect 5311 -1163 8178 -1160
rect 5311 -1194 5317 -1163
rect 8172 -1181 8178 -1163
rect 8212 -1181 8255 -1147
rect 8289 -1181 8295 -1147
rect 8172 -1193 8295 -1181
rect 5194 -1206 5317 -1194
rect 6681 -1423 6727 -1411
rect 5083 -1657 5174 -1613
rect 5096 -1661 5174 -1657
rect 6441 -1668 6475 -1440
rect 6681 -1457 6687 -1423
rect 6721 -1457 6727 -1423
rect 6681 -1495 6727 -1457
rect 6681 -1501 6759 -1495
rect 6681 -1535 6687 -1501
rect 6721 -1535 6759 -1501
rect 6681 -1549 6759 -1535
rect 6510 -1586 6646 -1585
rect 6510 -1591 6782 -1586
rect 6510 -1625 6522 -1591
rect 6556 -1625 6600 -1591
rect 6634 -1624 6782 -1591
rect 6634 -1625 6646 -1624
rect 6510 -1631 6646 -1625
rect 8043 -1666 8228 -1658
rect 6441 -1702 6761 -1668
rect 8043 -1700 8099 -1666
rect 8133 -1700 8177 -1666
rect 8211 -1700 8228 -1666
rect 8043 -1711 8228 -1700
rect 8391 -1708 8430 -954
rect 8466 -1070 8589 -1058
rect 8466 -1104 8472 -1070
rect 8506 -1104 8549 -1070
rect 8583 -1104 8589 -1070
rect 8466 -1148 8589 -1104
rect 9729 -1110 9844 -384
rect 12140 -392 12146 -358
rect 12180 -392 12186 -358
rect 12140 -436 12186 -392
rect 12140 -470 12146 -436
rect 12180 -470 12186 -436
rect 12140 -482 12186 -470
rect 12292 -404 12415 -392
rect 12292 -438 12298 -404
rect 12332 -438 12375 -404
rect 12409 -438 12415 -404
rect 12292 -482 12415 -438
rect 12143 -735 12183 -482
rect 12292 -516 12298 -482
rect 12332 -516 12375 -482
rect 12409 -516 12415 -482
rect 12292 -528 12415 -516
rect 12047 -741 12183 -735
rect 12047 -775 12059 -741
rect 12093 -775 12137 -741
rect 12171 -775 12183 -741
rect 12047 -781 12183 -775
rect 12295 -1127 12410 -528
rect 14589 -808 14623 723
rect 14527 -814 14663 -808
rect 14527 -848 14539 -814
rect 14573 -848 14617 -814
rect 14651 -848 14663 -814
rect 14527 -854 14663 -848
rect 8466 -1182 8472 -1148
rect 8506 -1182 8549 -1148
rect 8583 -1182 8589 -1148
rect 8466 -1194 8589 -1182
rect 4998 -1755 5138 -1715
rect 8966 -2074 9122 -2073
rect 4833 -2246 4969 -2240
rect 4833 -2280 4845 -2246
rect 4879 -2280 4923 -2246
rect 4957 -2280 4969 -2246
rect 4833 -2286 4969 -2280
rect 5252 -2682 5376 -2181
rect 5582 -2682 5706 -2166
rect 5932 -2682 6083 -2157
rect 6877 -2682 7007 -2354
rect 7323 -2682 7453 -2378
rect 7640 -2682 7770 -2368
rect 7946 -2682 8076 -2368
rect 8824 -2682 9122 -2074
rect -737 -2943 9122 -2682
<< viali >>
rect 1796 310 1830 344
rect 1796 232 1830 266
rect 4701 310 4735 344
rect 4701 232 4735 266
rect 7118 310 7152 344
rect 7118 232 7152 266
rect 7247 294 7281 328
rect 7324 294 7358 328
rect 7247 216 7281 250
rect 7324 216 7358 250
rect 9598 310 9632 344
rect 9598 232 9632 266
rect 9730 294 9764 328
rect 9807 294 9841 328
rect 9730 216 9764 250
rect 9807 216 9841 250
rect 12146 314 12180 348
rect 12146 236 12180 270
rect 12297 329 12331 363
rect 12374 329 12408 363
rect 12297 251 12331 285
rect 12374 251 12408 285
rect 1764 -116 1798 -82
rect 1842 -116 1876 -82
rect 610 -1096 644 -1062
rect 687 -1096 721 -1062
rect 610 -1174 644 -1140
rect 687 -1174 721 -1140
rect 4669 -132 4703 -98
rect 4747 -132 4781 -98
rect 6852 -69 6886 -35
rect 6930 -69 6964 -35
rect 9349 -56 9383 -22
rect 9427 -56 9461 -22
rect 1826 -1095 1860 -1061
rect 1903 -1095 1937 -1061
rect 1826 -1173 1860 -1139
rect 1903 -1173 1937 -1139
rect 3182 -1090 3216 -1056
rect 3259 -1090 3293 -1056
rect 3182 -1168 3216 -1134
rect 3259 -1168 3293 -1134
rect 1788 -1534 1822 -1500
rect 1866 -1534 1900 -1500
rect 7065 -264 7099 -230
rect 7142 -264 7176 -230
rect 7248 -264 7282 -230
rect 7325 -264 7359 -230
rect 5010 -773 5044 -739
rect 5088 -773 5122 -739
rect 3583 -1092 3617 -1058
rect 3660 -1092 3694 -1058
rect 3583 -1170 3617 -1136
rect 3660 -1170 3694 -1136
rect 4811 -1115 4845 -1081
rect 4888 -1115 4922 -1081
rect 4811 -1193 4845 -1159
rect 4888 -1193 4922 -1159
rect 3277 -2392 3311 -2358
rect 3355 -2392 3389 -2358
rect 5095 -857 5129 -823
rect 5173 -857 5207 -823
rect 5200 -1116 5234 -1082
rect 5277 -1116 5311 -1082
rect 9731 -294 9765 -260
rect 9808 -294 9842 -260
rect 9731 -372 9765 -338
rect 9808 -372 9842 -338
rect 8305 -944 8339 -910
rect 8383 -944 8417 -910
rect 8178 -1103 8212 -1069
rect 8255 -1103 8289 -1069
rect 5200 -1194 5234 -1160
rect 5277 -1194 5311 -1160
rect 8178 -1181 8212 -1147
rect 8255 -1181 8289 -1147
rect 6687 -1457 6721 -1423
rect 6687 -1535 6721 -1501
rect 6522 -1625 6556 -1591
rect 6600 -1625 6634 -1591
rect 8099 -1700 8133 -1666
rect 8177 -1700 8211 -1666
rect 8472 -1104 8506 -1070
rect 8549 -1104 8583 -1070
rect 12146 -392 12180 -358
rect 12146 -470 12180 -436
rect 12298 -438 12332 -404
rect 12375 -438 12409 -404
rect 12298 -516 12332 -482
rect 12375 -516 12409 -482
rect 12059 -775 12093 -741
rect 12137 -775 12171 -741
rect 14539 -848 14573 -814
rect 14617 -848 14651 -814
rect 8472 -1182 8506 -1148
rect 8549 -1182 8583 -1148
rect 4845 -2280 4879 -2246
rect 4923 -2280 4957 -2246
<< metal1 >>
rect -619 641 -445 669
rect -6 641 63 669
rect 1627 641 2656 669
rect 4932 641 5065 669
rect 7407 641 7546 669
rect 9879 641 10028 669
rect 12450 641 12547 669
rect -619 504 -365 532
rect -6 504 155 532
rect 1627 -34 1655 641
rect -1330 -62 1655 -34
rect 1694 504 2753 532
rect 1694 -94 1722 504
rect 1790 344 1836 356
rect 1790 310 1796 344
rect 1830 310 1836 344
rect 1790 266 1836 310
rect 1790 232 1796 266
rect 1830 232 1836 266
rect 1790 220 1836 232
rect 4695 344 4741 356
rect 4695 310 4701 344
rect 4735 310 4741 344
rect 4695 266 4741 310
rect 4695 232 4701 266
rect 4735 232 4741 266
rect 4695 220 4741 232
rect 1791 -76 1835 220
rect -1330 -122 1722 -94
rect 1752 -82 1888 -76
rect 1752 -116 1764 -82
rect 1798 -116 1842 -82
rect 1876 -116 1888 -82
rect 4696 -92 4740 220
rect 1752 -122 1888 -116
rect 4657 -98 4793 -92
rect 4657 -132 4669 -98
rect 4703 -132 4747 -98
rect 4781 -132 4793 -98
rect 4657 -138 4793 -132
rect 4932 -167 4960 641
rect -1333 -195 4960 -167
rect -738 -205 4960 -195
rect 5015 504 5136 532
rect 5015 -241 5043 504
rect 7112 344 7158 356
rect 7112 310 7118 344
rect 7152 310 7158 344
rect 7112 266 7158 310
rect 7112 232 7118 266
rect 7152 232 7158 266
rect 7112 220 7158 232
rect 7241 328 7364 340
rect 7241 294 7247 328
rect 7281 294 7324 328
rect 7358 294 7364 328
rect 7241 250 7364 294
rect 6840 -30 6976 -29
rect 7113 -30 7157 220
rect 7241 216 7247 250
rect 7281 216 7324 250
rect 7358 216 7364 250
rect 7241 204 7364 216
rect 6840 -35 7157 -30
rect 6840 -69 6852 -35
rect 6886 -69 6930 -35
rect 6964 -69 7157 -35
rect 6840 -74 7157 -69
rect 6840 -75 6976 -74
rect 7246 -213 7360 204
rect 7242 -214 7365 -213
rect -1330 -269 5043 -241
rect 7059 -230 7365 -214
rect 7059 -264 7065 -230
rect 7099 -264 7142 -230
rect 7176 -264 7248 -230
rect 7282 -264 7325 -230
rect 7359 -264 7365 -230
rect 7059 -276 7365 -264
rect 7407 -304 7435 641
rect -1330 -332 7435 -304
rect 7481 504 7616 532
rect 7481 -361 7509 504
rect 9592 344 9638 356
rect 9592 310 9598 344
rect 9632 310 9638 344
rect 9592 266 9638 310
rect 9592 232 9598 266
rect 9632 232 9638 266
rect 9592 220 9638 232
rect 9724 328 9847 340
rect 9724 294 9730 328
rect 9764 294 9807 328
rect 9841 294 9847 328
rect 9724 250 9847 294
rect 9337 -17 9473 -16
rect 9593 -17 9637 220
rect 9724 216 9730 250
rect 9764 216 9807 250
rect 9841 216 9847 250
rect 9724 204 9847 216
rect 9337 -22 9638 -17
rect 9337 -56 9349 -22
rect 9383 -56 9427 -22
rect 9461 -56 9638 -22
rect 9337 -61 9638 -56
rect 9337 -62 9473 -61
rect 9729 -248 9843 204
rect -1330 -389 7509 -361
rect 9725 -260 9848 -248
rect 9725 -294 9731 -260
rect 9765 -294 9808 -260
rect 9842 -294 9848 -260
rect 9725 -338 9848 -294
rect 9725 -372 9731 -338
rect 9765 -372 9808 -338
rect 9842 -372 9848 -338
rect 9725 -384 9848 -372
rect 9879 -417 9907 641
rect -1330 -468 9907 -417
rect 9965 504 10137 532
rect 9965 -500 9993 504
rect 12291 363 12414 375
rect 12140 348 12186 360
rect 12140 314 12146 348
rect 12180 314 12186 348
rect 12140 270 12186 314
rect 12140 236 12146 270
rect 12180 236 12186 270
rect 12291 329 12297 363
rect 12331 329 12374 363
rect 12408 329 12414 363
rect 12291 285 12414 329
rect 12291 251 12297 285
rect 12331 251 12374 285
rect 12408 251 12414 285
rect 12291 239 12414 251
rect 12140 224 12186 236
rect 12141 -346 12185 224
rect 12140 -358 12186 -346
rect 12140 -392 12146 -358
rect 12180 -392 12186 -358
rect 12296 -392 12410 239
rect 12140 -436 12186 -392
rect 12140 -470 12146 -436
rect 12180 -470 12186 -436
rect 12140 -482 12186 -470
rect 12292 -404 12415 -392
rect 12292 -438 12298 -404
rect 12332 -438 12375 -404
rect 12409 -438 12415 -404
rect 12292 -482 12415 -438
rect -1330 -536 9993 -500
rect 12292 -516 12298 -482
rect 12332 -516 12375 -482
rect 12409 -516 12415 -482
rect 12292 -528 12415 -516
rect 12450 -567 12478 641
rect -1330 -618 12478 -567
rect 12522 504 12634 532
rect 12522 -646 12550 504
rect -1330 -697 12550 -646
rect 4998 -737 5134 -733
rect 12047 -737 12183 -735
rect 4998 -739 12183 -737
rect 4998 -773 5010 -739
rect 5044 -773 5088 -739
rect 5122 -741 12183 -739
rect 5122 -773 12059 -741
rect 4998 -775 12059 -773
rect 12093 -775 12137 -741
rect 12171 -775 12183 -741
rect 4998 -779 12183 -775
rect 12047 -781 12183 -779
rect 14527 -814 14663 -808
rect 5083 -819 5238 -817
rect 14527 -819 14539 -814
rect 5083 -823 14539 -819
rect 5083 -857 5095 -823
rect 5129 -857 5173 -823
rect 5207 -848 14539 -823
rect 14573 -848 14617 -814
rect 14651 -848 14663 -814
rect 5207 -854 14663 -848
rect 5207 -857 14539 -854
rect 5083 -861 14539 -857
rect 5083 -863 5238 -861
rect -1330 -910 8430 -903
rect -1330 -944 8305 -910
rect 8339 -944 8383 -910
rect 8417 -944 8430 -910
rect -1330 -954 8430 -944
rect 604 -1062 727 -1050
rect 1820 -1061 1943 -1049
rect 1820 -1062 1826 -1061
rect 604 -1096 610 -1062
rect 644 -1096 687 -1062
rect 721 -1095 1826 -1062
rect 1860 -1095 1903 -1061
rect 1937 -1095 1943 -1061
rect 721 -1096 1943 -1095
rect 604 -1139 1943 -1096
rect 604 -1140 1826 -1139
rect 604 -1174 610 -1140
rect 644 -1174 687 -1140
rect 721 -1167 1826 -1140
rect 721 -1174 727 -1167
rect 604 -1186 727 -1174
rect 1820 -1173 1826 -1167
rect 1860 -1173 1903 -1139
rect 1937 -1173 1943 -1139
rect 1820 -1185 1943 -1173
rect 3176 -1055 3299 -1044
rect 3577 -1055 3700 -1046
rect 3176 -1056 3700 -1055
rect 3176 -1090 3182 -1056
rect 3216 -1090 3259 -1056
rect 3293 -1058 3700 -1056
rect 3293 -1090 3583 -1058
rect 3176 -1092 3583 -1090
rect 3617 -1092 3660 -1058
rect 3694 -1092 3700 -1058
rect 8172 -1069 8295 -1057
rect 3176 -1134 3700 -1092
rect 3176 -1168 3182 -1134
rect 3216 -1168 3259 -1134
rect 3293 -1136 3700 -1134
rect 3293 -1162 3583 -1136
rect 3293 -1168 3299 -1162
rect 3176 -1180 3299 -1168
rect 3577 -1170 3583 -1162
rect 3617 -1170 3660 -1136
rect 3694 -1170 3700 -1136
rect 3577 -1182 3700 -1170
rect 4805 -1081 4928 -1069
rect 4805 -1115 4811 -1081
rect 4845 -1115 4888 -1081
rect 4922 -1085 4928 -1081
rect 5194 -1082 5317 -1070
rect 5194 -1085 5200 -1082
rect 4922 -1115 5200 -1085
rect 4805 -1116 5200 -1115
rect 5234 -1116 5277 -1082
rect 5311 -1116 5317 -1082
rect 4805 -1159 5317 -1116
rect 4805 -1193 4811 -1159
rect 4845 -1193 4888 -1159
rect 4922 -1160 5317 -1159
rect 4922 -1192 5200 -1160
rect 4922 -1193 4928 -1192
rect 4805 -1205 4928 -1193
rect 5194 -1194 5200 -1192
rect 5234 -1194 5277 -1160
rect 5311 -1194 5317 -1160
rect 8172 -1103 8178 -1069
rect 8212 -1103 8255 -1069
rect 8289 -1070 8295 -1069
rect 8466 -1070 8589 -1058
rect 8289 -1103 8472 -1070
rect 8172 -1104 8472 -1103
rect 8506 -1104 8549 -1070
rect 8583 -1104 8589 -1070
rect 8172 -1147 8589 -1104
rect 8172 -1181 8178 -1147
rect 8212 -1181 8255 -1147
rect 8289 -1148 8589 -1147
rect 8289 -1181 8472 -1148
rect 8172 -1182 8472 -1181
rect 8506 -1182 8549 -1148
rect 8583 -1182 8589 -1148
rect 8172 -1185 8589 -1182
rect 8172 -1193 8295 -1185
rect 8466 -1194 8589 -1185
rect 5194 -1206 5317 -1194
rect 6681 -1413 6727 -1411
rect 6681 -1423 6735 -1413
rect 1364 -1485 1410 -1431
rect 6681 -1457 6687 -1423
rect 6721 -1457 6735 -1423
rect 1364 -1500 1916 -1485
rect 1364 -1531 1788 -1500
rect 1776 -1534 1788 -1531
rect 1822 -1534 1866 -1500
rect 1900 -1531 1916 -1500
rect 6681 -1501 6735 -1457
rect 1900 -1534 1912 -1531
rect 1776 -1540 1912 -1534
rect 6681 -1535 6687 -1501
rect 6721 -1535 6735 -1501
rect 6681 -1547 6735 -1535
rect -1330 -1603 -383 -1575
rect 6510 -1591 6646 -1585
rect 6510 -1625 6522 -1591
rect 6556 -1625 6600 -1591
rect 6634 -1625 6646 -1591
rect 6510 -1631 6646 -1625
rect -1330 -1747 -363 -1719
rect 6536 -2240 6582 -1631
rect 4833 -2246 6582 -2240
rect 4833 -2280 4845 -2246
rect 4879 -2280 4923 -2246
rect 4957 -2280 6582 -2246
rect 4833 -2286 6582 -2280
rect 6689 -2352 6735 -1547
rect 8087 -1666 8228 -1658
rect 8087 -1700 8099 -1666
rect 8133 -1700 8177 -1666
rect 8211 -1700 8228 -1666
rect 8087 -1711 8228 -1700
rect 8171 -2160 8228 -1711
rect 14490 -1992 14790 -1928
rect 8171 -2217 8412 -2160
rect 3265 -2358 6735 -2352
rect 3265 -2392 3277 -2358
rect 3311 -2392 3355 -2358
rect 3389 -2392 6735 -2358
rect 3265 -2398 6735 -2392
use 3AND_MAGIC#0  3AND_MAGIC_0
timestamp 1717691374
transform 1 0 6767 0 1 -1514
box -48 -929 1456 459
use 3AND_MAGIC#0  3AND_MAGIC_1
timestamp 1717691374
transform 1 0 1805 0 1 -1505
box -48 -929 1456 459
use AND_1#0  AND_1_0
timestamp 1717691374
transform 1 0 5103 0 1 -2225
box -45 -99 1479 1172
use AND_1#0  AND_1_1
timestamp 1717691374
transform 1 0 3498 0 1 -2227
box -45 -99 1479 1172
use DFF_MAG  DFF_MAG_0
timestamp 1717691374
transform 1 0 11001 0 1 -1840
box -2652 -1119 3660 811
use XNOR_MAGIC  XNOR_MAGIC_0
timestamp 1717691374
transform 1 0 10241 0 1 612
box -241 -624 1822 598
use XNOR_MAGIC  XNOR_MAGIC_1
timestamp 1717691374
transform 1 0 -259 0 1 612
box -241 -624 1822 598
use XNOR_MAGIC  XNOR_MAGIC_2
timestamp 1717691374
transform 1 0 2741 0 1 612
box -241 -624 1822 598
use XNOR_MAGIC  XNOR_MAGIC_3
timestamp 1717691374
transform 1 0 5241 0 1 612
box -241 -624 1822 598
use XNOR_MAGIC  XNOR_MAGIC_4
timestamp 1717691374
transform 1 0 7741 0 1 612
box -241 -624 1822 598
use XNOR_MAGIC  XNOR_MAGIC_5
timestamp 1717691374
transform 1 0 12741 0 1 612
box -241 -624 1822 598
use XNOR_MAGIC  XNOR_MAGIC_6
timestamp 1717691374
transform 1 0 -269 0 1 -1639
box -241 -624 1822 598
<< labels >>
flabel locali s 3305 -2219 3305 -2219 0 FreeSans 600 0 0 0 3_in_and_out
flabel metal1 s -678 -1588 -678 -1588 0 FreeSans 1000 0 0 0 Q3
flabel metal1 s -674 -1743 -674 -1743 0 FreeSans 1000 0 0 0 D2_4
flabel metal1 s -571 521 -571 521 0 FreeSans 1000 0 0 0 D2_2
flabel metal1 s -588 656 -588 656 0 FreeSans 1000 0 0 0 Q1
flabel metal1 s -310 -109 -310 -109 0 FreeSans 1000 0 0 0 D2_3
flabel metal1 s -114 -177 -114 -177 0 FreeSans 1000 0 0 0 Q4
flabel metal1 s 12 -256 12 -256 0 FreeSans 1000 0 0 0 D2_5
flabel metal1 s 231 -316 231 -316 0 FreeSans 1000 0 0 0 Q5
flabel metal1 s 454 -453 454 -453 0 FreeSans 1000 0 0 0 Q6
flabel metal1 s 633 -588 633 -588 0 FreeSans 1000 0 0 0 Q7
flabel metal1 s 402 -372 402 -372 0 FreeSans 1000 0 0 0 D2_6
flabel metal1 s 624 -520 624 -520 0 FreeSans 1000 0 0 0 D2_7
flabel metal1 s 820 -660 820 -660 0 FreeSans 1000 0 0 0 D2_1
flabel metal1 s 14758 -1962 14758 -1962 0 FreeSans 1600 0 0 0 P2
flabel locali s 8554 1307 8554 1307 0 FreeSans 1600 0 0 0 VDD
flabel locali s 5926 -2804 5926 -2804 0 FreeSans 1600 0 0 0 VSS
flabel metal1 s 235 -929 235 -929 0 FreeSans 1600 0 0 0 CLK
flabel metal1 s -392 -44 -392 -44 0 FreeSans 1600 0 0 0 Q2
<< end >>
