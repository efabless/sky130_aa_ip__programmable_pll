magic
tech sky130A
magscale 1 2
timestamp 1717691374
<< nwell >>
rect -523 -462 523 462
<< pmos >>
rect -429 -400 -29 400
rect 29 -400 429 400
<< pdiff >>
rect -487 357 -429 400
rect -487 323 -475 357
rect -441 323 -429 357
rect -487 289 -429 323
rect -487 255 -475 289
rect -441 255 -429 289
rect -487 221 -429 255
rect -487 187 -475 221
rect -441 187 -429 221
rect -487 153 -429 187
rect -487 119 -475 153
rect -441 119 -429 153
rect -487 85 -429 119
rect -487 51 -475 85
rect -441 51 -429 85
rect -487 17 -429 51
rect -487 -17 -475 17
rect -441 -17 -429 17
rect -487 -51 -429 -17
rect -487 -85 -475 -51
rect -441 -85 -429 -51
rect -487 -119 -429 -85
rect -487 -153 -475 -119
rect -441 -153 -429 -119
rect -487 -187 -429 -153
rect -487 -221 -475 -187
rect -441 -221 -429 -187
rect -487 -255 -429 -221
rect -487 -289 -475 -255
rect -441 -289 -429 -255
rect -487 -323 -429 -289
rect -487 -357 -475 -323
rect -441 -357 -429 -323
rect -487 -400 -429 -357
rect -29 357 29 400
rect -29 323 -17 357
rect 17 323 29 357
rect -29 289 29 323
rect -29 255 -17 289
rect 17 255 29 289
rect -29 221 29 255
rect -29 187 -17 221
rect 17 187 29 221
rect -29 153 29 187
rect -29 119 -17 153
rect 17 119 29 153
rect -29 85 29 119
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -119 29 -85
rect -29 -153 -17 -119
rect 17 -153 29 -119
rect -29 -187 29 -153
rect -29 -221 -17 -187
rect 17 -221 29 -187
rect -29 -255 29 -221
rect -29 -289 -17 -255
rect 17 -289 29 -255
rect -29 -323 29 -289
rect -29 -357 -17 -323
rect 17 -357 29 -323
rect -29 -400 29 -357
rect 429 357 487 400
rect 429 323 441 357
rect 475 323 487 357
rect 429 289 487 323
rect 429 255 441 289
rect 475 255 487 289
rect 429 221 487 255
rect 429 187 441 221
rect 475 187 487 221
rect 429 153 487 187
rect 429 119 441 153
rect 475 119 487 153
rect 429 85 487 119
rect 429 51 441 85
rect 475 51 487 85
rect 429 17 487 51
rect 429 -17 441 17
rect 475 -17 487 17
rect 429 -51 487 -17
rect 429 -85 441 -51
rect 475 -85 487 -51
rect 429 -119 487 -85
rect 429 -153 441 -119
rect 475 -153 487 -119
rect 429 -187 487 -153
rect 429 -221 441 -187
rect 475 -221 487 -187
rect 429 -255 487 -221
rect 429 -289 441 -255
rect 475 -289 487 -255
rect 429 -323 487 -289
rect 429 -357 441 -323
rect 475 -357 487 -323
rect 429 -400 487 -357
<< pdiffc >>
rect -475 323 -441 357
rect -475 255 -441 289
rect -475 187 -441 221
rect -475 119 -441 153
rect -475 51 -441 85
rect -475 -17 -441 17
rect -475 -85 -441 -51
rect -475 -153 -441 -119
rect -475 -221 -441 -187
rect -475 -289 -441 -255
rect -475 -357 -441 -323
rect -17 323 17 357
rect -17 255 17 289
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect -17 -289 17 -255
rect -17 -357 17 -323
rect 441 323 475 357
rect 441 255 475 289
rect 441 187 475 221
rect 441 119 475 153
rect 441 51 475 85
rect 441 -17 475 17
rect 441 -85 475 -51
rect 441 -153 475 -119
rect 441 -221 475 -187
rect 441 -289 475 -255
rect 441 -357 475 -323
<< poly >>
rect -429 400 -29 426
rect 29 400 429 426
rect -429 -426 -29 -400
rect 29 -426 429 -400
<< locali >>
rect -475 377 -441 404
rect -475 305 -441 323
rect -475 233 -441 255
rect -475 161 -441 187
rect -475 89 -441 119
rect -475 17 -441 51
rect -475 -51 -441 -17
rect -475 -119 -441 -89
rect -475 -187 -441 -161
rect -475 -255 -441 -233
rect -475 -323 -441 -305
rect -475 -404 -441 -377
rect -17 377 17 404
rect -17 305 17 323
rect -17 233 17 255
rect -17 161 17 187
rect -17 89 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -89
rect -17 -187 17 -161
rect -17 -255 17 -233
rect -17 -323 17 -305
rect -17 -404 17 -377
rect 441 377 475 404
rect 441 305 475 323
rect 441 233 475 255
rect 441 161 475 187
rect 441 89 475 119
rect 441 17 475 51
rect 441 -51 475 -17
rect 441 -119 475 -89
rect 441 -187 475 -161
rect 441 -255 475 -233
rect 441 -323 475 -305
rect 441 -404 475 -377
<< viali >>
rect -475 357 -441 377
rect -475 343 -441 357
rect -475 289 -441 305
rect -475 271 -441 289
rect -475 221 -441 233
rect -475 199 -441 221
rect -475 153 -441 161
rect -475 127 -441 153
rect -475 85 -441 89
rect -475 55 -441 85
rect -475 -17 -441 17
rect -475 -85 -441 -55
rect -475 -89 -441 -85
rect -475 -153 -441 -127
rect -475 -161 -441 -153
rect -475 -221 -441 -199
rect -475 -233 -441 -221
rect -475 -289 -441 -271
rect -475 -305 -441 -289
rect -475 -357 -441 -343
rect -475 -377 -441 -357
rect -17 357 17 377
rect -17 343 17 357
rect -17 289 17 305
rect -17 271 17 289
rect -17 221 17 233
rect -17 199 17 221
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect -17 -221 17 -199
rect -17 -233 17 -221
rect -17 -289 17 -271
rect -17 -305 17 -289
rect -17 -357 17 -343
rect -17 -377 17 -357
rect 441 357 475 377
rect 441 343 475 357
rect 441 289 475 305
rect 441 271 475 289
rect 441 221 475 233
rect 441 199 475 221
rect 441 153 475 161
rect 441 127 475 153
rect 441 85 475 89
rect 441 55 475 85
rect 441 -17 475 17
rect 441 -85 475 -55
rect 441 -89 475 -85
rect 441 -153 475 -127
rect 441 -161 475 -153
rect 441 -221 475 -199
rect 441 -233 475 -221
rect 441 -289 475 -271
rect 441 -305 475 -289
rect 441 -357 475 -343
rect 441 -377 475 -357
<< metal1 >>
rect -481 377 -435 400
rect -481 343 -475 377
rect -441 343 -435 377
rect -481 305 -435 343
rect -481 271 -475 305
rect -441 271 -435 305
rect -481 233 -435 271
rect -481 199 -475 233
rect -441 199 -435 233
rect -481 161 -435 199
rect -481 127 -475 161
rect -441 127 -435 161
rect -481 89 -435 127
rect -481 55 -475 89
rect -441 55 -435 89
rect -481 17 -435 55
rect -481 -17 -475 17
rect -441 -17 -435 17
rect -481 -55 -435 -17
rect -481 -89 -475 -55
rect -441 -89 -435 -55
rect -481 -127 -435 -89
rect -481 -161 -475 -127
rect -441 -161 -435 -127
rect -481 -199 -435 -161
rect -481 -233 -475 -199
rect -441 -233 -435 -199
rect -481 -271 -435 -233
rect -481 -305 -475 -271
rect -441 -305 -435 -271
rect -481 -343 -435 -305
rect -481 -377 -475 -343
rect -441 -377 -435 -343
rect -481 -400 -435 -377
rect -23 377 23 400
rect -23 343 -17 377
rect 17 343 23 377
rect -23 305 23 343
rect -23 271 -17 305
rect 17 271 23 305
rect -23 233 23 271
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -271 23 -233
rect -23 -305 -17 -271
rect 17 -305 23 -271
rect -23 -343 23 -305
rect -23 -377 -17 -343
rect 17 -377 23 -343
rect -23 -400 23 -377
rect 435 377 481 400
rect 435 343 441 377
rect 475 343 481 377
rect 435 305 481 343
rect 435 271 441 305
rect 475 271 481 305
rect 435 233 481 271
rect 435 199 441 233
rect 475 199 481 233
rect 435 161 481 199
rect 435 127 441 161
rect 475 127 481 161
rect 435 89 481 127
rect 435 55 441 89
rect 475 55 481 89
rect 435 17 481 55
rect 435 -17 441 17
rect 475 -17 481 17
rect 435 -55 481 -17
rect 435 -89 441 -55
rect 475 -89 481 -55
rect 435 -127 481 -89
rect 435 -161 441 -127
rect 475 -161 481 -127
rect 435 -199 481 -161
rect 435 -233 441 -199
rect 475 -233 481 -199
rect 435 -271 481 -233
rect 435 -305 441 -271
rect 475 -305 481 -271
rect 435 -343 481 -305
rect 435 -377 441 -343
rect 475 -377 481 -343
rect 435 -400 481 -377
<< end >>
