magic
tech sky130A
magscale 1 2
timestamp 1717691374
<< nwell >>
rect -2036 2206 -1189 2359
rect -1798 2133 -1753 2206
rect -1376 2132 -1331 2206
rect -1633 1482 -1495 1523
<< pwell >>
rect -2005 715 -1206 849
<< psubdiff >>
rect -1979 798 -1232 823
rect -1979 764 -1936 798
rect -1902 764 -1868 798
rect -1834 764 -1800 798
rect -1766 764 -1732 798
rect -1698 764 -1664 798
rect -1630 764 -1596 798
rect -1562 764 -1528 798
rect -1494 764 -1460 798
rect -1426 764 -1392 798
rect -1358 764 -1324 798
rect -1290 764 -1232 798
rect -1979 741 -1232 764
<< nsubdiff >>
rect -1999 2306 -1230 2322
rect -1999 2272 -1939 2306
rect -1905 2272 -1871 2306
rect -1837 2272 -1803 2306
rect -1769 2272 -1735 2306
rect -1701 2272 -1667 2306
rect -1633 2272 -1599 2306
rect -1565 2272 -1531 2306
rect -1497 2272 -1463 2306
rect -1429 2272 -1395 2306
rect -1361 2272 -1327 2306
rect -1293 2272 -1230 2306
rect -1999 2256 -1230 2272
<< psubdiffcont >>
rect -1936 764 -1902 798
rect -1868 764 -1834 798
rect -1800 764 -1766 798
rect -1732 764 -1698 798
rect -1664 764 -1630 798
rect -1596 764 -1562 798
rect -1528 764 -1494 798
rect -1460 764 -1426 798
rect -1392 764 -1358 798
rect -1324 764 -1290 798
<< nsubdiffcont >>
rect -1939 2272 -1905 2306
rect -1871 2272 -1837 2306
rect -1803 2272 -1769 2306
rect -1735 2272 -1701 2306
rect -1667 2272 -1633 2306
rect -1599 2272 -1565 2306
rect -1531 2272 -1497 2306
rect -1463 2272 -1429 2306
rect -1395 2272 -1361 2306
rect -1327 2272 -1293 2306
<< poly >>
rect -1942 1482 -1804 1523
rect -1844 1325 -1804 1482
rect -1999 1314 -1804 1325
rect -1999 1280 -1983 1314
rect -1949 1280 -1897 1314
rect -1863 1280 -1804 1314
rect -1999 1270 -1804 1280
rect -1844 1258 -1804 1270
rect -1746 1482 -1495 1523
rect -1746 1433 -1706 1482
rect -1323 1455 -1283 1532
rect -1462 1444 -1283 1455
rect -1746 1422 -1574 1433
rect -1746 1388 -1713 1422
rect -1679 1388 -1627 1422
rect -1593 1388 -1574 1422
rect -1462 1410 -1445 1444
rect -1411 1410 -1359 1444
rect -1325 1410 -1283 1444
rect -1462 1400 -1283 1410
rect -1746 1378 -1574 1388
rect -1746 1257 -1706 1378
rect -1323 1310 -1283 1400
rect -1406 1270 -1283 1310
rect -1406 1258 -1365 1270
<< polycont >>
rect -1983 1280 -1949 1314
rect -1897 1280 -1863 1314
rect -1713 1388 -1679 1422
rect -1627 1388 -1593 1422
rect -1445 1410 -1411 1444
rect -1359 1410 -1325 1444
<< locali >>
rect -1999 2306 -1230 2322
rect -1999 2272 -1939 2306
rect -1905 2272 -1871 2306
rect -1837 2272 -1803 2306
rect -1769 2272 -1735 2306
rect -1701 2272 -1667 2306
rect -1633 2272 -1599 2306
rect -1565 2272 -1531 2306
rect -1497 2272 -1463 2306
rect -1429 2272 -1395 2306
rect -1361 2272 -1327 2306
rect -1293 2272 -1230 2306
rect -1999 2256 -1230 2272
rect -1993 2130 -1948 2256
rect -1798 2133 -1753 2256
rect -1683 2182 -1443 2216
rect -1683 2140 -1641 2182
rect -1485 2138 -1443 2182
rect -1376 2132 -1331 2256
rect -1894 1505 -1852 1564
rect -1682 1505 -1640 1558
rect -1894 1469 -1640 1505
rect -1585 1506 -1543 1560
rect -1585 1467 -1444 1506
rect -1487 1455 -1444 1467
rect -1487 1444 -1306 1455
rect -1729 1423 -1574 1433
rect -2033 1422 -1574 1423
rect -2033 1388 -1713 1422
rect -1679 1388 -1627 1422
rect -1593 1388 -1574 1422
rect -2033 1387 -1574 1388
rect -1729 1378 -1574 1387
rect -1487 1410 -1445 1444
rect -1411 1410 -1359 1444
rect -1325 1410 -1306 1444
rect -1487 1400 -1306 1410
rect -1487 1330 -1444 1400
rect -1999 1316 -1844 1325
rect -2036 1314 -1844 1316
rect -2036 1282 -1983 1314
rect -1999 1280 -1983 1282
rect -1949 1280 -1897 1314
rect -1863 1280 -1844 1314
rect -1999 1270 -1844 1280
rect -1798 1290 -1444 1330
rect -1272 1310 -1229 1554
rect -1798 1220 -1753 1290
rect -1406 1270 -1191 1310
rect -1358 1267 -1191 1270
rect -1358 1227 -1314 1267
rect -1897 823 -1850 942
rect -1701 823 -1654 943
rect -1459 823 -1412 953
rect -1979 798 -1232 823
rect -1979 764 -1936 798
rect -1902 764 -1868 798
rect -1834 764 -1800 798
rect -1766 764 -1732 798
rect -1698 764 -1664 798
rect -1630 764 -1596 798
rect -1562 764 -1528 798
rect -1494 764 -1460 798
rect -1426 764 -1392 798
rect -1358 764 -1324 798
rect -1290 764 -1232 798
rect -1979 741 -1232 764
use sky130_fd_pr__nfet_01v8_FQGQPX  sky130_fd_pr__nfet_01v8_FQGQPX_0
timestamp 1717691374
transform 1 0 -1386 0 1 1082
box -104 -176 104 176
use sky130_fd_pr__nfet_01v8_FQGQPX  sky130_fd_pr__nfet_01v8_FQGQPX_1
timestamp 1717691374
transform 1 0 -1824 0 1 1082
box -104 -176 104 176
use sky130_fd_pr__nfet_01v8_FQGQPX  sky130_fd_pr__nfet_01v8_FQGQPX_2
timestamp 1717691374
transform 1 0 -1726 0 1 1082
box -104 -176 104 176
use sky130_fd_pr__pfet_01v8_6WH9DB  sky130_fd_pr__pfet_01v8_6WH9DB_0
timestamp 1717691374
transform 1 0 -1303 0 1 1844
box -114 -362 114 362
use sky130_fd_pr__pfet_01v8_6WH9DB  sky130_fd_pr__pfet_01v8_6WH9DB_1
timestamp 1717691374
transform 1 0 -1613 0 1 1844
box -114 -362 114 362
use sky130_fd_pr__pfet_01v8_6WH9DB  sky130_fd_pr__pfet_01v8_6WH9DB_2
timestamp 1717691374
transform 1 0 -1824 0 1 1844
box -114 -362 114 362
use sky130_fd_pr__pfet_01v8_6WH9DB  sky130_fd_pr__pfet_01v8_6WH9DB_3
timestamp 1717691374
transform 1 0 -1922 0 1 1844
box -114 -362 114 362
use sky130_fd_pr__pfet_01v8_6WH9DB  sky130_fd_pr__pfet_01v8_6WH9DB_4
timestamp 1717691374
transform 1 0 -1515 0 1 1844
box -114 -362 114 362
<< labels >>
flabel locali s -1635 2316 -1635 2316 0 FreeSans 1000 0 0 0 VDD
flabel locali s -1208 1292 -1208 1292 0 FreeSans 1000 0 0 0 VOUT
flabel locali s -2025 1400 -2025 1400 0 FreeSans 1000 0 0 0 A
flabel locali s -2024 1295 -2024 1295 0 FreeSans 1000 0 0 0 B
flabel locali s -1635 748 -1635 748 0 FreeSans 1000 0 0 0 VSS
<< end >>
