magic
tech sky130A
magscale 1 2
timestamp 1717691374
<< locali >>
rect -289 9526 60859 10629
rect -9356 8898 -9159 8933
rect -9356 8792 -9314 8898
rect -9208 8792 -9159 8898
rect -9356 8752 -9159 8792
rect -9700 8438 -9419 8486
rect -9700 8332 -9649 8438
rect -9471 8332 -9419 8438
rect -9700 8277 -9419 8332
rect -10060 8017 -9698 8120
rect -10060 7911 -9951 8017
rect -9773 7911 -9698 8017
rect -10060 7849 -9698 7911
rect -10247 6573 -10012 6596
rect -15441 6508 -10012 6573
rect -15441 6402 -10179 6508
rect -10073 6402 -10012 6508
rect -15441 6328 -10012 6402
rect -15441 6326 -10136 6328
rect -10333 6157 -10066 6193
rect -15678 6090 -10066 6157
rect -15678 5984 -10248 6090
rect -10142 5984 -10066 6090
rect -15678 5922 -10066 5984
rect -10333 5895 -10066 5922
rect -9835 4937 -9707 7849
rect -9582 5026 -9450 8277
rect -9340 5118 -9251 8752
rect -7831 7032 58142 7538
rect -8476 6564 -8258 6639
rect -8476 6458 -8430 6564
rect -8324 6458 -8258 6564
rect -8476 6393 -8258 6458
rect -8437 5536 -8295 6393
rect -8474 5487 -8295 5536
rect -7248 5513 -6703 7032
rect -235 6563 95 6616
rect -235 6385 -193 6563
rect 57 6533 95 6563
rect 2498 6534 2781 7032
rect 7866 6577 8223 6623
rect 57 6488 944 6533
rect 57 6385 698 6488
rect -235 6382 698 6385
rect 876 6382 944 6488
rect -235 6354 944 6382
rect 7866 6399 7918 6577
rect 8168 6556 8223 6577
rect 9044 6556 9401 6589
rect 8168 6543 9401 6556
rect 8168 6399 9096 6543
rect 7866 6367 9096 6399
rect 7866 6356 8223 6367
rect 9044 6365 9096 6367
rect 9346 6365 9401 6543
rect 10897 6497 11180 7032
rect -235 6322 95 6354
rect 9044 6322 9401 6365
rect 16422 6467 16687 6498
rect 17948 6467 18245 6500
rect 19809 6470 20092 7032
rect 26939 6475 27185 6544
rect 29028 6515 29311 7032
rect 34377 6612 34753 6682
rect 16422 6455 18245 6467
rect 16422 6277 16459 6455
rect 16637 6445 18245 6455
rect 16637 6339 18005 6445
rect 18183 6339 18245 6445
rect 16637 6300 18245 6339
rect 16637 6277 16687 6300
rect 17948 6278 18245 6300
rect 25286 6464 25512 6473
rect 26939 6464 27011 6475
rect 25286 6443 27011 6464
rect 16422 6233 16687 6277
rect 25286 6265 25339 6443
rect 25445 6369 27011 6443
rect 27117 6369 27185 6475
rect 25445 6331 27185 6369
rect 34377 6434 34450 6612
rect 34700 6587 34753 6612
rect 35978 6587 36228 6614
rect 34700 6549 36228 6587
rect 37823 6580 38130 7032
rect 43153 6616 43491 6677
rect 34700 6443 36003 6549
rect 36181 6443 36228 6549
rect 34700 6436 36228 6443
rect 34700 6434 34753 6436
rect 34377 6368 34753 6434
rect 35978 6385 36228 6436
rect 43153 6438 43235 6616
rect 43413 6581 43491 6616
rect 45141 6581 45409 6622
rect 46929 6601 47269 7032
rect 52383 6650 52653 6763
rect 43413 6551 45409 6581
rect 43413 6450 45233 6551
rect 43413 6438 43491 6450
rect 43153 6386 43491 6438
rect 45141 6445 45233 6450
rect 45339 6445 45409 6551
rect 52383 6544 52479 6650
rect 52585 6642 52653 6650
rect 54396 6642 54691 6684
rect 52585 6612 54691 6642
rect 56265 6625 56476 7032
rect 52585 6544 54506 6612
rect 52383 6506 54506 6544
rect 54612 6506 54691 6612
rect 52383 6503 54691 6506
rect 52383 6478 52653 6503
rect 45141 6382 45409 6445
rect 54396 6411 54691 6503
rect 25445 6265 25512 6331
rect 26939 6324 27185 6331
rect 25286 6239 25512 6265
rect -8474 5381 -8440 5487
rect -8334 5381 -8295 5487
rect -8474 5347 -8295 5381
rect -735 5316 1578 5610
rect 7197 5221 10085 5374
rect 14666 5286 18962 5540
rect 23517 5276 28145 5590
rect 32700 5308 36859 5687
rect 41447 5402 46033 5666
rect 50609 5393 55441 5735
rect 60384 5550 60859 9526
rect -9340 5077 -8304 5118
rect -9582 4985 -8160 5026
rect -9835 4896 -8130 4937
rect 684 4763 943 4806
rect -182 4720 943 4763
rect -182 4706 762 4720
rect -182 4600 -159 4706
rect 19 4614 762 4706
rect 868 4614 943 4720
rect 19 4600 943 4614
rect -182 4558 943 4600
rect 684 4543 943 4558
rect 8685 4549 9333 4695
rect -11964 3482 -11450 3576
rect -11964 3232 -11787 3482
rect -11537 3413 -11450 3482
rect -10204 3413 -9983 3441
rect -11537 3395 -9983 3413
rect -11537 3289 -10147 3395
rect -10041 3289 -9983 3395
rect -11537 3283 -9983 3289
rect -11537 3232 -11450 3283
rect -10204 3261 -9983 3283
rect 375 3415 1219 3446
rect 375 3339 1247 3415
rect 375 3300 1219 3339
rect -11964 3151 -11450 3232
rect -13434 2549 -13149 2570
rect -13434 2371 -13417 2549
rect -13167 2512 -13149 2549
rect -13167 2484 -8474 2512
rect -13167 2448 -8191 2484
rect -13167 2418 -8474 2448
rect -13167 2371 -13149 2418
rect -13434 2351 -13149 2371
rect -8371 2359 -8166 2395
rect -8371 2306 -8335 2359
rect -12452 2280 -8335 2306
rect -12452 2174 -12350 2280
rect -12244 2174 -8335 2280
rect -12452 2144 -8335 2174
rect 375 -450 521 3300
rect 7973 833 8196 868
rect 7921 735 7962 742
rect 7973 727 8028 833
rect 8134 727 8196 833
rect 7973 698 8196 727
rect -1491 -452 521 -450
rect -1491 -486 540 -452
rect -1491 -592 -1267 -486
rect -1017 -487 540 -486
rect -1017 -592 402 -487
rect -1491 -593 402 -592
rect 508 -593 540 -487
rect -1491 -620 540 -593
rect -1491 -621 464 -620
rect 390 -865 611 -819
rect 390 -971 442 -865
rect 548 -971 611 -865
rect 390 -1014 611 -971
rect 960 -1226 1096 159
rect 8685 -834 8831 4549
rect 17367 4463 18134 4609
rect 26686 4555 27415 4701
rect 35213 4587 36139 4826
rect 44541 4613 45205 4798
rect 53458 4646 54666 4940
rect 8955 3625 9680 3657
rect 8955 3549 9687 3625
rect 8955 3511 9680 3549
rect 8955 -472 9101 3511
rect 16422 878 16759 930
rect 16422 628 16482 878
rect 16660 628 16759 878
rect 16422 599 16759 628
rect 8932 -492 9135 -472
rect 8932 -598 8973 -492
rect 9079 -598 9135 -492
rect 8932 -619 9135 -598
rect 8616 -880 8890 -834
rect 8616 -986 8658 -880
rect 8836 -986 8890 -880
rect 8616 -1037 8890 -986
rect -14981 -1362 1096 -1226
rect 9400 -1425 9536 173
rect 16063 -447 16380 -362
rect 16063 -625 16126 -447
rect 16304 -625 16380 -447
rect 16063 -653 16380 -625
rect -14886 -1561 9536 -1425
rect 16080 -1242 16346 -653
rect 17367 -852 17513 4463
rect 17824 3494 18540 3530
rect 17824 3418 18550 3494
rect 17824 3384 18540 3418
rect 17824 -494 17970 3384
rect 25300 822 25514 843
rect 25300 644 25318 822
rect 25496 644 25514 822
rect 25300 623 25514 644
rect 17824 -600 17841 -494
rect 17947 -600 17970 -494
rect 17824 -617 17970 -600
rect 17313 -869 17565 -852
rect 17313 -975 17348 -869
rect 17526 -975 17565 -869
rect 17313 -991 17565 -975
rect 16080 -1420 16128 -1242
rect 16306 -1420 16346 -1242
rect 16080 -1433 16346 -1420
rect 16097 -1442 16337 -1433
rect 18310 -1658 18446 100
rect 26686 -813 26832 4555
rect 26961 3596 27738 3631
rect 26961 3520 27748 3596
rect 26961 3470 27738 3520
rect 26961 -451 27122 3470
rect 34426 840 34718 931
rect 34426 662 34496 840
rect 34674 662 34718 840
rect 34426 632 34718 662
rect 26943 -484 27137 -451
rect 26943 -590 26991 -484
rect 27097 -590 27137 -484
rect 26943 -618 27137 -590
rect 26652 -863 26884 -813
rect 26652 -969 26712 -863
rect 26818 -969 26884 -863
rect 26652 -1018 26884 -969
rect -14862 -1794 18446 -1658
rect 27461 -1913 27597 220
rect 35213 -798 35452 4587
rect 35713 3568 36463 3604
rect 35713 3492 36502 3568
rect 35713 3387 36463 3492
rect 35151 -816 35499 -798
rect 35151 -994 35203 -816
rect 35453 -994 35499 -816
rect 35151 -1030 35499 -994
rect 35713 -1183 35930 3387
rect 43191 918 43452 989
rect 43191 740 43246 918
rect 43424 740 43452 918
rect 43191 685 43452 740
rect 35656 -1194 36000 -1183
rect 35656 -1444 35703 -1194
rect 35953 -1444 36000 -1194
rect 35656 -1466 36000 -1444
rect -15052 -2049 27597 -1913
rect 36215 -2199 36351 250
rect 44541 -795 44726 4613
rect 44904 3393 45621 3563
rect 44904 -443 45074 3393
rect 52477 841 52579 883
rect 52477 807 52506 841
rect 52540 807 52579 841
rect 52477 772 52579 807
rect 44865 -483 45111 -443
rect 44865 -589 44897 -483
rect 45075 -589 45111 -483
rect 44865 -623 45111 -589
rect 44456 -831 44838 -795
rect 44456 -1009 44513 -831
rect 44763 -1009 44838 -831
rect 44456 -1040 44838 -1009
rect -15052 -2335 36351 -2199
rect 45368 -2498 45504 222
rect 53458 -798 53752 4646
rect 54180 3416 55061 3642
rect 53409 -828 53809 -798
rect 53409 -1006 53437 -828
rect 53759 -1006 53809 -828
rect 53409 -1036 53809 -1006
rect 54180 -1186 54406 3416
rect 61868 957 62227 1033
rect 61868 779 61973 957
rect 62151 779 62227 957
rect 61868 690 62227 779
rect 54091 -1235 54478 -1186
rect 54091 -1413 54164 -1235
rect 54414 -1413 54478 -1235
rect 54091 -1462 54478 -1413
rect -14981 -2634 45504 -2498
rect 54756 -2868 54892 241
rect -14933 -3004 54892 -2868
<< viali >>
rect -9314 8792 -9208 8898
rect -9649 8332 -9471 8438
rect -9951 7911 -9773 8017
rect -10179 6402 -10073 6508
rect -10248 5984 -10142 6090
rect -8430 6458 -8324 6564
rect -193 6385 57 6563
rect 698 6382 876 6488
rect 7918 6399 8168 6577
rect 9096 6365 9346 6543
rect 16459 6277 16637 6455
rect 18005 6339 18183 6445
rect 25339 6265 25445 6443
rect 27011 6369 27117 6475
rect 34450 6434 34700 6612
rect 36003 6443 36181 6549
rect 43235 6438 43413 6616
rect 45233 6445 45339 6551
rect 52479 6544 52585 6650
rect 54506 6506 54612 6612
rect -8440 5381 -8334 5487
rect -159 4600 19 4706
rect 762 4614 868 4720
rect -11787 3232 -11537 3482
rect -10147 3289 -10041 3395
rect -13417 2371 -13167 2549
rect -12350 2174 -12244 2280
rect 8028 727 8134 833
rect -1267 -592 -1017 -486
rect 402 -593 508 -487
rect 442 -971 548 -865
rect 16482 628 16660 878
rect 8973 -598 9079 -492
rect 8658 -986 8836 -880
rect 16126 -625 16304 -447
rect 25318 644 25496 822
rect 17841 -600 17947 -494
rect 17348 -975 17526 -869
rect 16128 -1420 16306 -1242
rect 34496 662 34674 840
rect 26991 -590 27097 -484
rect 26712 -969 26818 -863
rect 35203 -994 35453 -816
rect 43246 740 43424 918
rect 35703 -1444 35953 -1194
rect 52506 807 52540 841
rect 44897 -589 45075 -483
rect 44513 -1009 44763 -831
rect 53437 -1006 53759 -828
rect 61973 779 62151 957
rect 54164 -1413 54414 -1235
<< metal1 >>
rect -13439 11242 62182 11526
rect -13439 2616 -13170 11242
rect -12447 10309 52678 10620
rect -13500 2549 -13114 2616
rect -13500 2371 -13417 2549
rect -13167 2371 -13114 2549
rect -13500 2275 -13114 2371
rect -12447 2326 -12196 10309
rect -11860 9859 43410 10036
rect -11860 3576 -11529 9859
rect -10748 9300 34701 9521
rect -11964 3482 -11450 3576
rect -11964 3232 -11787 3482
rect -11537 3232 -11450 3482
rect -11964 3151 -11450 3232
rect -10748 3027 -10658 9300
rect -9367 8898 25512 8969
rect -9367 8792 -9314 8898
rect -9208 8792 25512 8898
rect -9367 8743 25512 8792
rect -9759 8438 16687 8528
rect -9759 8332 -9649 8438
rect -9471 8332 16687 8438
rect -9759 8263 16687 8332
rect -10041 8017 8206 8106
rect -10041 7911 -9951 8017
rect -9773 7911 8206 8017
rect -10041 7857 8206 7911
rect 385 6745 6850 6914
rect -10318 6616 -85 6656
rect -10318 6564 95 6616
rect -10318 6508 -8430 6564
rect -10318 6402 -10179 6508
rect -10073 6458 -8430 6508
rect -8324 6563 95 6564
rect -8324 6458 -193 6563
rect -10073 6402 -193 6458
rect -10318 6385 -193 6402
rect 57 6385 95 6563
rect -10318 6322 95 6385
rect -10318 6304 60 6322
rect -10333 6115 -10066 6193
rect -10333 6090 -419 6115
rect -10333 5984 -10248 6090
rect -10142 5984 -419 6090
rect -10333 5960 -419 5984
rect -10333 5895 -10066 5960
rect -8474 5487 -8295 5536
rect -8474 5381 -8440 5487
rect -8334 5460 -8295 5487
rect -8334 5385 -8115 5460
rect -8334 5381 -8295 5385
rect -8474 5347 -8295 5381
rect -574 3571 -419 5960
rect -649 3501 -419 3571
rect -185 4706 60 6304
rect -185 4600 -159 4706
rect 19 4600 60 4706
rect -10208 3395 -8098 3444
rect -10208 3289 -10147 3395
rect -10041 3289 -8098 3395
rect -10208 3248 -8098 3289
rect -8294 3242 -8098 3248
rect -8294 3053 -8096 3242
rect -8294 3046 -8098 3053
rect -10748 3014 -8765 3027
rect -10748 2972 -8093 3014
rect -10748 2937 -8765 2972
rect -409 2711 -288 2734
rect -692 2666 -288 2711
rect -12463 2280 -12175 2326
rect -12463 2174 -12350 2280
rect -12244 2174 -12175 2280
rect -12463 2096 -12175 2174
rect -683 1814 -542 1848
rect -1203 -422 -1133 1781
rect -576 1686 -542 1814
rect -1322 -486 -951 -422
rect -1322 -592 -1267 -486
rect -1017 -592 -951 -486
rect -1322 -642 -951 -592
rect -637 -971 -516 1686
rect -1917 -1092 -516 -971
rect -1917 -3935 -1796 -1092
rect -409 -3333 -288 2666
rect -185 -795 60 4600
rect 385 3097 554 6745
rect 683 6488 896 6503
rect 683 6382 698 6488
rect 876 6382 896 6488
rect 683 6370 896 6382
rect 684 4720 943 4806
rect 684 4614 762 4720
rect 868 4614 943 4720
rect 684 4543 943 4614
rect 6681 4465 6850 6745
rect 7957 6623 8206 7857
rect 8368 6797 15450 6988
rect 7866 6577 8223 6623
rect 7866 6399 7918 6577
rect 8168 6487 8223 6577
rect 8168 6433 8229 6487
rect 8168 6399 8223 6433
rect 7866 6356 8223 6399
rect 385 2928 735 3097
rect 7957 867 8206 6356
rect 8368 3083 8559 6797
rect 9044 6543 9401 6589
rect 9044 6365 9096 6543
rect 9346 6365 9401 6543
rect 9044 6322 9401 6365
rect 15234 4470 15450 6797
rect 16422 6455 16687 8263
rect 16422 6277 16459 6455
rect 16637 6277 16687 6455
rect 8368 2892 9218 3083
rect 16422 930 16687 6277
rect 16864 6804 24825 7006
rect 16864 3014 17066 6804
rect 17948 6445 18245 6500
rect 17948 6339 18005 6445
rect 18183 6339 18245 6445
rect 17948 6278 18245 6339
rect 24623 4411 24825 6804
rect 25286 6443 25512 8743
rect 25286 6265 25339 6443
rect 25445 6265 25512 6443
rect 16864 2812 18194 3014
rect 25286 1069 25512 6265
rect 26143 6739 34129 6998
rect 26143 3135 26402 6739
rect 26939 6475 27185 6544
rect 26939 6369 27011 6475
rect 27117 6448 27185 6475
rect 27117 6394 27478 6448
rect 27117 6369 27185 6394
rect 26939 6324 27185 6369
rect 33870 4421 34129 6739
rect 34480 6682 34701 9300
rect 34932 6719 42916 6957
rect 34377 6612 34753 6682
rect 34377 6434 34450 6612
rect 34700 6434 34753 6612
rect 34377 6368 34753 6434
rect 26143 2876 27351 3135
rect 16422 878 16759 930
rect 7973 833 8196 867
rect 7973 727 8028 833
rect 8134 727 8196 833
rect 7973 698 8196 727
rect 16422 628 16482 878
rect 16660 628 16759 878
rect 16422 599 16759 628
rect 25264 822 25562 1069
rect 34480 931 34701 6368
rect 34932 3195 35170 6719
rect 35978 6549 36228 6614
rect 35978 6443 36003 6549
rect 36181 6443 36228 6549
rect 35978 6385 36228 6443
rect 42678 4495 42916 6719
rect 43233 6677 43410 9859
rect 43718 6711 52106 7011
rect 43153 6616 43491 6677
rect 43153 6438 43235 6616
rect 43413 6438 43491 6616
rect 43153 6386 43491 6438
rect 34932 2957 36068 3195
rect 43233 989 43410 6386
rect 43718 3261 44018 6711
rect 45141 6551 45409 6622
rect 45141 6445 45233 6551
rect 45339 6445 45409 6551
rect 45141 6382 45409 6445
rect 51799 4526 52106 6711
rect 52367 6650 52678 10309
rect 52367 6544 52479 6650
rect 52585 6544 52678 6650
rect 43718 2961 45208 3261
rect 25264 644 25318 822
rect 25496 644 25562 822
rect 25264 569 25562 644
rect 34426 840 34718 931
rect 34426 662 34496 840
rect 34674 662 34718 840
rect 43191 918 43452 989
rect 43191 740 43246 918
rect 43424 740 43452 918
rect 43191 685 43452 740
rect 52367 841 52678 6544
rect 52943 6793 61462 7012
rect 52943 3155 53162 6793
rect 54396 6612 54691 6684
rect 54396 6506 54506 6612
rect 54612 6506 54691 6612
rect 54396 6411 54691 6506
rect 61243 4566 61462 6793
rect 52943 2936 54722 3155
rect 61898 1033 62182 11242
rect 52367 807 52506 841
rect 52540 807 52678 841
rect 52367 665 52678 807
rect 61868 957 62227 1033
rect 61868 779 61973 957
rect 62151 779 62227 957
rect 61868 690 62227 779
rect 34426 632 34718 662
rect 16063 -445 16380 -362
rect 363 -487 9163 -445
rect 363 -593 402 -487
rect 508 -492 9163 -487
rect 508 -593 8973 -492
rect 363 -598 8973 -593
rect 9079 -598 9163 -492
rect 363 -626 9163 -598
rect 16063 -447 55813 -445
rect 16063 -625 16126 -447
rect 16304 -483 55813 -447
rect 16304 -484 44897 -483
rect 16304 -494 26991 -484
rect 16304 -600 17841 -494
rect 17947 -590 26991 -494
rect 27097 -589 44897 -484
rect 45075 -589 55813 -483
rect 27097 -590 55813 -589
rect 17947 -600 55813 -590
rect 16304 -625 55813 -600
rect 16063 -626 55813 -625
rect 16063 -653 16380 -626
rect -185 -816 55813 -795
rect -185 -863 35203 -816
rect -185 -865 26712 -863
rect -185 -971 442 -865
rect 548 -869 26712 -865
rect 548 -880 17348 -869
rect 548 -971 8658 -880
rect -185 -986 8658 -971
rect 8836 -975 17348 -880
rect 17526 -969 26712 -869
rect 26818 -969 35203 -863
rect 17526 -975 35203 -969
rect 8836 -986 35203 -975
rect -185 -994 35203 -986
rect 35453 -828 55813 -816
rect 35453 -831 53437 -828
rect 35453 -994 44513 -831
rect -185 -1009 44513 -994
rect 44763 -1006 53437 -831
rect 53759 -1006 55813 -828
rect 44763 -1009 55813 -1006
rect -185 -1040 55813 -1009
rect 16020 -1242 16389 -1168
rect 16020 -1420 16128 -1242
rect 16306 -1420 16389 -1242
rect 16020 -1545 16389 -1420
rect 17340 -1194 55813 -1181
rect 17340 -1444 35703 -1194
rect 35953 -1235 55813 -1194
rect 35953 -1413 54164 -1235
rect 54414 -1413 55813 -1235
rect 35953 -1444 55813 -1413
rect 17340 -1466 55813 -1444
rect 16029 -3333 16329 -1545
rect -1449 -3633 16329 -3333
rect 17340 -3876 17625 -1466
rect -1654 -3935 17625 -3876
rect -1917 -4056 17625 -3935
rect -1654 -4161 17625 -4056
use LD_GEN_MAGIC  LD_GEN_MAGIC_0
timestamp 1717691374
transform 1 0 -8105 0 -1 5859
box -266 70 7553 4277
use mod_dff_magic  mod_dff_magic_0
timestamp 1717691374
transform 1 0 54694 0 1 3754
box -305 -3649 7647 3049
use mod_dff_magic  mod_dff_magic_1
timestamp 1717691374
transform 1 0 922 0 1 3649
box -305 -3649 7647 3049
use mod_dff_magic  mod_dff_magic_2
timestamp 1717691374
transform 1 0 9362 0 1 3638
box -305 -3649 7647 3049
use mod_dff_magic  mod_dff_magic_3
timestamp 1717691374
transform 1 0 18225 0 1 3599
box -305 -3649 7647 3049
use mod_dff_magic  mod_dff_magic_4
timestamp 1717691374
transform 1 0 27423 0 1 3633
box -305 -3649 7647 3049
use mod_dff_magic  mod_dff_magic_5
timestamp 1717691374
transform 1 0 36177 0 1 3699
box -305 -3649 7647 3049
use mod_dff_magic  mod_dff_magic_6
timestamp 1717691374
transform 1 0 45330 0 1 3716
box -305 -3649 7647 3049
<< labels >>
flabel metal1 s -1076 -3483 -1076 -3483 0 FreeSans 3125 0 0 0 LD1
flabel metal1 s -1265 -4068 -1265 -4068 0 FreeSans 3125 0 0 0 LD2
flabel locali s -1375 -550 -1375 -550 0 FreeSans 3125 0 0 0 LD3
flabel metal1 s -1025 6451 -1025 6451 0 FreeSans 3125 0 0 0 G-CLK
flabel metal1 s 8101 7971 8101 7971 0 FreeSans 3125 0 0 0 Q1
flabel metal1 s 16529 7857 16529 7857 0 FreeSans 3125 0 0 0 Q2
flabel metal1 s 25411 7890 25411 7890 0 FreeSans 3125 0 0 0 Q3
flabel metal1 s 34618 7776 34618 7776 0 FreeSans 3125 0 0 0 Q4
flabel metal1 s 43354 7938 43354 7938 0 FreeSans 3125 0 0 0 Q5
flabel metal1 s 52512 7857 52512 7857 0 FreeSans 3125 0 0 0 Q6
flabel metal1 s 62011 8247 62011 8247 0 FreeSans 3125 0 0 0 Q7
flabel locali s 22073 7310 22073 7310 0 FreeSans 3125 0 0 0 VSS
flabel locali s 60613 7795 60613 7795 0 FreeSans 3125 0 0 0 VDD
flabel locali s -679 -1308 -679 -1308 0 FreeSans 3125 0 0 0 D2_1
flabel locali s 27 -1521 27 -1521 0 FreeSans 3125 0 0 0 D2_2
flabel locali s 619 -1751 619 -1751 0 FreeSans 3125 0 0 0 D2_3
flabel locali s 1358 -1998 1358 -1998 0 FreeSans 3125 0 0 0 D2_4
flabel locali s 1752 -2277 1752 -2277 0 FreeSans 3125 0 0 0 D2_5
flabel locali s 2097 -2589 2097 -2589 0 FreeSans 3125 0 0 0 D2_6
flabel locali s 2212 -2917 2212 -2917 0 FreeSans 3125 0 0 0 D2_7
flabel metal1 s -8865 6018 -8865 6018 0 FreeSans 3125 0 0 0 LD
<< end >>
